module SRAM(
  input          clock,
  input          io_en,
  input  [8:0]   io_addr,
  input  [273:0] io_wdata,
  input          io_wen,
  output [273:0] io_rdata
);
`ifdef RANDOMIZE_MEM_INIT
  reg [287:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [273:0] array [0:511]; // @[SRAM.scala 13:26]
  wire  array_io_rdata_MPORT_en; // @[SRAM.scala 13:26]
  wire [8:0] array_io_rdata_MPORT_addr; // @[SRAM.scala 13:26]
  wire [273:0] array_io_rdata_MPORT_data; // @[SRAM.scala 13:26]
  wire [273:0] array_MPORT_data; // @[SRAM.scala 13:26]
  wire [8:0] array_MPORT_addr; // @[SRAM.scala 13:26]
  wire  array_MPORT_mask; // @[SRAM.scala 13:26]
  wire  array_MPORT_en; // @[SRAM.scala 13:26]
  reg  array_io_rdata_MPORT_en_pipe_0;
  reg [8:0] array_io_rdata_MPORT_addr_pipe_0;
  reg  io_rdata_REG; // @[SRAM.scala 15:26]
  assign array_io_rdata_MPORT_en = array_io_rdata_MPORT_en_pipe_0;
  assign array_io_rdata_MPORT_addr = array_io_rdata_MPORT_addr_pipe_0;
  assign array_io_rdata_MPORT_data = array[array_io_rdata_MPORT_addr]; // @[SRAM.scala 13:26]
  assign array_MPORT_data = io_wdata;
  assign array_MPORT_addr = io_addr;
  assign array_MPORT_mask = 1'h1;
  assign array_MPORT_en = io_en & io_wen;
  assign io_rdata = io_rdata_REG ? array_io_rdata_MPORT_data : 274'h0; // @[SRAM.scala 15:18]
  always @(posedge clock) begin
    if (array_MPORT_en & array_MPORT_mask) begin
      array[array_MPORT_addr] <= array_MPORT_data; // @[SRAM.scala 13:26]
    end
    array_io_rdata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      array_io_rdata_MPORT_addr_pipe_0 <= io_addr;
    end
    io_rdata_REG <= io_en; // @[SRAM.scala 15:26]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {9{`RANDOM}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    array[initvar] = _RAND_0[273:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  array_io_rdata_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  array_io_rdata_MPORT_addr_pipe_0 = _RAND_2[8:0];
  _RAND_3 = {1{`RANDOM}};
  io_rdata_REG = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ICache(
  input          clock,
  input          reset,
  input          auto_out_a_ready,
  output         auto_out_a_valid,
  output [1:0]   auto_out_a_bits_source,
  output [31:0]  auto_out_a_bits_address,
  output         auto_out_d_ready,
  input          auto_out_d_valid,
  input  [255:0] auto_out_d_bits_data,
  output         io_cache_req_ready,
  input          io_cache_req_valid,
  input  [38:0]  io_cache_req_bits_addr,
  input          io_cache_resp_ready,
  output         io_cache_resp_valid,
  output [63:0]  io_cache_resp_bits_rdata,
  input          io_fence_i
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [287:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [63:0] _RAND_517;
  reg [255:0] _RAND_518;
  reg [31:0] _RAND_519;
`endif // RANDOMIZE_REG_INIT
  wire  array_clock; // @[ICache.scala 50:21]
  wire  array_io_en; // @[ICache.scala 50:21]
  wire [8:0] array_io_addr; // @[ICache.scala 50:21]
  wire [273:0] array_io_wdata; // @[ICache.scala 50:21]
  wire  array_io_wen; // @[ICache.scala 50:21]
  wire [273:0] array_io_rdata; // @[ICache.scala 50:21]
  reg [38:0] req_r_addr; // @[ICache.scala 48:22]
  reg  valid_0; // @[ICache.scala 51:22]
  reg  valid_1; // @[ICache.scala 51:22]
  reg  valid_2; // @[ICache.scala 51:22]
  reg  valid_3; // @[ICache.scala 51:22]
  reg  valid_4; // @[ICache.scala 51:22]
  reg  valid_5; // @[ICache.scala 51:22]
  reg  valid_6; // @[ICache.scala 51:22]
  reg  valid_7; // @[ICache.scala 51:22]
  reg  valid_8; // @[ICache.scala 51:22]
  reg  valid_9; // @[ICache.scala 51:22]
  reg  valid_10; // @[ICache.scala 51:22]
  reg  valid_11; // @[ICache.scala 51:22]
  reg  valid_12; // @[ICache.scala 51:22]
  reg  valid_13; // @[ICache.scala 51:22]
  reg  valid_14; // @[ICache.scala 51:22]
  reg  valid_15; // @[ICache.scala 51:22]
  reg  valid_16; // @[ICache.scala 51:22]
  reg  valid_17; // @[ICache.scala 51:22]
  reg  valid_18; // @[ICache.scala 51:22]
  reg  valid_19; // @[ICache.scala 51:22]
  reg  valid_20; // @[ICache.scala 51:22]
  reg  valid_21; // @[ICache.scala 51:22]
  reg  valid_22; // @[ICache.scala 51:22]
  reg  valid_23; // @[ICache.scala 51:22]
  reg  valid_24; // @[ICache.scala 51:22]
  reg  valid_25; // @[ICache.scala 51:22]
  reg  valid_26; // @[ICache.scala 51:22]
  reg  valid_27; // @[ICache.scala 51:22]
  reg  valid_28; // @[ICache.scala 51:22]
  reg  valid_29; // @[ICache.scala 51:22]
  reg  valid_30; // @[ICache.scala 51:22]
  reg  valid_31; // @[ICache.scala 51:22]
  reg  valid_32; // @[ICache.scala 51:22]
  reg  valid_33; // @[ICache.scala 51:22]
  reg  valid_34; // @[ICache.scala 51:22]
  reg  valid_35; // @[ICache.scala 51:22]
  reg  valid_36; // @[ICache.scala 51:22]
  reg  valid_37; // @[ICache.scala 51:22]
  reg  valid_38; // @[ICache.scala 51:22]
  reg  valid_39; // @[ICache.scala 51:22]
  reg  valid_40; // @[ICache.scala 51:22]
  reg  valid_41; // @[ICache.scala 51:22]
  reg  valid_42; // @[ICache.scala 51:22]
  reg  valid_43; // @[ICache.scala 51:22]
  reg  valid_44; // @[ICache.scala 51:22]
  reg  valid_45; // @[ICache.scala 51:22]
  reg  valid_46; // @[ICache.scala 51:22]
  reg  valid_47; // @[ICache.scala 51:22]
  reg  valid_48; // @[ICache.scala 51:22]
  reg  valid_49; // @[ICache.scala 51:22]
  reg  valid_50; // @[ICache.scala 51:22]
  reg  valid_51; // @[ICache.scala 51:22]
  reg  valid_52; // @[ICache.scala 51:22]
  reg  valid_53; // @[ICache.scala 51:22]
  reg  valid_54; // @[ICache.scala 51:22]
  reg  valid_55; // @[ICache.scala 51:22]
  reg  valid_56; // @[ICache.scala 51:22]
  reg  valid_57; // @[ICache.scala 51:22]
  reg  valid_58; // @[ICache.scala 51:22]
  reg  valid_59; // @[ICache.scala 51:22]
  reg  valid_60; // @[ICache.scala 51:22]
  reg  valid_61; // @[ICache.scala 51:22]
  reg  valid_62; // @[ICache.scala 51:22]
  reg  valid_63; // @[ICache.scala 51:22]
  reg  valid_64; // @[ICache.scala 51:22]
  reg  valid_65; // @[ICache.scala 51:22]
  reg  valid_66; // @[ICache.scala 51:22]
  reg  valid_67; // @[ICache.scala 51:22]
  reg  valid_68; // @[ICache.scala 51:22]
  reg  valid_69; // @[ICache.scala 51:22]
  reg  valid_70; // @[ICache.scala 51:22]
  reg  valid_71; // @[ICache.scala 51:22]
  reg  valid_72; // @[ICache.scala 51:22]
  reg  valid_73; // @[ICache.scala 51:22]
  reg  valid_74; // @[ICache.scala 51:22]
  reg  valid_75; // @[ICache.scala 51:22]
  reg  valid_76; // @[ICache.scala 51:22]
  reg  valid_77; // @[ICache.scala 51:22]
  reg  valid_78; // @[ICache.scala 51:22]
  reg  valid_79; // @[ICache.scala 51:22]
  reg  valid_80; // @[ICache.scala 51:22]
  reg  valid_81; // @[ICache.scala 51:22]
  reg  valid_82; // @[ICache.scala 51:22]
  reg  valid_83; // @[ICache.scala 51:22]
  reg  valid_84; // @[ICache.scala 51:22]
  reg  valid_85; // @[ICache.scala 51:22]
  reg  valid_86; // @[ICache.scala 51:22]
  reg  valid_87; // @[ICache.scala 51:22]
  reg  valid_88; // @[ICache.scala 51:22]
  reg  valid_89; // @[ICache.scala 51:22]
  reg  valid_90; // @[ICache.scala 51:22]
  reg  valid_91; // @[ICache.scala 51:22]
  reg  valid_92; // @[ICache.scala 51:22]
  reg  valid_93; // @[ICache.scala 51:22]
  reg  valid_94; // @[ICache.scala 51:22]
  reg  valid_95; // @[ICache.scala 51:22]
  reg  valid_96; // @[ICache.scala 51:22]
  reg  valid_97; // @[ICache.scala 51:22]
  reg  valid_98; // @[ICache.scala 51:22]
  reg  valid_99; // @[ICache.scala 51:22]
  reg  valid_100; // @[ICache.scala 51:22]
  reg  valid_101; // @[ICache.scala 51:22]
  reg  valid_102; // @[ICache.scala 51:22]
  reg  valid_103; // @[ICache.scala 51:22]
  reg  valid_104; // @[ICache.scala 51:22]
  reg  valid_105; // @[ICache.scala 51:22]
  reg  valid_106; // @[ICache.scala 51:22]
  reg  valid_107; // @[ICache.scala 51:22]
  reg  valid_108; // @[ICache.scala 51:22]
  reg  valid_109; // @[ICache.scala 51:22]
  reg  valid_110; // @[ICache.scala 51:22]
  reg  valid_111; // @[ICache.scala 51:22]
  reg  valid_112; // @[ICache.scala 51:22]
  reg  valid_113; // @[ICache.scala 51:22]
  reg  valid_114; // @[ICache.scala 51:22]
  reg  valid_115; // @[ICache.scala 51:22]
  reg  valid_116; // @[ICache.scala 51:22]
  reg  valid_117; // @[ICache.scala 51:22]
  reg  valid_118; // @[ICache.scala 51:22]
  reg  valid_119; // @[ICache.scala 51:22]
  reg  valid_120; // @[ICache.scala 51:22]
  reg  valid_121; // @[ICache.scala 51:22]
  reg  valid_122; // @[ICache.scala 51:22]
  reg  valid_123; // @[ICache.scala 51:22]
  reg  valid_124; // @[ICache.scala 51:22]
  reg  valid_125; // @[ICache.scala 51:22]
  reg  valid_126; // @[ICache.scala 51:22]
  reg  valid_127; // @[ICache.scala 51:22]
  reg  valid_128; // @[ICache.scala 51:22]
  reg  valid_129; // @[ICache.scala 51:22]
  reg  valid_130; // @[ICache.scala 51:22]
  reg  valid_131; // @[ICache.scala 51:22]
  reg  valid_132; // @[ICache.scala 51:22]
  reg  valid_133; // @[ICache.scala 51:22]
  reg  valid_134; // @[ICache.scala 51:22]
  reg  valid_135; // @[ICache.scala 51:22]
  reg  valid_136; // @[ICache.scala 51:22]
  reg  valid_137; // @[ICache.scala 51:22]
  reg  valid_138; // @[ICache.scala 51:22]
  reg  valid_139; // @[ICache.scala 51:22]
  reg  valid_140; // @[ICache.scala 51:22]
  reg  valid_141; // @[ICache.scala 51:22]
  reg  valid_142; // @[ICache.scala 51:22]
  reg  valid_143; // @[ICache.scala 51:22]
  reg  valid_144; // @[ICache.scala 51:22]
  reg  valid_145; // @[ICache.scala 51:22]
  reg  valid_146; // @[ICache.scala 51:22]
  reg  valid_147; // @[ICache.scala 51:22]
  reg  valid_148; // @[ICache.scala 51:22]
  reg  valid_149; // @[ICache.scala 51:22]
  reg  valid_150; // @[ICache.scala 51:22]
  reg  valid_151; // @[ICache.scala 51:22]
  reg  valid_152; // @[ICache.scala 51:22]
  reg  valid_153; // @[ICache.scala 51:22]
  reg  valid_154; // @[ICache.scala 51:22]
  reg  valid_155; // @[ICache.scala 51:22]
  reg  valid_156; // @[ICache.scala 51:22]
  reg  valid_157; // @[ICache.scala 51:22]
  reg  valid_158; // @[ICache.scala 51:22]
  reg  valid_159; // @[ICache.scala 51:22]
  reg  valid_160; // @[ICache.scala 51:22]
  reg  valid_161; // @[ICache.scala 51:22]
  reg  valid_162; // @[ICache.scala 51:22]
  reg  valid_163; // @[ICache.scala 51:22]
  reg  valid_164; // @[ICache.scala 51:22]
  reg  valid_165; // @[ICache.scala 51:22]
  reg  valid_166; // @[ICache.scala 51:22]
  reg  valid_167; // @[ICache.scala 51:22]
  reg  valid_168; // @[ICache.scala 51:22]
  reg  valid_169; // @[ICache.scala 51:22]
  reg  valid_170; // @[ICache.scala 51:22]
  reg  valid_171; // @[ICache.scala 51:22]
  reg  valid_172; // @[ICache.scala 51:22]
  reg  valid_173; // @[ICache.scala 51:22]
  reg  valid_174; // @[ICache.scala 51:22]
  reg  valid_175; // @[ICache.scala 51:22]
  reg  valid_176; // @[ICache.scala 51:22]
  reg  valid_177; // @[ICache.scala 51:22]
  reg  valid_178; // @[ICache.scala 51:22]
  reg  valid_179; // @[ICache.scala 51:22]
  reg  valid_180; // @[ICache.scala 51:22]
  reg  valid_181; // @[ICache.scala 51:22]
  reg  valid_182; // @[ICache.scala 51:22]
  reg  valid_183; // @[ICache.scala 51:22]
  reg  valid_184; // @[ICache.scala 51:22]
  reg  valid_185; // @[ICache.scala 51:22]
  reg  valid_186; // @[ICache.scala 51:22]
  reg  valid_187; // @[ICache.scala 51:22]
  reg  valid_188; // @[ICache.scala 51:22]
  reg  valid_189; // @[ICache.scala 51:22]
  reg  valid_190; // @[ICache.scala 51:22]
  reg  valid_191; // @[ICache.scala 51:22]
  reg  valid_192; // @[ICache.scala 51:22]
  reg  valid_193; // @[ICache.scala 51:22]
  reg  valid_194; // @[ICache.scala 51:22]
  reg  valid_195; // @[ICache.scala 51:22]
  reg  valid_196; // @[ICache.scala 51:22]
  reg  valid_197; // @[ICache.scala 51:22]
  reg  valid_198; // @[ICache.scala 51:22]
  reg  valid_199; // @[ICache.scala 51:22]
  reg  valid_200; // @[ICache.scala 51:22]
  reg  valid_201; // @[ICache.scala 51:22]
  reg  valid_202; // @[ICache.scala 51:22]
  reg  valid_203; // @[ICache.scala 51:22]
  reg  valid_204; // @[ICache.scala 51:22]
  reg  valid_205; // @[ICache.scala 51:22]
  reg  valid_206; // @[ICache.scala 51:22]
  reg  valid_207; // @[ICache.scala 51:22]
  reg  valid_208; // @[ICache.scala 51:22]
  reg  valid_209; // @[ICache.scala 51:22]
  reg  valid_210; // @[ICache.scala 51:22]
  reg  valid_211; // @[ICache.scala 51:22]
  reg  valid_212; // @[ICache.scala 51:22]
  reg  valid_213; // @[ICache.scala 51:22]
  reg  valid_214; // @[ICache.scala 51:22]
  reg  valid_215; // @[ICache.scala 51:22]
  reg  valid_216; // @[ICache.scala 51:22]
  reg  valid_217; // @[ICache.scala 51:22]
  reg  valid_218; // @[ICache.scala 51:22]
  reg  valid_219; // @[ICache.scala 51:22]
  reg  valid_220; // @[ICache.scala 51:22]
  reg  valid_221; // @[ICache.scala 51:22]
  reg  valid_222; // @[ICache.scala 51:22]
  reg  valid_223; // @[ICache.scala 51:22]
  reg  valid_224; // @[ICache.scala 51:22]
  reg  valid_225; // @[ICache.scala 51:22]
  reg  valid_226; // @[ICache.scala 51:22]
  reg  valid_227; // @[ICache.scala 51:22]
  reg  valid_228; // @[ICache.scala 51:22]
  reg  valid_229; // @[ICache.scala 51:22]
  reg  valid_230; // @[ICache.scala 51:22]
  reg  valid_231; // @[ICache.scala 51:22]
  reg  valid_232; // @[ICache.scala 51:22]
  reg  valid_233; // @[ICache.scala 51:22]
  reg  valid_234; // @[ICache.scala 51:22]
  reg  valid_235; // @[ICache.scala 51:22]
  reg  valid_236; // @[ICache.scala 51:22]
  reg  valid_237; // @[ICache.scala 51:22]
  reg  valid_238; // @[ICache.scala 51:22]
  reg  valid_239; // @[ICache.scala 51:22]
  reg  valid_240; // @[ICache.scala 51:22]
  reg  valid_241; // @[ICache.scala 51:22]
  reg  valid_242; // @[ICache.scala 51:22]
  reg  valid_243; // @[ICache.scala 51:22]
  reg  valid_244; // @[ICache.scala 51:22]
  reg  valid_245; // @[ICache.scala 51:22]
  reg  valid_246; // @[ICache.scala 51:22]
  reg  valid_247; // @[ICache.scala 51:22]
  reg  valid_248; // @[ICache.scala 51:22]
  reg  valid_249; // @[ICache.scala 51:22]
  reg  valid_250; // @[ICache.scala 51:22]
  reg  valid_251; // @[ICache.scala 51:22]
  reg  valid_252; // @[ICache.scala 51:22]
  reg  valid_253; // @[ICache.scala 51:22]
  reg  valid_254; // @[ICache.scala 51:22]
  reg  valid_255; // @[ICache.scala 51:22]
  reg  valid_256; // @[ICache.scala 51:22]
  reg  valid_257; // @[ICache.scala 51:22]
  reg  valid_258; // @[ICache.scala 51:22]
  reg  valid_259; // @[ICache.scala 51:22]
  reg  valid_260; // @[ICache.scala 51:22]
  reg  valid_261; // @[ICache.scala 51:22]
  reg  valid_262; // @[ICache.scala 51:22]
  reg  valid_263; // @[ICache.scala 51:22]
  reg  valid_264; // @[ICache.scala 51:22]
  reg  valid_265; // @[ICache.scala 51:22]
  reg  valid_266; // @[ICache.scala 51:22]
  reg  valid_267; // @[ICache.scala 51:22]
  reg  valid_268; // @[ICache.scala 51:22]
  reg  valid_269; // @[ICache.scala 51:22]
  reg  valid_270; // @[ICache.scala 51:22]
  reg  valid_271; // @[ICache.scala 51:22]
  reg  valid_272; // @[ICache.scala 51:22]
  reg  valid_273; // @[ICache.scala 51:22]
  reg  valid_274; // @[ICache.scala 51:22]
  reg  valid_275; // @[ICache.scala 51:22]
  reg  valid_276; // @[ICache.scala 51:22]
  reg  valid_277; // @[ICache.scala 51:22]
  reg  valid_278; // @[ICache.scala 51:22]
  reg  valid_279; // @[ICache.scala 51:22]
  reg  valid_280; // @[ICache.scala 51:22]
  reg  valid_281; // @[ICache.scala 51:22]
  reg  valid_282; // @[ICache.scala 51:22]
  reg  valid_283; // @[ICache.scala 51:22]
  reg  valid_284; // @[ICache.scala 51:22]
  reg  valid_285; // @[ICache.scala 51:22]
  reg  valid_286; // @[ICache.scala 51:22]
  reg  valid_287; // @[ICache.scala 51:22]
  reg  valid_288; // @[ICache.scala 51:22]
  reg  valid_289; // @[ICache.scala 51:22]
  reg  valid_290; // @[ICache.scala 51:22]
  reg  valid_291; // @[ICache.scala 51:22]
  reg  valid_292; // @[ICache.scala 51:22]
  reg  valid_293; // @[ICache.scala 51:22]
  reg  valid_294; // @[ICache.scala 51:22]
  reg  valid_295; // @[ICache.scala 51:22]
  reg  valid_296; // @[ICache.scala 51:22]
  reg  valid_297; // @[ICache.scala 51:22]
  reg  valid_298; // @[ICache.scala 51:22]
  reg  valid_299; // @[ICache.scala 51:22]
  reg  valid_300; // @[ICache.scala 51:22]
  reg  valid_301; // @[ICache.scala 51:22]
  reg  valid_302; // @[ICache.scala 51:22]
  reg  valid_303; // @[ICache.scala 51:22]
  reg  valid_304; // @[ICache.scala 51:22]
  reg  valid_305; // @[ICache.scala 51:22]
  reg  valid_306; // @[ICache.scala 51:22]
  reg  valid_307; // @[ICache.scala 51:22]
  reg  valid_308; // @[ICache.scala 51:22]
  reg  valid_309; // @[ICache.scala 51:22]
  reg  valid_310; // @[ICache.scala 51:22]
  reg  valid_311; // @[ICache.scala 51:22]
  reg  valid_312; // @[ICache.scala 51:22]
  reg  valid_313; // @[ICache.scala 51:22]
  reg  valid_314; // @[ICache.scala 51:22]
  reg  valid_315; // @[ICache.scala 51:22]
  reg  valid_316; // @[ICache.scala 51:22]
  reg  valid_317; // @[ICache.scala 51:22]
  reg  valid_318; // @[ICache.scala 51:22]
  reg  valid_319; // @[ICache.scala 51:22]
  reg  valid_320; // @[ICache.scala 51:22]
  reg  valid_321; // @[ICache.scala 51:22]
  reg  valid_322; // @[ICache.scala 51:22]
  reg  valid_323; // @[ICache.scala 51:22]
  reg  valid_324; // @[ICache.scala 51:22]
  reg  valid_325; // @[ICache.scala 51:22]
  reg  valid_326; // @[ICache.scala 51:22]
  reg  valid_327; // @[ICache.scala 51:22]
  reg  valid_328; // @[ICache.scala 51:22]
  reg  valid_329; // @[ICache.scala 51:22]
  reg  valid_330; // @[ICache.scala 51:22]
  reg  valid_331; // @[ICache.scala 51:22]
  reg  valid_332; // @[ICache.scala 51:22]
  reg  valid_333; // @[ICache.scala 51:22]
  reg  valid_334; // @[ICache.scala 51:22]
  reg  valid_335; // @[ICache.scala 51:22]
  reg  valid_336; // @[ICache.scala 51:22]
  reg  valid_337; // @[ICache.scala 51:22]
  reg  valid_338; // @[ICache.scala 51:22]
  reg  valid_339; // @[ICache.scala 51:22]
  reg  valid_340; // @[ICache.scala 51:22]
  reg  valid_341; // @[ICache.scala 51:22]
  reg  valid_342; // @[ICache.scala 51:22]
  reg  valid_343; // @[ICache.scala 51:22]
  reg  valid_344; // @[ICache.scala 51:22]
  reg  valid_345; // @[ICache.scala 51:22]
  reg  valid_346; // @[ICache.scala 51:22]
  reg  valid_347; // @[ICache.scala 51:22]
  reg  valid_348; // @[ICache.scala 51:22]
  reg  valid_349; // @[ICache.scala 51:22]
  reg  valid_350; // @[ICache.scala 51:22]
  reg  valid_351; // @[ICache.scala 51:22]
  reg  valid_352; // @[ICache.scala 51:22]
  reg  valid_353; // @[ICache.scala 51:22]
  reg  valid_354; // @[ICache.scala 51:22]
  reg  valid_355; // @[ICache.scala 51:22]
  reg  valid_356; // @[ICache.scala 51:22]
  reg  valid_357; // @[ICache.scala 51:22]
  reg  valid_358; // @[ICache.scala 51:22]
  reg  valid_359; // @[ICache.scala 51:22]
  reg  valid_360; // @[ICache.scala 51:22]
  reg  valid_361; // @[ICache.scala 51:22]
  reg  valid_362; // @[ICache.scala 51:22]
  reg  valid_363; // @[ICache.scala 51:22]
  reg  valid_364; // @[ICache.scala 51:22]
  reg  valid_365; // @[ICache.scala 51:22]
  reg  valid_366; // @[ICache.scala 51:22]
  reg  valid_367; // @[ICache.scala 51:22]
  reg  valid_368; // @[ICache.scala 51:22]
  reg  valid_369; // @[ICache.scala 51:22]
  reg  valid_370; // @[ICache.scala 51:22]
  reg  valid_371; // @[ICache.scala 51:22]
  reg  valid_372; // @[ICache.scala 51:22]
  reg  valid_373; // @[ICache.scala 51:22]
  reg  valid_374; // @[ICache.scala 51:22]
  reg  valid_375; // @[ICache.scala 51:22]
  reg  valid_376; // @[ICache.scala 51:22]
  reg  valid_377; // @[ICache.scala 51:22]
  reg  valid_378; // @[ICache.scala 51:22]
  reg  valid_379; // @[ICache.scala 51:22]
  reg  valid_380; // @[ICache.scala 51:22]
  reg  valid_381; // @[ICache.scala 51:22]
  reg  valid_382; // @[ICache.scala 51:22]
  reg  valid_383; // @[ICache.scala 51:22]
  reg  valid_384; // @[ICache.scala 51:22]
  reg  valid_385; // @[ICache.scala 51:22]
  reg  valid_386; // @[ICache.scala 51:22]
  reg  valid_387; // @[ICache.scala 51:22]
  reg  valid_388; // @[ICache.scala 51:22]
  reg  valid_389; // @[ICache.scala 51:22]
  reg  valid_390; // @[ICache.scala 51:22]
  reg  valid_391; // @[ICache.scala 51:22]
  reg  valid_392; // @[ICache.scala 51:22]
  reg  valid_393; // @[ICache.scala 51:22]
  reg  valid_394; // @[ICache.scala 51:22]
  reg  valid_395; // @[ICache.scala 51:22]
  reg  valid_396; // @[ICache.scala 51:22]
  reg  valid_397; // @[ICache.scala 51:22]
  reg  valid_398; // @[ICache.scala 51:22]
  reg  valid_399; // @[ICache.scala 51:22]
  reg  valid_400; // @[ICache.scala 51:22]
  reg  valid_401; // @[ICache.scala 51:22]
  reg  valid_402; // @[ICache.scala 51:22]
  reg  valid_403; // @[ICache.scala 51:22]
  reg  valid_404; // @[ICache.scala 51:22]
  reg  valid_405; // @[ICache.scala 51:22]
  reg  valid_406; // @[ICache.scala 51:22]
  reg  valid_407; // @[ICache.scala 51:22]
  reg  valid_408; // @[ICache.scala 51:22]
  reg  valid_409; // @[ICache.scala 51:22]
  reg  valid_410; // @[ICache.scala 51:22]
  reg  valid_411; // @[ICache.scala 51:22]
  reg  valid_412; // @[ICache.scala 51:22]
  reg  valid_413; // @[ICache.scala 51:22]
  reg  valid_414; // @[ICache.scala 51:22]
  reg  valid_415; // @[ICache.scala 51:22]
  reg  valid_416; // @[ICache.scala 51:22]
  reg  valid_417; // @[ICache.scala 51:22]
  reg  valid_418; // @[ICache.scala 51:22]
  reg  valid_419; // @[ICache.scala 51:22]
  reg  valid_420; // @[ICache.scala 51:22]
  reg  valid_421; // @[ICache.scala 51:22]
  reg  valid_422; // @[ICache.scala 51:22]
  reg  valid_423; // @[ICache.scala 51:22]
  reg  valid_424; // @[ICache.scala 51:22]
  reg  valid_425; // @[ICache.scala 51:22]
  reg  valid_426; // @[ICache.scala 51:22]
  reg  valid_427; // @[ICache.scala 51:22]
  reg  valid_428; // @[ICache.scala 51:22]
  reg  valid_429; // @[ICache.scala 51:22]
  reg  valid_430; // @[ICache.scala 51:22]
  reg  valid_431; // @[ICache.scala 51:22]
  reg  valid_432; // @[ICache.scala 51:22]
  reg  valid_433; // @[ICache.scala 51:22]
  reg  valid_434; // @[ICache.scala 51:22]
  reg  valid_435; // @[ICache.scala 51:22]
  reg  valid_436; // @[ICache.scala 51:22]
  reg  valid_437; // @[ICache.scala 51:22]
  reg  valid_438; // @[ICache.scala 51:22]
  reg  valid_439; // @[ICache.scala 51:22]
  reg  valid_440; // @[ICache.scala 51:22]
  reg  valid_441; // @[ICache.scala 51:22]
  reg  valid_442; // @[ICache.scala 51:22]
  reg  valid_443; // @[ICache.scala 51:22]
  reg  valid_444; // @[ICache.scala 51:22]
  reg  valid_445; // @[ICache.scala 51:22]
  reg  valid_446; // @[ICache.scala 51:22]
  reg  valid_447; // @[ICache.scala 51:22]
  reg  valid_448; // @[ICache.scala 51:22]
  reg  valid_449; // @[ICache.scala 51:22]
  reg  valid_450; // @[ICache.scala 51:22]
  reg  valid_451; // @[ICache.scala 51:22]
  reg  valid_452; // @[ICache.scala 51:22]
  reg  valid_453; // @[ICache.scala 51:22]
  reg  valid_454; // @[ICache.scala 51:22]
  reg  valid_455; // @[ICache.scala 51:22]
  reg  valid_456; // @[ICache.scala 51:22]
  reg  valid_457; // @[ICache.scala 51:22]
  reg  valid_458; // @[ICache.scala 51:22]
  reg  valid_459; // @[ICache.scala 51:22]
  reg  valid_460; // @[ICache.scala 51:22]
  reg  valid_461; // @[ICache.scala 51:22]
  reg  valid_462; // @[ICache.scala 51:22]
  reg  valid_463; // @[ICache.scala 51:22]
  reg  valid_464; // @[ICache.scala 51:22]
  reg  valid_465; // @[ICache.scala 51:22]
  reg  valid_466; // @[ICache.scala 51:22]
  reg  valid_467; // @[ICache.scala 51:22]
  reg  valid_468; // @[ICache.scala 51:22]
  reg  valid_469; // @[ICache.scala 51:22]
  reg  valid_470; // @[ICache.scala 51:22]
  reg  valid_471; // @[ICache.scala 51:22]
  reg  valid_472; // @[ICache.scala 51:22]
  reg  valid_473; // @[ICache.scala 51:22]
  reg  valid_474; // @[ICache.scala 51:22]
  reg  valid_475; // @[ICache.scala 51:22]
  reg  valid_476; // @[ICache.scala 51:22]
  reg  valid_477; // @[ICache.scala 51:22]
  reg  valid_478; // @[ICache.scala 51:22]
  reg  valid_479; // @[ICache.scala 51:22]
  reg  valid_480; // @[ICache.scala 51:22]
  reg  valid_481; // @[ICache.scala 51:22]
  reg  valid_482; // @[ICache.scala 51:22]
  reg  valid_483; // @[ICache.scala 51:22]
  reg  valid_484; // @[ICache.scala 51:22]
  reg  valid_485; // @[ICache.scala 51:22]
  reg  valid_486; // @[ICache.scala 51:22]
  reg  valid_487; // @[ICache.scala 51:22]
  reg  valid_488; // @[ICache.scala 51:22]
  reg  valid_489; // @[ICache.scala 51:22]
  reg  valid_490; // @[ICache.scala 51:22]
  reg  valid_491; // @[ICache.scala 51:22]
  reg  valid_492; // @[ICache.scala 51:22]
  reg  valid_493; // @[ICache.scala 51:22]
  reg  valid_494; // @[ICache.scala 51:22]
  reg  valid_495; // @[ICache.scala 51:22]
  reg  valid_496; // @[ICache.scala 51:22]
  reg  valid_497; // @[ICache.scala 51:22]
  reg  valid_498; // @[ICache.scala 51:22]
  reg  valid_499; // @[ICache.scala 51:22]
  reg  valid_500; // @[ICache.scala 51:22]
  reg  valid_501; // @[ICache.scala 51:22]
  reg  valid_502; // @[ICache.scala 51:22]
  reg  valid_503; // @[ICache.scala 51:22]
  reg  valid_504; // @[ICache.scala 51:22]
  reg  valid_505; // @[ICache.scala 51:22]
  reg  valid_506; // @[ICache.scala 51:22]
  reg  valid_507; // @[ICache.scala 51:22]
  reg  valid_508; // @[ICache.scala 51:22]
  reg  valid_509; // @[ICache.scala 51:22]
  reg  valid_510; // @[ICache.scala 51:22]
  reg  valid_511; // @[ICache.scala 51:22]
  reg [2:0] state; // @[ICache.scala 78:68]
  wire  _GEN_2 = 9'h1 == req_r_addr[13:5] ? valid_1 : valid_0; // @[ICache.scala 68:{44,44}]
  wire  _GEN_3 = 9'h2 == req_r_addr[13:5] ? valid_2 : _GEN_2; // @[ICache.scala 68:{44,44}]
  wire  _GEN_4 = 9'h3 == req_r_addr[13:5] ? valid_3 : _GEN_3; // @[ICache.scala 68:{44,44}]
  wire  _GEN_5 = 9'h4 == req_r_addr[13:5] ? valid_4 : _GEN_4; // @[ICache.scala 68:{44,44}]
  wire  _GEN_6 = 9'h5 == req_r_addr[13:5] ? valid_5 : _GEN_5; // @[ICache.scala 68:{44,44}]
  wire  _GEN_7 = 9'h6 == req_r_addr[13:5] ? valid_6 : _GEN_6; // @[ICache.scala 68:{44,44}]
  wire  _GEN_8 = 9'h7 == req_r_addr[13:5] ? valid_7 : _GEN_7; // @[ICache.scala 68:{44,44}]
  wire  _GEN_9 = 9'h8 == req_r_addr[13:5] ? valid_8 : _GEN_8; // @[ICache.scala 68:{44,44}]
  wire  _GEN_10 = 9'h9 == req_r_addr[13:5] ? valid_9 : _GEN_9; // @[ICache.scala 68:{44,44}]
  wire  _GEN_11 = 9'ha == req_r_addr[13:5] ? valid_10 : _GEN_10; // @[ICache.scala 68:{44,44}]
  wire  _GEN_12 = 9'hb == req_r_addr[13:5] ? valid_11 : _GEN_11; // @[ICache.scala 68:{44,44}]
  wire  _GEN_13 = 9'hc == req_r_addr[13:5] ? valid_12 : _GEN_12; // @[ICache.scala 68:{44,44}]
  wire  _GEN_14 = 9'hd == req_r_addr[13:5] ? valid_13 : _GEN_13; // @[ICache.scala 68:{44,44}]
  wire  _GEN_15 = 9'he == req_r_addr[13:5] ? valid_14 : _GEN_14; // @[ICache.scala 68:{44,44}]
  wire  _GEN_16 = 9'hf == req_r_addr[13:5] ? valid_15 : _GEN_15; // @[ICache.scala 68:{44,44}]
  wire  _GEN_17 = 9'h10 == req_r_addr[13:5] ? valid_16 : _GEN_16; // @[ICache.scala 68:{44,44}]
  wire  _GEN_18 = 9'h11 == req_r_addr[13:5] ? valid_17 : _GEN_17; // @[ICache.scala 68:{44,44}]
  wire  _GEN_19 = 9'h12 == req_r_addr[13:5] ? valid_18 : _GEN_18; // @[ICache.scala 68:{44,44}]
  wire  _GEN_20 = 9'h13 == req_r_addr[13:5] ? valid_19 : _GEN_19; // @[ICache.scala 68:{44,44}]
  wire  _GEN_21 = 9'h14 == req_r_addr[13:5] ? valid_20 : _GEN_20; // @[ICache.scala 68:{44,44}]
  wire  _GEN_22 = 9'h15 == req_r_addr[13:5] ? valid_21 : _GEN_21; // @[ICache.scala 68:{44,44}]
  wire  _GEN_23 = 9'h16 == req_r_addr[13:5] ? valid_22 : _GEN_22; // @[ICache.scala 68:{44,44}]
  wire  _GEN_24 = 9'h17 == req_r_addr[13:5] ? valid_23 : _GEN_23; // @[ICache.scala 68:{44,44}]
  wire  _GEN_25 = 9'h18 == req_r_addr[13:5] ? valid_24 : _GEN_24; // @[ICache.scala 68:{44,44}]
  wire  _GEN_26 = 9'h19 == req_r_addr[13:5] ? valid_25 : _GEN_25; // @[ICache.scala 68:{44,44}]
  wire  _GEN_27 = 9'h1a == req_r_addr[13:5] ? valid_26 : _GEN_26; // @[ICache.scala 68:{44,44}]
  wire  _GEN_28 = 9'h1b == req_r_addr[13:5] ? valid_27 : _GEN_27; // @[ICache.scala 68:{44,44}]
  wire  _GEN_29 = 9'h1c == req_r_addr[13:5] ? valid_28 : _GEN_28; // @[ICache.scala 68:{44,44}]
  wire  _GEN_30 = 9'h1d == req_r_addr[13:5] ? valid_29 : _GEN_29; // @[ICache.scala 68:{44,44}]
  wire  _GEN_31 = 9'h1e == req_r_addr[13:5] ? valid_30 : _GEN_30; // @[ICache.scala 68:{44,44}]
  wire  _GEN_32 = 9'h1f == req_r_addr[13:5] ? valid_31 : _GEN_31; // @[ICache.scala 68:{44,44}]
  wire  _GEN_33 = 9'h20 == req_r_addr[13:5] ? valid_32 : _GEN_32; // @[ICache.scala 68:{44,44}]
  wire  _GEN_34 = 9'h21 == req_r_addr[13:5] ? valid_33 : _GEN_33; // @[ICache.scala 68:{44,44}]
  wire  _GEN_35 = 9'h22 == req_r_addr[13:5] ? valid_34 : _GEN_34; // @[ICache.scala 68:{44,44}]
  wire  _GEN_36 = 9'h23 == req_r_addr[13:5] ? valid_35 : _GEN_35; // @[ICache.scala 68:{44,44}]
  wire  _GEN_37 = 9'h24 == req_r_addr[13:5] ? valid_36 : _GEN_36; // @[ICache.scala 68:{44,44}]
  wire  _GEN_38 = 9'h25 == req_r_addr[13:5] ? valid_37 : _GEN_37; // @[ICache.scala 68:{44,44}]
  wire  _GEN_39 = 9'h26 == req_r_addr[13:5] ? valid_38 : _GEN_38; // @[ICache.scala 68:{44,44}]
  wire  _GEN_40 = 9'h27 == req_r_addr[13:5] ? valid_39 : _GEN_39; // @[ICache.scala 68:{44,44}]
  wire  _GEN_41 = 9'h28 == req_r_addr[13:5] ? valid_40 : _GEN_40; // @[ICache.scala 68:{44,44}]
  wire  _GEN_42 = 9'h29 == req_r_addr[13:5] ? valid_41 : _GEN_41; // @[ICache.scala 68:{44,44}]
  wire  _GEN_43 = 9'h2a == req_r_addr[13:5] ? valid_42 : _GEN_42; // @[ICache.scala 68:{44,44}]
  wire  _GEN_44 = 9'h2b == req_r_addr[13:5] ? valid_43 : _GEN_43; // @[ICache.scala 68:{44,44}]
  wire  _GEN_45 = 9'h2c == req_r_addr[13:5] ? valid_44 : _GEN_44; // @[ICache.scala 68:{44,44}]
  wire  _GEN_46 = 9'h2d == req_r_addr[13:5] ? valid_45 : _GEN_45; // @[ICache.scala 68:{44,44}]
  wire  _GEN_47 = 9'h2e == req_r_addr[13:5] ? valid_46 : _GEN_46; // @[ICache.scala 68:{44,44}]
  wire  _GEN_48 = 9'h2f == req_r_addr[13:5] ? valid_47 : _GEN_47; // @[ICache.scala 68:{44,44}]
  wire  _GEN_49 = 9'h30 == req_r_addr[13:5] ? valid_48 : _GEN_48; // @[ICache.scala 68:{44,44}]
  wire  _GEN_50 = 9'h31 == req_r_addr[13:5] ? valid_49 : _GEN_49; // @[ICache.scala 68:{44,44}]
  wire  _GEN_51 = 9'h32 == req_r_addr[13:5] ? valid_50 : _GEN_50; // @[ICache.scala 68:{44,44}]
  wire  _GEN_52 = 9'h33 == req_r_addr[13:5] ? valid_51 : _GEN_51; // @[ICache.scala 68:{44,44}]
  wire  _GEN_53 = 9'h34 == req_r_addr[13:5] ? valid_52 : _GEN_52; // @[ICache.scala 68:{44,44}]
  wire  _GEN_54 = 9'h35 == req_r_addr[13:5] ? valid_53 : _GEN_53; // @[ICache.scala 68:{44,44}]
  wire  _GEN_55 = 9'h36 == req_r_addr[13:5] ? valid_54 : _GEN_54; // @[ICache.scala 68:{44,44}]
  wire  _GEN_56 = 9'h37 == req_r_addr[13:5] ? valid_55 : _GEN_55; // @[ICache.scala 68:{44,44}]
  wire  _GEN_57 = 9'h38 == req_r_addr[13:5] ? valid_56 : _GEN_56; // @[ICache.scala 68:{44,44}]
  wire  _GEN_58 = 9'h39 == req_r_addr[13:5] ? valid_57 : _GEN_57; // @[ICache.scala 68:{44,44}]
  wire  _GEN_59 = 9'h3a == req_r_addr[13:5] ? valid_58 : _GEN_58; // @[ICache.scala 68:{44,44}]
  wire  _GEN_60 = 9'h3b == req_r_addr[13:5] ? valid_59 : _GEN_59; // @[ICache.scala 68:{44,44}]
  wire  _GEN_61 = 9'h3c == req_r_addr[13:5] ? valid_60 : _GEN_60; // @[ICache.scala 68:{44,44}]
  wire  _GEN_62 = 9'h3d == req_r_addr[13:5] ? valid_61 : _GEN_61; // @[ICache.scala 68:{44,44}]
  wire  _GEN_63 = 9'h3e == req_r_addr[13:5] ? valid_62 : _GEN_62; // @[ICache.scala 68:{44,44}]
  wire  _GEN_64 = 9'h3f == req_r_addr[13:5] ? valid_63 : _GEN_63; // @[ICache.scala 68:{44,44}]
  wire  _GEN_65 = 9'h40 == req_r_addr[13:5] ? valid_64 : _GEN_64; // @[ICache.scala 68:{44,44}]
  wire  _GEN_66 = 9'h41 == req_r_addr[13:5] ? valid_65 : _GEN_65; // @[ICache.scala 68:{44,44}]
  wire  _GEN_67 = 9'h42 == req_r_addr[13:5] ? valid_66 : _GEN_66; // @[ICache.scala 68:{44,44}]
  wire  _GEN_68 = 9'h43 == req_r_addr[13:5] ? valid_67 : _GEN_67; // @[ICache.scala 68:{44,44}]
  wire  _GEN_69 = 9'h44 == req_r_addr[13:5] ? valid_68 : _GEN_68; // @[ICache.scala 68:{44,44}]
  wire  _GEN_70 = 9'h45 == req_r_addr[13:5] ? valid_69 : _GEN_69; // @[ICache.scala 68:{44,44}]
  wire  _GEN_71 = 9'h46 == req_r_addr[13:5] ? valid_70 : _GEN_70; // @[ICache.scala 68:{44,44}]
  wire  _GEN_72 = 9'h47 == req_r_addr[13:5] ? valid_71 : _GEN_71; // @[ICache.scala 68:{44,44}]
  wire  _GEN_73 = 9'h48 == req_r_addr[13:5] ? valid_72 : _GEN_72; // @[ICache.scala 68:{44,44}]
  wire  _GEN_74 = 9'h49 == req_r_addr[13:5] ? valid_73 : _GEN_73; // @[ICache.scala 68:{44,44}]
  wire  _GEN_75 = 9'h4a == req_r_addr[13:5] ? valid_74 : _GEN_74; // @[ICache.scala 68:{44,44}]
  wire  _GEN_76 = 9'h4b == req_r_addr[13:5] ? valid_75 : _GEN_75; // @[ICache.scala 68:{44,44}]
  wire  _GEN_77 = 9'h4c == req_r_addr[13:5] ? valid_76 : _GEN_76; // @[ICache.scala 68:{44,44}]
  wire  _GEN_78 = 9'h4d == req_r_addr[13:5] ? valid_77 : _GEN_77; // @[ICache.scala 68:{44,44}]
  wire  _GEN_79 = 9'h4e == req_r_addr[13:5] ? valid_78 : _GEN_78; // @[ICache.scala 68:{44,44}]
  wire  _GEN_80 = 9'h4f == req_r_addr[13:5] ? valid_79 : _GEN_79; // @[ICache.scala 68:{44,44}]
  wire  _GEN_81 = 9'h50 == req_r_addr[13:5] ? valid_80 : _GEN_80; // @[ICache.scala 68:{44,44}]
  wire  _GEN_82 = 9'h51 == req_r_addr[13:5] ? valid_81 : _GEN_81; // @[ICache.scala 68:{44,44}]
  wire  _GEN_83 = 9'h52 == req_r_addr[13:5] ? valid_82 : _GEN_82; // @[ICache.scala 68:{44,44}]
  wire  _GEN_84 = 9'h53 == req_r_addr[13:5] ? valid_83 : _GEN_83; // @[ICache.scala 68:{44,44}]
  wire  _GEN_85 = 9'h54 == req_r_addr[13:5] ? valid_84 : _GEN_84; // @[ICache.scala 68:{44,44}]
  wire  _GEN_86 = 9'h55 == req_r_addr[13:5] ? valid_85 : _GEN_85; // @[ICache.scala 68:{44,44}]
  wire  _GEN_87 = 9'h56 == req_r_addr[13:5] ? valid_86 : _GEN_86; // @[ICache.scala 68:{44,44}]
  wire  _GEN_88 = 9'h57 == req_r_addr[13:5] ? valid_87 : _GEN_87; // @[ICache.scala 68:{44,44}]
  wire  _GEN_89 = 9'h58 == req_r_addr[13:5] ? valid_88 : _GEN_88; // @[ICache.scala 68:{44,44}]
  wire  _GEN_90 = 9'h59 == req_r_addr[13:5] ? valid_89 : _GEN_89; // @[ICache.scala 68:{44,44}]
  wire  _GEN_91 = 9'h5a == req_r_addr[13:5] ? valid_90 : _GEN_90; // @[ICache.scala 68:{44,44}]
  wire  _GEN_92 = 9'h5b == req_r_addr[13:5] ? valid_91 : _GEN_91; // @[ICache.scala 68:{44,44}]
  wire  _GEN_93 = 9'h5c == req_r_addr[13:5] ? valid_92 : _GEN_92; // @[ICache.scala 68:{44,44}]
  wire  _GEN_94 = 9'h5d == req_r_addr[13:5] ? valid_93 : _GEN_93; // @[ICache.scala 68:{44,44}]
  wire  _GEN_95 = 9'h5e == req_r_addr[13:5] ? valid_94 : _GEN_94; // @[ICache.scala 68:{44,44}]
  wire  _GEN_96 = 9'h5f == req_r_addr[13:5] ? valid_95 : _GEN_95; // @[ICache.scala 68:{44,44}]
  wire  _GEN_97 = 9'h60 == req_r_addr[13:5] ? valid_96 : _GEN_96; // @[ICache.scala 68:{44,44}]
  wire  _GEN_98 = 9'h61 == req_r_addr[13:5] ? valid_97 : _GEN_97; // @[ICache.scala 68:{44,44}]
  wire  _GEN_99 = 9'h62 == req_r_addr[13:5] ? valid_98 : _GEN_98; // @[ICache.scala 68:{44,44}]
  wire  _GEN_100 = 9'h63 == req_r_addr[13:5] ? valid_99 : _GEN_99; // @[ICache.scala 68:{44,44}]
  wire  _GEN_101 = 9'h64 == req_r_addr[13:5] ? valid_100 : _GEN_100; // @[ICache.scala 68:{44,44}]
  wire  _GEN_102 = 9'h65 == req_r_addr[13:5] ? valid_101 : _GEN_101; // @[ICache.scala 68:{44,44}]
  wire  _GEN_103 = 9'h66 == req_r_addr[13:5] ? valid_102 : _GEN_102; // @[ICache.scala 68:{44,44}]
  wire  _GEN_104 = 9'h67 == req_r_addr[13:5] ? valid_103 : _GEN_103; // @[ICache.scala 68:{44,44}]
  wire  _GEN_105 = 9'h68 == req_r_addr[13:5] ? valid_104 : _GEN_104; // @[ICache.scala 68:{44,44}]
  wire  _GEN_106 = 9'h69 == req_r_addr[13:5] ? valid_105 : _GEN_105; // @[ICache.scala 68:{44,44}]
  wire  _GEN_107 = 9'h6a == req_r_addr[13:5] ? valid_106 : _GEN_106; // @[ICache.scala 68:{44,44}]
  wire  _GEN_108 = 9'h6b == req_r_addr[13:5] ? valid_107 : _GEN_107; // @[ICache.scala 68:{44,44}]
  wire  _GEN_109 = 9'h6c == req_r_addr[13:5] ? valid_108 : _GEN_108; // @[ICache.scala 68:{44,44}]
  wire  _GEN_110 = 9'h6d == req_r_addr[13:5] ? valid_109 : _GEN_109; // @[ICache.scala 68:{44,44}]
  wire  _GEN_111 = 9'h6e == req_r_addr[13:5] ? valid_110 : _GEN_110; // @[ICache.scala 68:{44,44}]
  wire  _GEN_112 = 9'h6f == req_r_addr[13:5] ? valid_111 : _GEN_111; // @[ICache.scala 68:{44,44}]
  wire  _GEN_113 = 9'h70 == req_r_addr[13:5] ? valid_112 : _GEN_112; // @[ICache.scala 68:{44,44}]
  wire  _GEN_114 = 9'h71 == req_r_addr[13:5] ? valid_113 : _GEN_113; // @[ICache.scala 68:{44,44}]
  wire  _GEN_115 = 9'h72 == req_r_addr[13:5] ? valid_114 : _GEN_114; // @[ICache.scala 68:{44,44}]
  wire  _GEN_116 = 9'h73 == req_r_addr[13:5] ? valid_115 : _GEN_115; // @[ICache.scala 68:{44,44}]
  wire  _GEN_117 = 9'h74 == req_r_addr[13:5] ? valid_116 : _GEN_116; // @[ICache.scala 68:{44,44}]
  wire  _GEN_118 = 9'h75 == req_r_addr[13:5] ? valid_117 : _GEN_117; // @[ICache.scala 68:{44,44}]
  wire  _GEN_119 = 9'h76 == req_r_addr[13:5] ? valid_118 : _GEN_118; // @[ICache.scala 68:{44,44}]
  wire  _GEN_120 = 9'h77 == req_r_addr[13:5] ? valid_119 : _GEN_119; // @[ICache.scala 68:{44,44}]
  wire  _GEN_121 = 9'h78 == req_r_addr[13:5] ? valid_120 : _GEN_120; // @[ICache.scala 68:{44,44}]
  wire  _GEN_122 = 9'h79 == req_r_addr[13:5] ? valid_121 : _GEN_121; // @[ICache.scala 68:{44,44}]
  wire  _GEN_123 = 9'h7a == req_r_addr[13:5] ? valid_122 : _GEN_122; // @[ICache.scala 68:{44,44}]
  wire  _GEN_124 = 9'h7b == req_r_addr[13:5] ? valid_123 : _GEN_123; // @[ICache.scala 68:{44,44}]
  wire  _GEN_125 = 9'h7c == req_r_addr[13:5] ? valid_124 : _GEN_124; // @[ICache.scala 68:{44,44}]
  wire  _GEN_126 = 9'h7d == req_r_addr[13:5] ? valid_125 : _GEN_125; // @[ICache.scala 68:{44,44}]
  wire  _GEN_127 = 9'h7e == req_r_addr[13:5] ? valid_126 : _GEN_126; // @[ICache.scala 68:{44,44}]
  wire  _GEN_128 = 9'h7f == req_r_addr[13:5] ? valid_127 : _GEN_127; // @[ICache.scala 68:{44,44}]
  wire  _GEN_129 = 9'h80 == req_r_addr[13:5] ? valid_128 : _GEN_128; // @[ICache.scala 68:{44,44}]
  wire  _GEN_130 = 9'h81 == req_r_addr[13:5] ? valid_129 : _GEN_129; // @[ICache.scala 68:{44,44}]
  wire  _GEN_131 = 9'h82 == req_r_addr[13:5] ? valid_130 : _GEN_130; // @[ICache.scala 68:{44,44}]
  wire  _GEN_132 = 9'h83 == req_r_addr[13:5] ? valid_131 : _GEN_131; // @[ICache.scala 68:{44,44}]
  wire  _GEN_133 = 9'h84 == req_r_addr[13:5] ? valid_132 : _GEN_132; // @[ICache.scala 68:{44,44}]
  wire  _GEN_134 = 9'h85 == req_r_addr[13:5] ? valid_133 : _GEN_133; // @[ICache.scala 68:{44,44}]
  wire  _GEN_135 = 9'h86 == req_r_addr[13:5] ? valid_134 : _GEN_134; // @[ICache.scala 68:{44,44}]
  wire  _GEN_136 = 9'h87 == req_r_addr[13:5] ? valid_135 : _GEN_135; // @[ICache.scala 68:{44,44}]
  wire  _GEN_137 = 9'h88 == req_r_addr[13:5] ? valid_136 : _GEN_136; // @[ICache.scala 68:{44,44}]
  wire  _GEN_138 = 9'h89 == req_r_addr[13:5] ? valid_137 : _GEN_137; // @[ICache.scala 68:{44,44}]
  wire  _GEN_139 = 9'h8a == req_r_addr[13:5] ? valid_138 : _GEN_138; // @[ICache.scala 68:{44,44}]
  wire  _GEN_140 = 9'h8b == req_r_addr[13:5] ? valid_139 : _GEN_139; // @[ICache.scala 68:{44,44}]
  wire  _GEN_141 = 9'h8c == req_r_addr[13:5] ? valid_140 : _GEN_140; // @[ICache.scala 68:{44,44}]
  wire  _GEN_142 = 9'h8d == req_r_addr[13:5] ? valid_141 : _GEN_141; // @[ICache.scala 68:{44,44}]
  wire  _GEN_143 = 9'h8e == req_r_addr[13:5] ? valid_142 : _GEN_142; // @[ICache.scala 68:{44,44}]
  wire  _GEN_144 = 9'h8f == req_r_addr[13:5] ? valid_143 : _GEN_143; // @[ICache.scala 68:{44,44}]
  wire  _GEN_145 = 9'h90 == req_r_addr[13:5] ? valid_144 : _GEN_144; // @[ICache.scala 68:{44,44}]
  wire  _GEN_146 = 9'h91 == req_r_addr[13:5] ? valid_145 : _GEN_145; // @[ICache.scala 68:{44,44}]
  wire  _GEN_147 = 9'h92 == req_r_addr[13:5] ? valid_146 : _GEN_146; // @[ICache.scala 68:{44,44}]
  wire  _GEN_148 = 9'h93 == req_r_addr[13:5] ? valid_147 : _GEN_147; // @[ICache.scala 68:{44,44}]
  wire  _GEN_149 = 9'h94 == req_r_addr[13:5] ? valid_148 : _GEN_148; // @[ICache.scala 68:{44,44}]
  wire  _GEN_150 = 9'h95 == req_r_addr[13:5] ? valid_149 : _GEN_149; // @[ICache.scala 68:{44,44}]
  wire  _GEN_151 = 9'h96 == req_r_addr[13:5] ? valid_150 : _GEN_150; // @[ICache.scala 68:{44,44}]
  wire  _GEN_152 = 9'h97 == req_r_addr[13:5] ? valid_151 : _GEN_151; // @[ICache.scala 68:{44,44}]
  wire  _GEN_153 = 9'h98 == req_r_addr[13:5] ? valid_152 : _GEN_152; // @[ICache.scala 68:{44,44}]
  wire  _GEN_154 = 9'h99 == req_r_addr[13:5] ? valid_153 : _GEN_153; // @[ICache.scala 68:{44,44}]
  wire  _GEN_155 = 9'h9a == req_r_addr[13:5] ? valid_154 : _GEN_154; // @[ICache.scala 68:{44,44}]
  wire  _GEN_156 = 9'h9b == req_r_addr[13:5] ? valid_155 : _GEN_155; // @[ICache.scala 68:{44,44}]
  wire  _GEN_157 = 9'h9c == req_r_addr[13:5] ? valid_156 : _GEN_156; // @[ICache.scala 68:{44,44}]
  wire  _GEN_158 = 9'h9d == req_r_addr[13:5] ? valid_157 : _GEN_157; // @[ICache.scala 68:{44,44}]
  wire  _GEN_159 = 9'h9e == req_r_addr[13:5] ? valid_158 : _GEN_158; // @[ICache.scala 68:{44,44}]
  wire  _GEN_160 = 9'h9f == req_r_addr[13:5] ? valid_159 : _GEN_159; // @[ICache.scala 68:{44,44}]
  wire  _GEN_161 = 9'ha0 == req_r_addr[13:5] ? valid_160 : _GEN_160; // @[ICache.scala 68:{44,44}]
  wire  _GEN_162 = 9'ha1 == req_r_addr[13:5] ? valid_161 : _GEN_161; // @[ICache.scala 68:{44,44}]
  wire  _GEN_163 = 9'ha2 == req_r_addr[13:5] ? valid_162 : _GEN_162; // @[ICache.scala 68:{44,44}]
  wire  _GEN_164 = 9'ha3 == req_r_addr[13:5] ? valid_163 : _GEN_163; // @[ICache.scala 68:{44,44}]
  wire  _GEN_165 = 9'ha4 == req_r_addr[13:5] ? valid_164 : _GEN_164; // @[ICache.scala 68:{44,44}]
  wire  _GEN_166 = 9'ha5 == req_r_addr[13:5] ? valid_165 : _GEN_165; // @[ICache.scala 68:{44,44}]
  wire  _GEN_167 = 9'ha6 == req_r_addr[13:5] ? valid_166 : _GEN_166; // @[ICache.scala 68:{44,44}]
  wire  _GEN_168 = 9'ha7 == req_r_addr[13:5] ? valid_167 : _GEN_167; // @[ICache.scala 68:{44,44}]
  wire  _GEN_169 = 9'ha8 == req_r_addr[13:5] ? valid_168 : _GEN_168; // @[ICache.scala 68:{44,44}]
  wire  _GEN_170 = 9'ha9 == req_r_addr[13:5] ? valid_169 : _GEN_169; // @[ICache.scala 68:{44,44}]
  wire  _GEN_171 = 9'haa == req_r_addr[13:5] ? valid_170 : _GEN_170; // @[ICache.scala 68:{44,44}]
  wire  _GEN_172 = 9'hab == req_r_addr[13:5] ? valid_171 : _GEN_171; // @[ICache.scala 68:{44,44}]
  wire  _GEN_173 = 9'hac == req_r_addr[13:5] ? valid_172 : _GEN_172; // @[ICache.scala 68:{44,44}]
  wire  _GEN_174 = 9'had == req_r_addr[13:5] ? valid_173 : _GEN_173; // @[ICache.scala 68:{44,44}]
  wire  _GEN_175 = 9'hae == req_r_addr[13:5] ? valid_174 : _GEN_174; // @[ICache.scala 68:{44,44}]
  wire  _GEN_176 = 9'haf == req_r_addr[13:5] ? valid_175 : _GEN_175; // @[ICache.scala 68:{44,44}]
  wire  _GEN_177 = 9'hb0 == req_r_addr[13:5] ? valid_176 : _GEN_176; // @[ICache.scala 68:{44,44}]
  wire  _GEN_178 = 9'hb1 == req_r_addr[13:5] ? valid_177 : _GEN_177; // @[ICache.scala 68:{44,44}]
  wire  _GEN_179 = 9'hb2 == req_r_addr[13:5] ? valid_178 : _GEN_178; // @[ICache.scala 68:{44,44}]
  wire  _GEN_180 = 9'hb3 == req_r_addr[13:5] ? valid_179 : _GEN_179; // @[ICache.scala 68:{44,44}]
  wire  _GEN_181 = 9'hb4 == req_r_addr[13:5] ? valid_180 : _GEN_180; // @[ICache.scala 68:{44,44}]
  wire  _GEN_182 = 9'hb5 == req_r_addr[13:5] ? valid_181 : _GEN_181; // @[ICache.scala 68:{44,44}]
  wire  _GEN_183 = 9'hb6 == req_r_addr[13:5] ? valid_182 : _GEN_182; // @[ICache.scala 68:{44,44}]
  wire  _GEN_184 = 9'hb7 == req_r_addr[13:5] ? valid_183 : _GEN_183; // @[ICache.scala 68:{44,44}]
  wire  _GEN_185 = 9'hb8 == req_r_addr[13:5] ? valid_184 : _GEN_184; // @[ICache.scala 68:{44,44}]
  wire  _GEN_186 = 9'hb9 == req_r_addr[13:5] ? valid_185 : _GEN_185; // @[ICache.scala 68:{44,44}]
  wire  _GEN_187 = 9'hba == req_r_addr[13:5] ? valid_186 : _GEN_186; // @[ICache.scala 68:{44,44}]
  wire  _GEN_188 = 9'hbb == req_r_addr[13:5] ? valid_187 : _GEN_187; // @[ICache.scala 68:{44,44}]
  wire  _GEN_189 = 9'hbc == req_r_addr[13:5] ? valid_188 : _GEN_188; // @[ICache.scala 68:{44,44}]
  wire  _GEN_190 = 9'hbd == req_r_addr[13:5] ? valid_189 : _GEN_189; // @[ICache.scala 68:{44,44}]
  wire  _GEN_191 = 9'hbe == req_r_addr[13:5] ? valid_190 : _GEN_190; // @[ICache.scala 68:{44,44}]
  wire  _GEN_192 = 9'hbf == req_r_addr[13:5] ? valid_191 : _GEN_191; // @[ICache.scala 68:{44,44}]
  wire  _GEN_193 = 9'hc0 == req_r_addr[13:5] ? valid_192 : _GEN_192; // @[ICache.scala 68:{44,44}]
  wire  _GEN_194 = 9'hc1 == req_r_addr[13:5] ? valid_193 : _GEN_193; // @[ICache.scala 68:{44,44}]
  wire  _GEN_195 = 9'hc2 == req_r_addr[13:5] ? valid_194 : _GEN_194; // @[ICache.scala 68:{44,44}]
  wire  _GEN_196 = 9'hc3 == req_r_addr[13:5] ? valid_195 : _GEN_195; // @[ICache.scala 68:{44,44}]
  wire  _GEN_197 = 9'hc4 == req_r_addr[13:5] ? valid_196 : _GEN_196; // @[ICache.scala 68:{44,44}]
  wire  _GEN_198 = 9'hc5 == req_r_addr[13:5] ? valid_197 : _GEN_197; // @[ICache.scala 68:{44,44}]
  wire  _GEN_199 = 9'hc6 == req_r_addr[13:5] ? valid_198 : _GEN_198; // @[ICache.scala 68:{44,44}]
  wire  _GEN_200 = 9'hc7 == req_r_addr[13:5] ? valid_199 : _GEN_199; // @[ICache.scala 68:{44,44}]
  wire  _GEN_201 = 9'hc8 == req_r_addr[13:5] ? valid_200 : _GEN_200; // @[ICache.scala 68:{44,44}]
  wire  _GEN_202 = 9'hc9 == req_r_addr[13:5] ? valid_201 : _GEN_201; // @[ICache.scala 68:{44,44}]
  wire  _GEN_203 = 9'hca == req_r_addr[13:5] ? valid_202 : _GEN_202; // @[ICache.scala 68:{44,44}]
  wire  _GEN_204 = 9'hcb == req_r_addr[13:5] ? valid_203 : _GEN_203; // @[ICache.scala 68:{44,44}]
  wire  _GEN_205 = 9'hcc == req_r_addr[13:5] ? valid_204 : _GEN_204; // @[ICache.scala 68:{44,44}]
  wire  _GEN_206 = 9'hcd == req_r_addr[13:5] ? valid_205 : _GEN_205; // @[ICache.scala 68:{44,44}]
  wire  _GEN_207 = 9'hce == req_r_addr[13:5] ? valid_206 : _GEN_206; // @[ICache.scala 68:{44,44}]
  wire  _GEN_208 = 9'hcf == req_r_addr[13:5] ? valid_207 : _GEN_207; // @[ICache.scala 68:{44,44}]
  wire  _GEN_209 = 9'hd0 == req_r_addr[13:5] ? valid_208 : _GEN_208; // @[ICache.scala 68:{44,44}]
  wire  _GEN_210 = 9'hd1 == req_r_addr[13:5] ? valid_209 : _GEN_209; // @[ICache.scala 68:{44,44}]
  wire  _GEN_211 = 9'hd2 == req_r_addr[13:5] ? valid_210 : _GEN_210; // @[ICache.scala 68:{44,44}]
  wire  _GEN_212 = 9'hd3 == req_r_addr[13:5] ? valid_211 : _GEN_211; // @[ICache.scala 68:{44,44}]
  wire  _GEN_213 = 9'hd4 == req_r_addr[13:5] ? valid_212 : _GEN_212; // @[ICache.scala 68:{44,44}]
  wire  _GEN_214 = 9'hd5 == req_r_addr[13:5] ? valid_213 : _GEN_213; // @[ICache.scala 68:{44,44}]
  wire  _GEN_215 = 9'hd6 == req_r_addr[13:5] ? valid_214 : _GEN_214; // @[ICache.scala 68:{44,44}]
  wire  _GEN_216 = 9'hd7 == req_r_addr[13:5] ? valid_215 : _GEN_215; // @[ICache.scala 68:{44,44}]
  wire  _GEN_217 = 9'hd8 == req_r_addr[13:5] ? valid_216 : _GEN_216; // @[ICache.scala 68:{44,44}]
  wire  _GEN_218 = 9'hd9 == req_r_addr[13:5] ? valid_217 : _GEN_217; // @[ICache.scala 68:{44,44}]
  wire  _GEN_219 = 9'hda == req_r_addr[13:5] ? valid_218 : _GEN_218; // @[ICache.scala 68:{44,44}]
  wire  _GEN_220 = 9'hdb == req_r_addr[13:5] ? valid_219 : _GEN_219; // @[ICache.scala 68:{44,44}]
  wire  _GEN_221 = 9'hdc == req_r_addr[13:5] ? valid_220 : _GEN_220; // @[ICache.scala 68:{44,44}]
  wire  _GEN_222 = 9'hdd == req_r_addr[13:5] ? valid_221 : _GEN_221; // @[ICache.scala 68:{44,44}]
  wire  _GEN_223 = 9'hde == req_r_addr[13:5] ? valid_222 : _GEN_222; // @[ICache.scala 68:{44,44}]
  wire  _GEN_224 = 9'hdf == req_r_addr[13:5] ? valid_223 : _GEN_223; // @[ICache.scala 68:{44,44}]
  wire  _GEN_225 = 9'he0 == req_r_addr[13:5] ? valid_224 : _GEN_224; // @[ICache.scala 68:{44,44}]
  wire  _GEN_226 = 9'he1 == req_r_addr[13:5] ? valid_225 : _GEN_225; // @[ICache.scala 68:{44,44}]
  wire  _GEN_227 = 9'he2 == req_r_addr[13:5] ? valid_226 : _GEN_226; // @[ICache.scala 68:{44,44}]
  wire  _GEN_228 = 9'he3 == req_r_addr[13:5] ? valid_227 : _GEN_227; // @[ICache.scala 68:{44,44}]
  wire  _GEN_229 = 9'he4 == req_r_addr[13:5] ? valid_228 : _GEN_228; // @[ICache.scala 68:{44,44}]
  wire  _GEN_230 = 9'he5 == req_r_addr[13:5] ? valid_229 : _GEN_229; // @[ICache.scala 68:{44,44}]
  wire  _GEN_231 = 9'he6 == req_r_addr[13:5] ? valid_230 : _GEN_230; // @[ICache.scala 68:{44,44}]
  wire  _GEN_232 = 9'he7 == req_r_addr[13:5] ? valid_231 : _GEN_231; // @[ICache.scala 68:{44,44}]
  wire  _GEN_233 = 9'he8 == req_r_addr[13:5] ? valid_232 : _GEN_232; // @[ICache.scala 68:{44,44}]
  wire  _GEN_234 = 9'he9 == req_r_addr[13:5] ? valid_233 : _GEN_233; // @[ICache.scala 68:{44,44}]
  wire  _GEN_235 = 9'hea == req_r_addr[13:5] ? valid_234 : _GEN_234; // @[ICache.scala 68:{44,44}]
  wire  _GEN_236 = 9'heb == req_r_addr[13:5] ? valid_235 : _GEN_235; // @[ICache.scala 68:{44,44}]
  wire  _GEN_237 = 9'hec == req_r_addr[13:5] ? valid_236 : _GEN_236; // @[ICache.scala 68:{44,44}]
  wire  _GEN_238 = 9'hed == req_r_addr[13:5] ? valid_237 : _GEN_237; // @[ICache.scala 68:{44,44}]
  wire  _GEN_239 = 9'hee == req_r_addr[13:5] ? valid_238 : _GEN_238; // @[ICache.scala 68:{44,44}]
  wire  _GEN_240 = 9'hef == req_r_addr[13:5] ? valid_239 : _GEN_239; // @[ICache.scala 68:{44,44}]
  wire  _GEN_241 = 9'hf0 == req_r_addr[13:5] ? valid_240 : _GEN_240; // @[ICache.scala 68:{44,44}]
  wire  _GEN_242 = 9'hf1 == req_r_addr[13:5] ? valid_241 : _GEN_241; // @[ICache.scala 68:{44,44}]
  wire  _GEN_243 = 9'hf2 == req_r_addr[13:5] ? valid_242 : _GEN_242; // @[ICache.scala 68:{44,44}]
  wire  _GEN_244 = 9'hf3 == req_r_addr[13:5] ? valid_243 : _GEN_243; // @[ICache.scala 68:{44,44}]
  wire  _GEN_245 = 9'hf4 == req_r_addr[13:5] ? valid_244 : _GEN_244; // @[ICache.scala 68:{44,44}]
  wire  _GEN_246 = 9'hf5 == req_r_addr[13:5] ? valid_245 : _GEN_245; // @[ICache.scala 68:{44,44}]
  wire  _GEN_247 = 9'hf6 == req_r_addr[13:5] ? valid_246 : _GEN_246; // @[ICache.scala 68:{44,44}]
  wire  _GEN_248 = 9'hf7 == req_r_addr[13:5] ? valid_247 : _GEN_247; // @[ICache.scala 68:{44,44}]
  wire  _GEN_249 = 9'hf8 == req_r_addr[13:5] ? valid_248 : _GEN_248; // @[ICache.scala 68:{44,44}]
  wire  _GEN_250 = 9'hf9 == req_r_addr[13:5] ? valid_249 : _GEN_249; // @[ICache.scala 68:{44,44}]
  wire  _GEN_251 = 9'hfa == req_r_addr[13:5] ? valid_250 : _GEN_250; // @[ICache.scala 68:{44,44}]
  wire  _GEN_252 = 9'hfb == req_r_addr[13:5] ? valid_251 : _GEN_251; // @[ICache.scala 68:{44,44}]
  wire  _GEN_253 = 9'hfc == req_r_addr[13:5] ? valid_252 : _GEN_252; // @[ICache.scala 68:{44,44}]
  wire  _GEN_254 = 9'hfd == req_r_addr[13:5] ? valid_253 : _GEN_253; // @[ICache.scala 68:{44,44}]
  wire  _GEN_255 = 9'hfe == req_r_addr[13:5] ? valid_254 : _GEN_254; // @[ICache.scala 68:{44,44}]
  wire  _GEN_256 = 9'hff == req_r_addr[13:5] ? valid_255 : _GEN_255; // @[ICache.scala 68:{44,44}]
  wire  _GEN_257 = 9'h100 == req_r_addr[13:5] ? valid_256 : _GEN_256; // @[ICache.scala 68:{44,44}]
  wire  _GEN_258 = 9'h101 == req_r_addr[13:5] ? valid_257 : _GEN_257; // @[ICache.scala 68:{44,44}]
  wire  _GEN_259 = 9'h102 == req_r_addr[13:5] ? valid_258 : _GEN_258; // @[ICache.scala 68:{44,44}]
  wire  _GEN_260 = 9'h103 == req_r_addr[13:5] ? valid_259 : _GEN_259; // @[ICache.scala 68:{44,44}]
  wire  _GEN_261 = 9'h104 == req_r_addr[13:5] ? valid_260 : _GEN_260; // @[ICache.scala 68:{44,44}]
  wire  _GEN_262 = 9'h105 == req_r_addr[13:5] ? valid_261 : _GEN_261; // @[ICache.scala 68:{44,44}]
  wire  _GEN_263 = 9'h106 == req_r_addr[13:5] ? valid_262 : _GEN_262; // @[ICache.scala 68:{44,44}]
  wire  _GEN_264 = 9'h107 == req_r_addr[13:5] ? valid_263 : _GEN_263; // @[ICache.scala 68:{44,44}]
  wire  _GEN_265 = 9'h108 == req_r_addr[13:5] ? valid_264 : _GEN_264; // @[ICache.scala 68:{44,44}]
  wire  _GEN_266 = 9'h109 == req_r_addr[13:5] ? valid_265 : _GEN_265; // @[ICache.scala 68:{44,44}]
  wire  _GEN_267 = 9'h10a == req_r_addr[13:5] ? valid_266 : _GEN_266; // @[ICache.scala 68:{44,44}]
  wire  _GEN_268 = 9'h10b == req_r_addr[13:5] ? valid_267 : _GEN_267; // @[ICache.scala 68:{44,44}]
  wire  _GEN_269 = 9'h10c == req_r_addr[13:5] ? valid_268 : _GEN_268; // @[ICache.scala 68:{44,44}]
  wire  _GEN_270 = 9'h10d == req_r_addr[13:5] ? valid_269 : _GEN_269; // @[ICache.scala 68:{44,44}]
  wire  _GEN_271 = 9'h10e == req_r_addr[13:5] ? valid_270 : _GEN_270; // @[ICache.scala 68:{44,44}]
  wire  _GEN_272 = 9'h10f == req_r_addr[13:5] ? valid_271 : _GEN_271; // @[ICache.scala 68:{44,44}]
  wire  _GEN_273 = 9'h110 == req_r_addr[13:5] ? valid_272 : _GEN_272; // @[ICache.scala 68:{44,44}]
  wire  _GEN_274 = 9'h111 == req_r_addr[13:5] ? valid_273 : _GEN_273; // @[ICache.scala 68:{44,44}]
  wire  _GEN_275 = 9'h112 == req_r_addr[13:5] ? valid_274 : _GEN_274; // @[ICache.scala 68:{44,44}]
  wire  _GEN_276 = 9'h113 == req_r_addr[13:5] ? valid_275 : _GEN_275; // @[ICache.scala 68:{44,44}]
  wire  _GEN_277 = 9'h114 == req_r_addr[13:5] ? valid_276 : _GEN_276; // @[ICache.scala 68:{44,44}]
  wire  _GEN_278 = 9'h115 == req_r_addr[13:5] ? valid_277 : _GEN_277; // @[ICache.scala 68:{44,44}]
  wire  _GEN_279 = 9'h116 == req_r_addr[13:5] ? valid_278 : _GEN_278; // @[ICache.scala 68:{44,44}]
  wire  _GEN_280 = 9'h117 == req_r_addr[13:5] ? valid_279 : _GEN_279; // @[ICache.scala 68:{44,44}]
  wire  _GEN_281 = 9'h118 == req_r_addr[13:5] ? valid_280 : _GEN_280; // @[ICache.scala 68:{44,44}]
  wire  _GEN_282 = 9'h119 == req_r_addr[13:5] ? valid_281 : _GEN_281; // @[ICache.scala 68:{44,44}]
  wire  _GEN_283 = 9'h11a == req_r_addr[13:5] ? valid_282 : _GEN_282; // @[ICache.scala 68:{44,44}]
  wire  _GEN_284 = 9'h11b == req_r_addr[13:5] ? valid_283 : _GEN_283; // @[ICache.scala 68:{44,44}]
  wire  _GEN_285 = 9'h11c == req_r_addr[13:5] ? valid_284 : _GEN_284; // @[ICache.scala 68:{44,44}]
  wire  _GEN_286 = 9'h11d == req_r_addr[13:5] ? valid_285 : _GEN_285; // @[ICache.scala 68:{44,44}]
  wire  _GEN_287 = 9'h11e == req_r_addr[13:5] ? valid_286 : _GEN_286; // @[ICache.scala 68:{44,44}]
  wire  _GEN_288 = 9'h11f == req_r_addr[13:5] ? valid_287 : _GEN_287; // @[ICache.scala 68:{44,44}]
  wire  _GEN_289 = 9'h120 == req_r_addr[13:5] ? valid_288 : _GEN_288; // @[ICache.scala 68:{44,44}]
  wire  _GEN_290 = 9'h121 == req_r_addr[13:5] ? valid_289 : _GEN_289; // @[ICache.scala 68:{44,44}]
  wire  _GEN_291 = 9'h122 == req_r_addr[13:5] ? valid_290 : _GEN_290; // @[ICache.scala 68:{44,44}]
  wire  _GEN_292 = 9'h123 == req_r_addr[13:5] ? valid_291 : _GEN_291; // @[ICache.scala 68:{44,44}]
  wire  _GEN_293 = 9'h124 == req_r_addr[13:5] ? valid_292 : _GEN_292; // @[ICache.scala 68:{44,44}]
  wire  _GEN_294 = 9'h125 == req_r_addr[13:5] ? valid_293 : _GEN_293; // @[ICache.scala 68:{44,44}]
  wire  _GEN_295 = 9'h126 == req_r_addr[13:5] ? valid_294 : _GEN_294; // @[ICache.scala 68:{44,44}]
  wire  _GEN_296 = 9'h127 == req_r_addr[13:5] ? valid_295 : _GEN_295; // @[ICache.scala 68:{44,44}]
  wire  _GEN_297 = 9'h128 == req_r_addr[13:5] ? valid_296 : _GEN_296; // @[ICache.scala 68:{44,44}]
  wire  _GEN_298 = 9'h129 == req_r_addr[13:5] ? valid_297 : _GEN_297; // @[ICache.scala 68:{44,44}]
  wire  _GEN_299 = 9'h12a == req_r_addr[13:5] ? valid_298 : _GEN_298; // @[ICache.scala 68:{44,44}]
  wire  _GEN_300 = 9'h12b == req_r_addr[13:5] ? valid_299 : _GEN_299; // @[ICache.scala 68:{44,44}]
  wire  _GEN_301 = 9'h12c == req_r_addr[13:5] ? valid_300 : _GEN_300; // @[ICache.scala 68:{44,44}]
  wire  _GEN_302 = 9'h12d == req_r_addr[13:5] ? valid_301 : _GEN_301; // @[ICache.scala 68:{44,44}]
  wire  _GEN_303 = 9'h12e == req_r_addr[13:5] ? valid_302 : _GEN_302; // @[ICache.scala 68:{44,44}]
  wire  _GEN_304 = 9'h12f == req_r_addr[13:5] ? valid_303 : _GEN_303; // @[ICache.scala 68:{44,44}]
  wire  _GEN_305 = 9'h130 == req_r_addr[13:5] ? valid_304 : _GEN_304; // @[ICache.scala 68:{44,44}]
  wire  _GEN_306 = 9'h131 == req_r_addr[13:5] ? valid_305 : _GEN_305; // @[ICache.scala 68:{44,44}]
  wire  _GEN_307 = 9'h132 == req_r_addr[13:5] ? valid_306 : _GEN_306; // @[ICache.scala 68:{44,44}]
  wire  _GEN_308 = 9'h133 == req_r_addr[13:5] ? valid_307 : _GEN_307; // @[ICache.scala 68:{44,44}]
  wire  _GEN_309 = 9'h134 == req_r_addr[13:5] ? valid_308 : _GEN_308; // @[ICache.scala 68:{44,44}]
  wire  _GEN_310 = 9'h135 == req_r_addr[13:5] ? valid_309 : _GEN_309; // @[ICache.scala 68:{44,44}]
  wire  _GEN_311 = 9'h136 == req_r_addr[13:5] ? valid_310 : _GEN_310; // @[ICache.scala 68:{44,44}]
  wire  _GEN_312 = 9'h137 == req_r_addr[13:5] ? valid_311 : _GEN_311; // @[ICache.scala 68:{44,44}]
  wire  _GEN_313 = 9'h138 == req_r_addr[13:5] ? valid_312 : _GEN_312; // @[ICache.scala 68:{44,44}]
  wire  _GEN_314 = 9'h139 == req_r_addr[13:5] ? valid_313 : _GEN_313; // @[ICache.scala 68:{44,44}]
  wire  _GEN_315 = 9'h13a == req_r_addr[13:5] ? valid_314 : _GEN_314; // @[ICache.scala 68:{44,44}]
  wire  _GEN_316 = 9'h13b == req_r_addr[13:5] ? valid_315 : _GEN_315; // @[ICache.scala 68:{44,44}]
  wire  _GEN_317 = 9'h13c == req_r_addr[13:5] ? valid_316 : _GEN_316; // @[ICache.scala 68:{44,44}]
  wire  _GEN_318 = 9'h13d == req_r_addr[13:5] ? valid_317 : _GEN_317; // @[ICache.scala 68:{44,44}]
  wire  _GEN_319 = 9'h13e == req_r_addr[13:5] ? valid_318 : _GEN_318; // @[ICache.scala 68:{44,44}]
  wire  _GEN_320 = 9'h13f == req_r_addr[13:5] ? valid_319 : _GEN_319; // @[ICache.scala 68:{44,44}]
  wire  _GEN_321 = 9'h140 == req_r_addr[13:5] ? valid_320 : _GEN_320; // @[ICache.scala 68:{44,44}]
  wire  _GEN_322 = 9'h141 == req_r_addr[13:5] ? valid_321 : _GEN_321; // @[ICache.scala 68:{44,44}]
  wire  _GEN_323 = 9'h142 == req_r_addr[13:5] ? valid_322 : _GEN_322; // @[ICache.scala 68:{44,44}]
  wire  _GEN_324 = 9'h143 == req_r_addr[13:5] ? valid_323 : _GEN_323; // @[ICache.scala 68:{44,44}]
  wire  _GEN_325 = 9'h144 == req_r_addr[13:5] ? valid_324 : _GEN_324; // @[ICache.scala 68:{44,44}]
  wire  _GEN_326 = 9'h145 == req_r_addr[13:5] ? valid_325 : _GEN_325; // @[ICache.scala 68:{44,44}]
  wire  _GEN_327 = 9'h146 == req_r_addr[13:5] ? valid_326 : _GEN_326; // @[ICache.scala 68:{44,44}]
  wire  _GEN_328 = 9'h147 == req_r_addr[13:5] ? valid_327 : _GEN_327; // @[ICache.scala 68:{44,44}]
  wire  _GEN_329 = 9'h148 == req_r_addr[13:5] ? valid_328 : _GEN_328; // @[ICache.scala 68:{44,44}]
  wire  _GEN_330 = 9'h149 == req_r_addr[13:5] ? valid_329 : _GEN_329; // @[ICache.scala 68:{44,44}]
  wire  _GEN_331 = 9'h14a == req_r_addr[13:5] ? valid_330 : _GEN_330; // @[ICache.scala 68:{44,44}]
  wire  _GEN_332 = 9'h14b == req_r_addr[13:5] ? valid_331 : _GEN_331; // @[ICache.scala 68:{44,44}]
  wire  _GEN_333 = 9'h14c == req_r_addr[13:5] ? valid_332 : _GEN_332; // @[ICache.scala 68:{44,44}]
  wire  _GEN_334 = 9'h14d == req_r_addr[13:5] ? valid_333 : _GEN_333; // @[ICache.scala 68:{44,44}]
  wire  _GEN_335 = 9'h14e == req_r_addr[13:5] ? valid_334 : _GEN_334; // @[ICache.scala 68:{44,44}]
  wire  _GEN_336 = 9'h14f == req_r_addr[13:5] ? valid_335 : _GEN_335; // @[ICache.scala 68:{44,44}]
  wire  _GEN_337 = 9'h150 == req_r_addr[13:5] ? valid_336 : _GEN_336; // @[ICache.scala 68:{44,44}]
  wire  _GEN_338 = 9'h151 == req_r_addr[13:5] ? valid_337 : _GEN_337; // @[ICache.scala 68:{44,44}]
  wire  _GEN_339 = 9'h152 == req_r_addr[13:5] ? valid_338 : _GEN_338; // @[ICache.scala 68:{44,44}]
  wire  _GEN_340 = 9'h153 == req_r_addr[13:5] ? valid_339 : _GEN_339; // @[ICache.scala 68:{44,44}]
  wire  _GEN_341 = 9'h154 == req_r_addr[13:5] ? valid_340 : _GEN_340; // @[ICache.scala 68:{44,44}]
  wire  _GEN_342 = 9'h155 == req_r_addr[13:5] ? valid_341 : _GEN_341; // @[ICache.scala 68:{44,44}]
  wire  _GEN_343 = 9'h156 == req_r_addr[13:5] ? valid_342 : _GEN_342; // @[ICache.scala 68:{44,44}]
  wire  _GEN_344 = 9'h157 == req_r_addr[13:5] ? valid_343 : _GEN_343; // @[ICache.scala 68:{44,44}]
  wire  _GEN_345 = 9'h158 == req_r_addr[13:5] ? valid_344 : _GEN_344; // @[ICache.scala 68:{44,44}]
  wire  _GEN_346 = 9'h159 == req_r_addr[13:5] ? valid_345 : _GEN_345; // @[ICache.scala 68:{44,44}]
  wire  _GEN_347 = 9'h15a == req_r_addr[13:5] ? valid_346 : _GEN_346; // @[ICache.scala 68:{44,44}]
  wire  _GEN_348 = 9'h15b == req_r_addr[13:5] ? valid_347 : _GEN_347; // @[ICache.scala 68:{44,44}]
  wire  _GEN_349 = 9'h15c == req_r_addr[13:5] ? valid_348 : _GEN_348; // @[ICache.scala 68:{44,44}]
  wire  _GEN_350 = 9'h15d == req_r_addr[13:5] ? valid_349 : _GEN_349; // @[ICache.scala 68:{44,44}]
  wire  _GEN_351 = 9'h15e == req_r_addr[13:5] ? valid_350 : _GEN_350; // @[ICache.scala 68:{44,44}]
  wire  _GEN_352 = 9'h15f == req_r_addr[13:5] ? valid_351 : _GEN_351; // @[ICache.scala 68:{44,44}]
  wire  _GEN_353 = 9'h160 == req_r_addr[13:5] ? valid_352 : _GEN_352; // @[ICache.scala 68:{44,44}]
  wire  _GEN_354 = 9'h161 == req_r_addr[13:5] ? valid_353 : _GEN_353; // @[ICache.scala 68:{44,44}]
  wire  _GEN_355 = 9'h162 == req_r_addr[13:5] ? valid_354 : _GEN_354; // @[ICache.scala 68:{44,44}]
  wire  _GEN_356 = 9'h163 == req_r_addr[13:5] ? valid_355 : _GEN_355; // @[ICache.scala 68:{44,44}]
  wire  _GEN_357 = 9'h164 == req_r_addr[13:5] ? valid_356 : _GEN_356; // @[ICache.scala 68:{44,44}]
  wire  _GEN_358 = 9'h165 == req_r_addr[13:5] ? valid_357 : _GEN_357; // @[ICache.scala 68:{44,44}]
  wire  _GEN_359 = 9'h166 == req_r_addr[13:5] ? valid_358 : _GEN_358; // @[ICache.scala 68:{44,44}]
  wire  _GEN_360 = 9'h167 == req_r_addr[13:5] ? valid_359 : _GEN_359; // @[ICache.scala 68:{44,44}]
  wire  _GEN_361 = 9'h168 == req_r_addr[13:5] ? valid_360 : _GEN_360; // @[ICache.scala 68:{44,44}]
  wire  _GEN_362 = 9'h169 == req_r_addr[13:5] ? valid_361 : _GEN_361; // @[ICache.scala 68:{44,44}]
  wire  _GEN_363 = 9'h16a == req_r_addr[13:5] ? valid_362 : _GEN_362; // @[ICache.scala 68:{44,44}]
  wire  _GEN_364 = 9'h16b == req_r_addr[13:5] ? valid_363 : _GEN_363; // @[ICache.scala 68:{44,44}]
  wire  _GEN_365 = 9'h16c == req_r_addr[13:5] ? valid_364 : _GEN_364; // @[ICache.scala 68:{44,44}]
  wire  _GEN_366 = 9'h16d == req_r_addr[13:5] ? valid_365 : _GEN_365; // @[ICache.scala 68:{44,44}]
  wire  _GEN_367 = 9'h16e == req_r_addr[13:5] ? valid_366 : _GEN_366; // @[ICache.scala 68:{44,44}]
  wire  _GEN_368 = 9'h16f == req_r_addr[13:5] ? valid_367 : _GEN_367; // @[ICache.scala 68:{44,44}]
  wire  _GEN_369 = 9'h170 == req_r_addr[13:5] ? valid_368 : _GEN_368; // @[ICache.scala 68:{44,44}]
  wire  _GEN_370 = 9'h171 == req_r_addr[13:5] ? valid_369 : _GEN_369; // @[ICache.scala 68:{44,44}]
  wire  _GEN_371 = 9'h172 == req_r_addr[13:5] ? valid_370 : _GEN_370; // @[ICache.scala 68:{44,44}]
  wire  _GEN_372 = 9'h173 == req_r_addr[13:5] ? valid_371 : _GEN_371; // @[ICache.scala 68:{44,44}]
  wire  _GEN_373 = 9'h174 == req_r_addr[13:5] ? valid_372 : _GEN_372; // @[ICache.scala 68:{44,44}]
  wire  _GEN_374 = 9'h175 == req_r_addr[13:5] ? valid_373 : _GEN_373; // @[ICache.scala 68:{44,44}]
  wire  _GEN_375 = 9'h176 == req_r_addr[13:5] ? valid_374 : _GEN_374; // @[ICache.scala 68:{44,44}]
  wire  _GEN_376 = 9'h177 == req_r_addr[13:5] ? valid_375 : _GEN_375; // @[ICache.scala 68:{44,44}]
  wire  _GEN_377 = 9'h178 == req_r_addr[13:5] ? valid_376 : _GEN_376; // @[ICache.scala 68:{44,44}]
  wire  _GEN_378 = 9'h179 == req_r_addr[13:5] ? valid_377 : _GEN_377; // @[ICache.scala 68:{44,44}]
  wire  _GEN_379 = 9'h17a == req_r_addr[13:5] ? valid_378 : _GEN_378; // @[ICache.scala 68:{44,44}]
  wire  _GEN_380 = 9'h17b == req_r_addr[13:5] ? valid_379 : _GEN_379; // @[ICache.scala 68:{44,44}]
  wire  _GEN_381 = 9'h17c == req_r_addr[13:5] ? valid_380 : _GEN_380; // @[ICache.scala 68:{44,44}]
  wire  _GEN_382 = 9'h17d == req_r_addr[13:5] ? valid_381 : _GEN_381; // @[ICache.scala 68:{44,44}]
  wire  _GEN_383 = 9'h17e == req_r_addr[13:5] ? valid_382 : _GEN_382; // @[ICache.scala 68:{44,44}]
  wire  _GEN_384 = 9'h17f == req_r_addr[13:5] ? valid_383 : _GEN_383; // @[ICache.scala 68:{44,44}]
  wire  _GEN_385 = 9'h180 == req_r_addr[13:5] ? valid_384 : _GEN_384; // @[ICache.scala 68:{44,44}]
  wire  _GEN_386 = 9'h181 == req_r_addr[13:5] ? valid_385 : _GEN_385; // @[ICache.scala 68:{44,44}]
  wire  _GEN_387 = 9'h182 == req_r_addr[13:5] ? valid_386 : _GEN_386; // @[ICache.scala 68:{44,44}]
  wire  _GEN_388 = 9'h183 == req_r_addr[13:5] ? valid_387 : _GEN_387; // @[ICache.scala 68:{44,44}]
  wire  _GEN_389 = 9'h184 == req_r_addr[13:5] ? valid_388 : _GEN_388; // @[ICache.scala 68:{44,44}]
  wire  _GEN_390 = 9'h185 == req_r_addr[13:5] ? valid_389 : _GEN_389; // @[ICache.scala 68:{44,44}]
  wire  _GEN_391 = 9'h186 == req_r_addr[13:5] ? valid_390 : _GEN_390; // @[ICache.scala 68:{44,44}]
  wire  _GEN_392 = 9'h187 == req_r_addr[13:5] ? valid_391 : _GEN_391; // @[ICache.scala 68:{44,44}]
  wire  _GEN_393 = 9'h188 == req_r_addr[13:5] ? valid_392 : _GEN_392; // @[ICache.scala 68:{44,44}]
  wire  _GEN_394 = 9'h189 == req_r_addr[13:5] ? valid_393 : _GEN_393; // @[ICache.scala 68:{44,44}]
  wire  _GEN_395 = 9'h18a == req_r_addr[13:5] ? valid_394 : _GEN_394; // @[ICache.scala 68:{44,44}]
  wire  _GEN_396 = 9'h18b == req_r_addr[13:5] ? valid_395 : _GEN_395; // @[ICache.scala 68:{44,44}]
  wire  _GEN_397 = 9'h18c == req_r_addr[13:5] ? valid_396 : _GEN_396; // @[ICache.scala 68:{44,44}]
  wire  _GEN_398 = 9'h18d == req_r_addr[13:5] ? valid_397 : _GEN_397; // @[ICache.scala 68:{44,44}]
  wire  _GEN_399 = 9'h18e == req_r_addr[13:5] ? valid_398 : _GEN_398; // @[ICache.scala 68:{44,44}]
  wire  _GEN_400 = 9'h18f == req_r_addr[13:5] ? valid_399 : _GEN_399; // @[ICache.scala 68:{44,44}]
  wire  _GEN_401 = 9'h190 == req_r_addr[13:5] ? valid_400 : _GEN_400; // @[ICache.scala 68:{44,44}]
  wire  _GEN_402 = 9'h191 == req_r_addr[13:5] ? valid_401 : _GEN_401; // @[ICache.scala 68:{44,44}]
  wire  _GEN_403 = 9'h192 == req_r_addr[13:5] ? valid_402 : _GEN_402; // @[ICache.scala 68:{44,44}]
  wire  _GEN_404 = 9'h193 == req_r_addr[13:5] ? valid_403 : _GEN_403; // @[ICache.scala 68:{44,44}]
  wire  _GEN_405 = 9'h194 == req_r_addr[13:5] ? valid_404 : _GEN_404; // @[ICache.scala 68:{44,44}]
  wire  _GEN_406 = 9'h195 == req_r_addr[13:5] ? valid_405 : _GEN_405; // @[ICache.scala 68:{44,44}]
  wire  _GEN_407 = 9'h196 == req_r_addr[13:5] ? valid_406 : _GEN_406; // @[ICache.scala 68:{44,44}]
  wire  _GEN_408 = 9'h197 == req_r_addr[13:5] ? valid_407 : _GEN_407; // @[ICache.scala 68:{44,44}]
  wire  _GEN_409 = 9'h198 == req_r_addr[13:5] ? valid_408 : _GEN_408; // @[ICache.scala 68:{44,44}]
  wire  _GEN_410 = 9'h199 == req_r_addr[13:5] ? valid_409 : _GEN_409; // @[ICache.scala 68:{44,44}]
  wire  _GEN_411 = 9'h19a == req_r_addr[13:5] ? valid_410 : _GEN_410; // @[ICache.scala 68:{44,44}]
  wire  _GEN_412 = 9'h19b == req_r_addr[13:5] ? valid_411 : _GEN_411; // @[ICache.scala 68:{44,44}]
  wire  _GEN_413 = 9'h19c == req_r_addr[13:5] ? valid_412 : _GEN_412; // @[ICache.scala 68:{44,44}]
  wire  _GEN_414 = 9'h19d == req_r_addr[13:5] ? valid_413 : _GEN_413; // @[ICache.scala 68:{44,44}]
  wire  _GEN_415 = 9'h19e == req_r_addr[13:5] ? valid_414 : _GEN_414; // @[ICache.scala 68:{44,44}]
  wire  _GEN_416 = 9'h19f == req_r_addr[13:5] ? valid_415 : _GEN_415; // @[ICache.scala 68:{44,44}]
  wire  _GEN_417 = 9'h1a0 == req_r_addr[13:5] ? valid_416 : _GEN_416; // @[ICache.scala 68:{44,44}]
  wire  _GEN_418 = 9'h1a1 == req_r_addr[13:5] ? valid_417 : _GEN_417; // @[ICache.scala 68:{44,44}]
  wire  _GEN_419 = 9'h1a2 == req_r_addr[13:5] ? valid_418 : _GEN_418; // @[ICache.scala 68:{44,44}]
  wire  _GEN_420 = 9'h1a3 == req_r_addr[13:5] ? valid_419 : _GEN_419; // @[ICache.scala 68:{44,44}]
  wire  _GEN_421 = 9'h1a4 == req_r_addr[13:5] ? valid_420 : _GEN_420; // @[ICache.scala 68:{44,44}]
  wire  _GEN_422 = 9'h1a5 == req_r_addr[13:5] ? valid_421 : _GEN_421; // @[ICache.scala 68:{44,44}]
  wire  _GEN_423 = 9'h1a6 == req_r_addr[13:5] ? valid_422 : _GEN_422; // @[ICache.scala 68:{44,44}]
  wire  _GEN_424 = 9'h1a7 == req_r_addr[13:5] ? valid_423 : _GEN_423; // @[ICache.scala 68:{44,44}]
  wire  _GEN_425 = 9'h1a8 == req_r_addr[13:5] ? valid_424 : _GEN_424; // @[ICache.scala 68:{44,44}]
  wire  _GEN_426 = 9'h1a9 == req_r_addr[13:5] ? valid_425 : _GEN_425; // @[ICache.scala 68:{44,44}]
  wire  _GEN_427 = 9'h1aa == req_r_addr[13:5] ? valid_426 : _GEN_426; // @[ICache.scala 68:{44,44}]
  wire  _GEN_428 = 9'h1ab == req_r_addr[13:5] ? valid_427 : _GEN_427; // @[ICache.scala 68:{44,44}]
  wire  _GEN_429 = 9'h1ac == req_r_addr[13:5] ? valid_428 : _GEN_428; // @[ICache.scala 68:{44,44}]
  wire  _GEN_430 = 9'h1ad == req_r_addr[13:5] ? valid_429 : _GEN_429; // @[ICache.scala 68:{44,44}]
  wire  _GEN_431 = 9'h1ae == req_r_addr[13:5] ? valid_430 : _GEN_430; // @[ICache.scala 68:{44,44}]
  wire  _GEN_432 = 9'h1af == req_r_addr[13:5] ? valid_431 : _GEN_431; // @[ICache.scala 68:{44,44}]
  wire  _GEN_433 = 9'h1b0 == req_r_addr[13:5] ? valid_432 : _GEN_432; // @[ICache.scala 68:{44,44}]
  wire  _GEN_434 = 9'h1b1 == req_r_addr[13:5] ? valid_433 : _GEN_433; // @[ICache.scala 68:{44,44}]
  wire  _GEN_435 = 9'h1b2 == req_r_addr[13:5] ? valid_434 : _GEN_434; // @[ICache.scala 68:{44,44}]
  wire  _GEN_436 = 9'h1b3 == req_r_addr[13:5] ? valid_435 : _GEN_435; // @[ICache.scala 68:{44,44}]
  wire  _GEN_437 = 9'h1b4 == req_r_addr[13:5] ? valid_436 : _GEN_436; // @[ICache.scala 68:{44,44}]
  wire  _GEN_438 = 9'h1b5 == req_r_addr[13:5] ? valid_437 : _GEN_437; // @[ICache.scala 68:{44,44}]
  wire  _GEN_439 = 9'h1b6 == req_r_addr[13:5] ? valid_438 : _GEN_438; // @[ICache.scala 68:{44,44}]
  wire  _GEN_440 = 9'h1b7 == req_r_addr[13:5] ? valid_439 : _GEN_439; // @[ICache.scala 68:{44,44}]
  wire  _GEN_441 = 9'h1b8 == req_r_addr[13:5] ? valid_440 : _GEN_440; // @[ICache.scala 68:{44,44}]
  wire  _GEN_442 = 9'h1b9 == req_r_addr[13:5] ? valid_441 : _GEN_441; // @[ICache.scala 68:{44,44}]
  wire  _GEN_443 = 9'h1ba == req_r_addr[13:5] ? valid_442 : _GEN_442; // @[ICache.scala 68:{44,44}]
  wire  _GEN_444 = 9'h1bb == req_r_addr[13:5] ? valid_443 : _GEN_443; // @[ICache.scala 68:{44,44}]
  wire  _GEN_445 = 9'h1bc == req_r_addr[13:5] ? valid_444 : _GEN_444; // @[ICache.scala 68:{44,44}]
  wire  _GEN_446 = 9'h1bd == req_r_addr[13:5] ? valid_445 : _GEN_445; // @[ICache.scala 68:{44,44}]
  wire  _GEN_447 = 9'h1be == req_r_addr[13:5] ? valid_446 : _GEN_446; // @[ICache.scala 68:{44,44}]
  wire  _GEN_448 = 9'h1bf == req_r_addr[13:5] ? valid_447 : _GEN_447; // @[ICache.scala 68:{44,44}]
  wire  _GEN_449 = 9'h1c0 == req_r_addr[13:5] ? valid_448 : _GEN_448; // @[ICache.scala 68:{44,44}]
  wire  _GEN_450 = 9'h1c1 == req_r_addr[13:5] ? valid_449 : _GEN_449; // @[ICache.scala 68:{44,44}]
  wire  _GEN_451 = 9'h1c2 == req_r_addr[13:5] ? valid_450 : _GEN_450; // @[ICache.scala 68:{44,44}]
  wire  _GEN_452 = 9'h1c3 == req_r_addr[13:5] ? valid_451 : _GEN_451; // @[ICache.scala 68:{44,44}]
  wire  _GEN_453 = 9'h1c4 == req_r_addr[13:5] ? valid_452 : _GEN_452; // @[ICache.scala 68:{44,44}]
  wire  _GEN_454 = 9'h1c5 == req_r_addr[13:5] ? valid_453 : _GEN_453; // @[ICache.scala 68:{44,44}]
  wire  _GEN_455 = 9'h1c6 == req_r_addr[13:5] ? valid_454 : _GEN_454; // @[ICache.scala 68:{44,44}]
  wire  _GEN_456 = 9'h1c7 == req_r_addr[13:5] ? valid_455 : _GEN_455; // @[ICache.scala 68:{44,44}]
  wire  _GEN_457 = 9'h1c8 == req_r_addr[13:5] ? valid_456 : _GEN_456; // @[ICache.scala 68:{44,44}]
  wire  _GEN_458 = 9'h1c9 == req_r_addr[13:5] ? valid_457 : _GEN_457; // @[ICache.scala 68:{44,44}]
  wire  _GEN_459 = 9'h1ca == req_r_addr[13:5] ? valid_458 : _GEN_458; // @[ICache.scala 68:{44,44}]
  wire  _GEN_460 = 9'h1cb == req_r_addr[13:5] ? valid_459 : _GEN_459; // @[ICache.scala 68:{44,44}]
  wire  _GEN_461 = 9'h1cc == req_r_addr[13:5] ? valid_460 : _GEN_460; // @[ICache.scala 68:{44,44}]
  wire  _GEN_462 = 9'h1cd == req_r_addr[13:5] ? valid_461 : _GEN_461; // @[ICache.scala 68:{44,44}]
  wire  _GEN_463 = 9'h1ce == req_r_addr[13:5] ? valid_462 : _GEN_462; // @[ICache.scala 68:{44,44}]
  wire  _GEN_464 = 9'h1cf == req_r_addr[13:5] ? valid_463 : _GEN_463; // @[ICache.scala 68:{44,44}]
  wire  _GEN_465 = 9'h1d0 == req_r_addr[13:5] ? valid_464 : _GEN_464; // @[ICache.scala 68:{44,44}]
  wire  _GEN_466 = 9'h1d1 == req_r_addr[13:5] ? valid_465 : _GEN_465; // @[ICache.scala 68:{44,44}]
  wire  _GEN_467 = 9'h1d2 == req_r_addr[13:5] ? valid_466 : _GEN_466; // @[ICache.scala 68:{44,44}]
  wire  _GEN_468 = 9'h1d3 == req_r_addr[13:5] ? valid_467 : _GEN_467; // @[ICache.scala 68:{44,44}]
  wire  _GEN_469 = 9'h1d4 == req_r_addr[13:5] ? valid_468 : _GEN_468; // @[ICache.scala 68:{44,44}]
  wire  _GEN_470 = 9'h1d5 == req_r_addr[13:5] ? valid_469 : _GEN_469; // @[ICache.scala 68:{44,44}]
  wire  _GEN_471 = 9'h1d6 == req_r_addr[13:5] ? valid_470 : _GEN_470; // @[ICache.scala 68:{44,44}]
  wire  _GEN_472 = 9'h1d7 == req_r_addr[13:5] ? valid_471 : _GEN_471; // @[ICache.scala 68:{44,44}]
  wire  _GEN_473 = 9'h1d8 == req_r_addr[13:5] ? valid_472 : _GEN_472; // @[ICache.scala 68:{44,44}]
  wire  _GEN_474 = 9'h1d9 == req_r_addr[13:5] ? valid_473 : _GEN_473; // @[ICache.scala 68:{44,44}]
  wire  _GEN_475 = 9'h1da == req_r_addr[13:5] ? valid_474 : _GEN_474; // @[ICache.scala 68:{44,44}]
  wire  _GEN_476 = 9'h1db == req_r_addr[13:5] ? valid_475 : _GEN_475; // @[ICache.scala 68:{44,44}]
  wire  _GEN_477 = 9'h1dc == req_r_addr[13:5] ? valid_476 : _GEN_476; // @[ICache.scala 68:{44,44}]
  wire  _GEN_478 = 9'h1dd == req_r_addr[13:5] ? valid_477 : _GEN_477; // @[ICache.scala 68:{44,44}]
  wire  _GEN_479 = 9'h1de == req_r_addr[13:5] ? valid_478 : _GEN_478; // @[ICache.scala 68:{44,44}]
  wire  _GEN_480 = 9'h1df == req_r_addr[13:5] ? valid_479 : _GEN_479; // @[ICache.scala 68:{44,44}]
  wire  _GEN_481 = 9'h1e0 == req_r_addr[13:5] ? valid_480 : _GEN_480; // @[ICache.scala 68:{44,44}]
  wire  _GEN_482 = 9'h1e1 == req_r_addr[13:5] ? valid_481 : _GEN_481; // @[ICache.scala 68:{44,44}]
  wire  _GEN_483 = 9'h1e2 == req_r_addr[13:5] ? valid_482 : _GEN_482; // @[ICache.scala 68:{44,44}]
  wire  _GEN_484 = 9'h1e3 == req_r_addr[13:5] ? valid_483 : _GEN_483; // @[ICache.scala 68:{44,44}]
  wire  _GEN_485 = 9'h1e4 == req_r_addr[13:5] ? valid_484 : _GEN_484; // @[ICache.scala 68:{44,44}]
  wire  _GEN_486 = 9'h1e5 == req_r_addr[13:5] ? valid_485 : _GEN_485; // @[ICache.scala 68:{44,44}]
  wire  _GEN_487 = 9'h1e6 == req_r_addr[13:5] ? valid_486 : _GEN_486; // @[ICache.scala 68:{44,44}]
  wire  _GEN_488 = 9'h1e7 == req_r_addr[13:5] ? valid_487 : _GEN_487; // @[ICache.scala 68:{44,44}]
  wire  _GEN_489 = 9'h1e8 == req_r_addr[13:5] ? valid_488 : _GEN_488; // @[ICache.scala 68:{44,44}]
  wire  _GEN_490 = 9'h1e9 == req_r_addr[13:5] ? valid_489 : _GEN_489; // @[ICache.scala 68:{44,44}]
  wire  _GEN_491 = 9'h1ea == req_r_addr[13:5] ? valid_490 : _GEN_490; // @[ICache.scala 68:{44,44}]
  wire  _GEN_492 = 9'h1eb == req_r_addr[13:5] ? valid_491 : _GEN_491; // @[ICache.scala 68:{44,44}]
  wire  _GEN_493 = 9'h1ec == req_r_addr[13:5] ? valid_492 : _GEN_492; // @[ICache.scala 68:{44,44}]
  wire  _GEN_494 = 9'h1ed == req_r_addr[13:5] ? valid_493 : _GEN_493; // @[ICache.scala 68:{44,44}]
  wire  _GEN_495 = 9'h1ee == req_r_addr[13:5] ? valid_494 : _GEN_494; // @[ICache.scala 68:{44,44}]
  wire  _GEN_496 = 9'h1ef == req_r_addr[13:5] ? valid_495 : _GEN_495; // @[ICache.scala 68:{44,44}]
  wire  _GEN_497 = 9'h1f0 == req_r_addr[13:5] ? valid_496 : _GEN_496; // @[ICache.scala 68:{44,44}]
  wire  _GEN_498 = 9'h1f1 == req_r_addr[13:5] ? valid_497 : _GEN_497; // @[ICache.scala 68:{44,44}]
  wire  _GEN_499 = 9'h1f2 == req_r_addr[13:5] ? valid_498 : _GEN_498; // @[ICache.scala 68:{44,44}]
  wire  _GEN_500 = 9'h1f3 == req_r_addr[13:5] ? valid_499 : _GEN_499; // @[ICache.scala 68:{44,44}]
  wire  _GEN_501 = 9'h1f4 == req_r_addr[13:5] ? valid_500 : _GEN_500; // @[ICache.scala 68:{44,44}]
  wire  _GEN_502 = 9'h1f5 == req_r_addr[13:5] ? valid_501 : _GEN_501; // @[ICache.scala 68:{44,44}]
  wire  _GEN_503 = 9'h1f6 == req_r_addr[13:5] ? valid_502 : _GEN_502; // @[ICache.scala 68:{44,44}]
  wire  _GEN_504 = 9'h1f7 == req_r_addr[13:5] ? valid_503 : _GEN_503; // @[ICache.scala 68:{44,44}]
  wire  _GEN_505 = 9'h1f8 == req_r_addr[13:5] ? valid_504 : _GEN_504; // @[ICache.scala 68:{44,44}]
  wire  _GEN_506 = 9'h1f9 == req_r_addr[13:5] ? valid_505 : _GEN_505; // @[ICache.scala 68:{44,44}]
  wire  _GEN_507 = 9'h1fa == req_r_addr[13:5] ? valid_506 : _GEN_506; // @[ICache.scala 68:{44,44}]
  wire  _GEN_508 = 9'h1fb == req_r_addr[13:5] ? valid_507 : _GEN_507; // @[ICache.scala 68:{44,44}]
  wire  _GEN_509 = 9'h1fc == req_r_addr[13:5] ? valid_508 : _GEN_508; // @[ICache.scala 68:{44,44}]
  wire  _GEN_510 = 9'h1fd == req_r_addr[13:5] ? valid_509 : _GEN_509; // @[ICache.scala 68:{44,44}]
  wire  _GEN_511 = 9'h1fe == req_r_addr[13:5] ? valid_510 : _GEN_510; // @[ICache.scala 68:{44,44}]
  wire  _GEN_512 = 9'h1ff == req_r_addr[13:5] ? valid_511 : _GEN_511; // @[ICache.scala 68:{44,44}]
  reg  array_out_REG; // @[ICache.scala 67:50]
  reg [273:0] array_out_r; // @[Reg.scala 35:20]
  wire [273:0] _array_out_T = array_out_REG ? array_io_rdata : array_out_r; // @[Utils.scala 50:8]
  wire [17:0] array_out_tag = _array_out_T[273:256]; // @[ICache.scala 67:66]
  wire  array_hit = _GEN_512 & req_r_addr[31:14] == array_out_tag; // @[ICache.scala 68:44]
  wire  _s2_ready_T_1 = state == 3'h0 & array_hit; // @[ICache.scala 143:35]
  wire  _s2_ready_T_2 = state == 3'h3; // @[ICache.scala 143:59]
  wire  s2_ready = (state == 3'h0 & array_hit | state == 3'h3 | state == 3'h4) & io_cache_resp_ready; // @[ICache.scala 143:92]
  wire  fire = io_cache_req_valid & s2_ready; // @[ICache.scala 56:27]
  wire  tl_d_ready = state == 3'h2; // @[ICache.scala 152:24]
  wire  _array_io_en_T = tl_d_ready & auto_out_d_valid; // @[Decoupled.scala 51:35]
  wire [255:0] array_out_data = _array_out_T[255:0]; // @[ICache.scala 67:66]
  wire [8:0] _GEN_513 = fire ? io_cache_req_bits_addr[13:5] : 9'h0; // @[ICache.scala 71:14 60:18 72:19]
  wire  _state_T = io_cache_resp_ready & io_cache_resp_valid; // @[Decoupled.scala 51:35]
  wire  _state_T_1 = io_cache_req_ready & io_cache_req_valid; // @[Decoupled.scala 51:35]
  wire  _state_T_2 = ~_state_T_1; // @[ICache.scala 82:33]
  wire  tl_a_valid = state == 3'h1; // @[ICache.scala 150:24]
  wire  _T_2 = auto_out_a_ready & tl_a_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_522 = _array_io_en_T ? 3'h3 : state; // @[ICache.scala 90:23 91:15 78:68]
  wire [2:0] _state_T_8 = _state_T_2 ? 3'h4 : 3'h0; // @[ICache.scala 96:21]
  wire [2:0] _GEN_523 = _state_T ? _state_T_8 : state; // @[ICache.scala 95:23 96:15 78:68]
  wire [2:0] _GEN_524 = _state_T_1 ? 3'h0 : state; // @[ICache.scala 100:22 101:15 78:68]
  wire [2:0] _GEN_525 = 3'h4 == state ? _GEN_524 : state; // @[ICache.scala 80:17 78:68]
  wire [2:0] _GEN_526 = 3'h3 == state ? _GEN_523 : _GEN_525; // @[ICache.scala 80:17]
  wire [63:0] _array_data_T_6 = 2'h1 == req_r_addr[4:3] ? array_out_data[127:64] : array_out_data[63:0]; // @[Mux.scala 81:58]
  wire [63:0] _array_data_T_8 = 2'h2 == req_r_addr[4:3] ? array_out_data[191:128] : _array_data_T_6; // @[Mux.scala 81:58]
  wire [63:0] _array_data_T_10 = 2'h3 == req_r_addr[4:3] ? array_out_data[255:192] : _array_data_T_8; // @[Mux.scala 81:58]
  reg  array_data_REG; // @[ICache.scala 118:12]
  reg [63:0] array_data_r; // @[Reg.scala 35:20]
  wire [63:0] _GEN_530 = array_data_REG ? _array_data_T_10 : array_data_r; // @[Reg.scala 36:18 35:20 36:22]
  reg [255:0] wdata; // @[Reg.scala 35:20]
  wire [273:0] _array_io_wdata_T_1 = {req_r_addr[31:14],auto_out_d_bits_data}; // @[Cat.scala 33:92]
  wire  _GEN_532 = 9'h0 == req_r_addr[13:5] | valid_0; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_533 = 9'h1 == req_r_addr[13:5] | valid_1; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_534 = 9'h2 == req_r_addr[13:5] | valid_2; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_535 = 9'h3 == req_r_addr[13:5] | valid_3; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_536 = 9'h4 == req_r_addr[13:5] | valid_4; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_537 = 9'h5 == req_r_addr[13:5] | valid_5; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_538 = 9'h6 == req_r_addr[13:5] | valid_6; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_539 = 9'h7 == req_r_addr[13:5] | valid_7; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_540 = 9'h8 == req_r_addr[13:5] | valid_8; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_541 = 9'h9 == req_r_addr[13:5] | valid_9; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_542 = 9'ha == req_r_addr[13:5] | valid_10; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_543 = 9'hb == req_r_addr[13:5] | valid_11; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_544 = 9'hc == req_r_addr[13:5] | valid_12; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_545 = 9'hd == req_r_addr[13:5] | valid_13; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_546 = 9'he == req_r_addr[13:5] | valid_14; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_547 = 9'hf == req_r_addr[13:5] | valid_15; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_548 = 9'h10 == req_r_addr[13:5] | valid_16; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_549 = 9'h11 == req_r_addr[13:5] | valid_17; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_550 = 9'h12 == req_r_addr[13:5] | valid_18; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_551 = 9'h13 == req_r_addr[13:5] | valid_19; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_552 = 9'h14 == req_r_addr[13:5] | valid_20; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_553 = 9'h15 == req_r_addr[13:5] | valid_21; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_554 = 9'h16 == req_r_addr[13:5] | valid_22; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_555 = 9'h17 == req_r_addr[13:5] | valid_23; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_556 = 9'h18 == req_r_addr[13:5] | valid_24; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_557 = 9'h19 == req_r_addr[13:5] | valid_25; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_558 = 9'h1a == req_r_addr[13:5] | valid_26; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_559 = 9'h1b == req_r_addr[13:5] | valid_27; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_560 = 9'h1c == req_r_addr[13:5] | valid_28; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_561 = 9'h1d == req_r_addr[13:5] | valid_29; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_562 = 9'h1e == req_r_addr[13:5] | valid_30; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_563 = 9'h1f == req_r_addr[13:5] | valid_31; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_564 = 9'h20 == req_r_addr[13:5] | valid_32; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_565 = 9'h21 == req_r_addr[13:5] | valid_33; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_566 = 9'h22 == req_r_addr[13:5] | valid_34; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_567 = 9'h23 == req_r_addr[13:5] | valid_35; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_568 = 9'h24 == req_r_addr[13:5] | valid_36; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_569 = 9'h25 == req_r_addr[13:5] | valid_37; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_570 = 9'h26 == req_r_addr[13:5] | valid_38; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_571 = 9'h27 == req_r_addr[13:5] | valid_39; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_572 = 9'h28 == req_r_addr[13:5] | valid_40; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_573 = 9'h29 == req_r_addr[13:5] | valid_41; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_574 = 9'h2a == req_r_addr[13:5] | valid_42; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_575 = 9'h2b == req_r_addr[13:5] | valid_43; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_576 = 9'h2c == req_r_addr[13:5] | valid_44; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_577 = 9'h2d == req_r_addr[13:5] | valid_45; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_578 = 9'h2e == req_r_addr[13:5] | valid_46; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_579 = 9'h2f == req_r_addr[13:5] | valid_47; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_580 = 9'h30 == req_r_addr[13:5] | valid_48; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_581 = 9'h31 == req_r_addr[13:5] | valid_49; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_582 = 9'h32 == req_r_addr[13:5] | valid_50; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_583 = 9'h33 == req_r_addr[13:5] | valid_51; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_584 = 9'h34 == req_r_addr[13:5] | valid_52; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_585 = 9'h35 == req_r_addr[13:5] | valid_53; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_586 = 9'h36 == req_r_addr[13:5] | valid_54; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_587 = 9'h37 == req_r_addr[13:5] | valid_55; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_588 = 9'h38 == req_r_addr[13:5] | valid_56; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_589 = 9'h39 == req_r_addr[13:5] | valid_57; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_590 = 9'h3a == req_r_addr[13:5] | valid_58; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_591 = 9'h3b == req_r_addr[13:5] | valid_59; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_592 = 9'h3c == req_r_addr[13:5] | valid_60; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_593 = 9'h3d == req_r_addr[13:5] | valid_61; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_594 = 9'h3e == req_r_addr[13:5] | valid_62; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_595 = 9'h3f == req_r_addr[13:5] | valid_63; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_596 = 9'h40 == req_r_addr[13:5] | valid_64; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_597 = 9'h41 == req_r_addr[13:5] | valid_65; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_598 = 9'h42 == req_r_addr[13:5] | valid_66; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_599 = 9'h43 == req_r_addr[13:5] | valid_67; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_600 = 9'h44 == req_r_addr[13:5] | valid_68; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_601 = 9'h45 == req_r_addr[13:5] | valid_69; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_602 = 9'h46 == req_r_addr[13:5] | valid_70; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_603 = 9'h47 == req_r_addr[13:5] | valid_71; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_604 = 9'h48 == req_r_addr[13:5] | valid_72; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_605 = 9'h49 == req_r_addr[13:5] | valid_73; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_606 = 9'h4a == req_r_addr[13:5] | valid_74; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_607 = 9'h4b == req_r_addr[13:5] | valid_75; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_608 = 9'h4c == req_r_addr[13:5] | valid_76; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_609 = 9'h4d == req_r_addr[13:5] | valid_77; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_610 = 9'h4e == req_r_addr[13:5] | valid_78; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_611 = 9'h4f == req_r_addr[13:5] | valid_79; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_612 = 9'h50 == req_r_addr[13:5] | valid_80; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_613 = 9'h51 == req_r_addr[13:5] | valid_81; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_614 = 9'h52 == req_r_addr[13:5] | valid_82; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_615 = 9'h53 == req_r_addr[13:5] | valid_83; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_616 = 9'h54 == req_r_addr[13:5] | valid_84; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_617 = 9'h55 == req_r_addr[13:5] | valid_85; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_618 = 9'h56 == req_r_addr[13:5] | valid_86; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_619 = 9'h57 == req_r_addr[13:5] | valid_87; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_620 = 9'h58 == req_r_addr[13:5] | valid_88; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_621 = 9'h59 == req_r_addr[13:5] | valid_89; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_622 = 9'h5a == req_r_addr[13:5] | valid_90; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_623 = 9'h5b == req_r_addr[13:5] | valid_91; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_624 = 9'h5c == req_r_addr[13:5] | valid_92; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_625 = 9'h5d == req_r_addr[13:5] | valid_93; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_626 = 9'h5e == req_r_addr[13:5] | valid_94; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_627 = 9'h5f == req_r_addr[13:5] | valid_95; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_628 = 9'h60 == req_r_addr[13:5] | valid_96; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_629 = 9'h61 == req_r_addr[13:5] | valid_97; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_630 = 9'h62 == req_r_addr[13:5] | valid_98; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_631 = 9'h63 == req_r_addr[13:5] | valid_99; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_632 = 9'h64 == req_r_addr[13:5] | valid_100; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_633 = 9'h65 == req_r_addr[13:5] | valid_101; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_634 = 9'h66 == req_r_addr[13:5] | valid_102; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_635 = 9'h67 == req_r_addr[13:5] | valid_103; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_636 = 9'h68 == req_r_addr[13:5] | valid_104; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_637 = 9'h69 == req_r_addr[13:5] | valid_105; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_638 = 9'h6a == req_r_addr[13:5] | valid_106; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_639 = 9'h6b == req_r_addr[13:5] | valid_107; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_640 = 9'h6c == req_r_addr[13:5] | valid_108; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_641 = 9'h6d == req_r_addr[13:5] | valid_109; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_642 = 9'h6e == req_r_addr[13:5] | valid_110; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_643 = 9'h6f == req_r_addr[13:5] | valid_111; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_644 = 9'h70 == req_r_addr[13:5] | valid_112; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_645 = 9'h71 == req_r_addr[13:5] | valid_113; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_646 = 9'h72 == req_r_addr[13:5] | valid_114; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_647 = 9'h73 == req_r_addr[13:5] | valid_115; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_648 = 9'h74 == req_r_addr[13:5] | valid_116; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_649 = 9'h75 == req_r_addr[13:5] | valid_117; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_650 = 9'h76 == req_r_addr[13:5] | valid_118; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_651 = 9'h77 == req_r_addr[13:5] | valid_119; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_652 = 9'h78 == req_r_addr[13:5] | valid_120; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_653 = 9'h79 == req_r_addr[13:5] | valid_121; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_654 = 9'h7a == req_r_addr[13:5] | valid_122; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_655 = 9'h7b == req_r_addr[13:5] | valid_123; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_656 = 9'h7c == req_r_addr[13:5] | valid_124; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_657 = 9'h7d == req_r_addr[13:5] | valid_125; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_658 = 9'h7e == req_r_addr[13:5] | valid_126; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_659 = 9'h7f == req_r_addr[13:5] | valid_127; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_660 = 9'h80 == req_r_addr[13:5] | valid_128; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_661 = 9'h81 == req_r_addr[13:5] | valid_129; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_662 = 9'h82 == req_r_addr[13:5] | valid_130; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_663 = 9'h83 == req_r_addr[13:5] | valid_131; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_664 = 9'h84 == req_r_addr[13:5] | valid_132; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_665 = 9'h85 == req_r_addr[13:5] | valid_133; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_666 = 9'h86 == req_r_addr[13:5] | valid_134; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_667 = 9'h87 == req_r_addr[13:5] | valid_135; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_668 = 9'h88 == req_r_addr[13:5] | valid_136; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_669 = 9'h89 == req_r_addr[13:5] | valid_137; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_670 = 9'h8a == req_r_addr[13:5] | valid_138; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_671 = 9'h8b == req_r_addr[13:5] | valid_139; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_672 = 9'h8c == req_r_addr[13:5] | valid_140; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_673 = 9'h8d == req_r_addr[13:5] | valid_141; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_674 = 9'h8e == req_r_addr[13:5] | valid_142; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_675 = 9'h8f == req_r_addr[13:5] | valid_143; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_676 = 9'h90 == req_r_addr[13:5] | valid_144; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_677 = 9'h91 == req_r_addr[13:5] | valid_145; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_678 = 9'h92 == req_r_addr[13:5] | valid_146; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_679 = 9'h93 == req_r_addr[13:5] | valid_147; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_680 = 9'h94 == req_r_addr[13:5] | valid_148; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_681 = 9'h95 == req_r_addr[13:5] | valid_149; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_682 = 9'h96 == req_r_addr[13:5] | valid_150; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_683 = 9'h97 == req_r_addr[13:5] | valid_151; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_684 = 9'h98 == req_r_addr[13:5] | valid_152; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_685 = 9'h99 == req_r_addr[13:5] | valid_153; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_686 = 9'h9a == req_r_addr[13:5] | valid_154; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_687 = 9'h9b == req_r_addr[13:5] | valid_155; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_688 = 9'h9c == req_r_addr[13:5] | valid_156; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_689 = 9'h9d == req_r_addr[13:5] | valid_157; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_690 = 9'h9e == req_r_addr[13:5] | valid_158; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_691 = 9'h9f == req_r_addr[13:5] | valid_159; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_692 = 9'ha0 == req_r_addr[13:5] | valid_160; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_693 = 9'ha1 == req_r_addr[13:5] | valid_161; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_694 = 9'ha2 == req_r_addr[13:5] | valid_162; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_695 = 9'ha3 == req_r_addr[13:5] | valid_163; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_696 = 9'ha4 == req_r_addr[13:5] | valid_164; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_697 = 9'ha5 == req_r_addr[13:5] | valid_165; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_698 = 9'ha6 == req_r_addr[13:5] | valid_166; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_699 = 9'ha7 == req_r_addr[13:5] | valid_167; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_700 = 9'ha8 == req_r_addr[13:5] | valid_168; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_701 = 9'ha9 == req_r_addr[13:5] | valid_169; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_702 = 9'haa == req_r_addr[13:5] | valid_170; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_703 = 9'hab == req_r_addr[13:5] | valid_171; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_704 = 9'hac == req_r_addr[13:5] | valid_172; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_705 = 9'had == req_r_addr[13:5] | valid_173; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_706 = 9'hae == req_r_addr[13:5] | valid_174; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_707 = 9'haf == req_r_addr[13:5] | valid_175; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_708 = 9'hb0 == req_r_addr[13:5] | valid_176; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_709 = 9'hb1 == req_r_addr[13:5] | valid_177; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_710 = 9'hb2 == req_r_addr[13:5] | valid_178; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_711 = 9'hb3 == req_r_addr[13:5] | valid_179; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_712 = 9'hb4 == req_r_addr[13:5] | valid_180; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_713 = 9'hb5 == req_r_addr[13:5] | valid_181; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_714 = 9'hb6 == req_r_addr[13:5] | valid_182; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_715 = 9'hb7 == req_r_addr[13:5] | valid_183; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_716 = 9'hb8 == req_r_addr[13:5] | valid_184; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_717 = 9'hb9 == req_r_addr[13:5] | valid_185; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_718 = 9'hba == req_r_addr[13:5] | valid_186; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_719 = 9'hbb == req_r_addr[13:5] | valid_187; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_720 = 9'hbc == req_r_addr[13:5] | valid_188; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_721 = 9'hbd == req_r_addr[13:5] | valid_189; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_722 = 9'hbe == req_r_addr[13:5] | valid_190; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_723 = 9'hbf == req_r_addr[13:5] | valid_191; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_724 = 9'hc0 == req_r_addr[13:5] | valid_192; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_725 = 9'hc1 == req_r_addr[13:5] | valid_193; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_726 = 9'hc2 == req_r_addr[13:5] | valid_194; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_727 = 9'hc3 == req_r_addr[13:5] | valid_195; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_728 = 9'hc4 == req_r_addr[13:5] | valid_196; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_729 = 9'hc5 == req_r_addr[13:5] | valid_197; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_730 = 9'hc6 == req_r_addr[13:5] | valid_198; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_731 = 9'hc7 == req_r_addr[13:5] | valid_199; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_732 = 9'hc8 == req_r_addr[13:5] | valid_200; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_733 = 9'hc9 == req_r_addr[13:5] | valid_201; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_734 = 9'hca == req_r_addr[13:5] | valid_202; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_735 = 9'hcb == req_r_addr[13:5] | valid_203; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_736 = 9'hcc == req_r_addr[13:5] | valid_204; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_737 = 9'hcd == req_r_addr[13:5] | valid_205; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_738 = 9'hce == req_r_addr[13:5] | valid_206; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_739 = 9'hcf == req_r_addr[13:5] | valid_207; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_740 = 9'hd0 == req_r_addr[13:5] | valid_208; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_741 = 9'hd1 == req_r_addr[13:5] | valid_209; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_742 = 9'hd2 == req_r_addr[13:5] | valid_210; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_743 = 9'hd3 == req_r_addr[13:5] | valid_211; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_744 = 9'hd4 == req_r_addr[13:5] | valid_212; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_745 = 9'hd5 == req_r_addr[13:5] | valid_213; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_746 = 9'hd6 == req_r_addr[13:5] | valid_214; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_747 = 9'hd7 == req_r_addr[13:5] | valid_215; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_748 = 9'hd8 == req_r_addr[13:5] | valid_216; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_749 = 9'hd9 == req_r_addr[13:5] | valid_217; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_750 = 9'hda == req_r_addr[13:5] | valid_218; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_751 = 9'hdb == req_r_addr[13:5] | valid_219; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_752 = 9'hdc == req_r_addr[13:5] | valid_220; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_753 = 9'hdd == req_r_addr[13:5] | valid_221; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_754 = 9'hde == req_r_addr[13:5] | valid_222; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_755 = 9'hdf == req_r_addr[13:5] | valid_223; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_756 = 9'he0 == req_r_addr[13:5] | valid_224; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_757 = 9'he1 == req_r_addr[13:5] | valid_225; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_758 = 9'he2 == req_r_addr[13:5] | valid_226; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_759 = 9'he3 == req_r_addr[13:5] | valid_227; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_760 = 9'he4 == req_r_addr[13:5] | valid_228; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_761 = 9'he5 == req_r_addr[13:5] | valid_229; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_762 = 9'he6 == req_r_addr[13:5] | valid_230; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_763 = 9'he7 == req_r_addr[13:5] | valid_231; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_764 = 9'he8 == req_r_addr[13:5] | valid_232; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_765 = 9'he9 == req_r_addr[13:5] | valid_233; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_766 = 9'hea == req_r_addr[13:5] | valid_234; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_767 = 9'heb == req_r_addr[13:5] | valid_235; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_768 = 9'hec == req_r_addr[13:5] | valid_236; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_769 = 9'hed == req_r_addr[13:5] | valid_237; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_770 = 9'hee == req_r_addr[13:5] | valid_238; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_771 = 9'hef == req_r_addr[13:5] | valid_239; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_772 = 9'hf0 == req_r_addr[13:5] | valid_240; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_773 = 9'hf1 == req_r_addr[13:5] | valid_241; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_774 = 9'hf2 == req_r_addr[13:5] | valid_242; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_775 = 9'hf3 == req_r_addr[13:5] | valid_243; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_776 = 9'hf4 == req_r_addr[13:5] | valid_244; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_777 = 9'hf5 == req_r_addr[13:5] | valid_245; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_778 = 9'hf6 == req_r_addr[13:5] | valid_246; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_779 = 9'hf7 == req_r_addr[13:5] | valid_247; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_780 = 9'hf8 == req_r_addr[13:5] | valid_248; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_781 = 9'hf9 == req_r_addr[13:5] | valid_249; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_782 = 9'hfa == req_r_addr[13:5] | valid_250; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_783 = 9'hfb == req_r_addr[13:5] | valid_251; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_784 = 9'hfc == req_r_addr[13:5] | valid_252; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_785 = 9'hfd == req_r_addr[13:5] | valid_253; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_786 = 9'hfe == req_r_addr[13:5] | valid_254; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_787 = 9'hff == req_r_addr[13:5] | valid_255; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_788 = 9'h100 == req_r_addr[13:5] | valid_256; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_789 = 9'h101 == req_r_addr[13:5] | valid_257; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_790 = 9'h102 == req_r_addr[13:5] | valid_258; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_791 = 9'h103 == req_r_addr[13:5] | valid_259; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_792 = 9'h104 == req_r_addr[13:5] | valid_260; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_793 = 9'h105 == req_r_addr[13:5] | valid_261; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_794 = 9'h106 == req_r_addr[13:5] | valid_262; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_795 = 9'h107 == req_r_addr[13:5] | valid_263; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_796 = 9'h108 == req_r_addr[13:5] | valid_264; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_797 = 9'h109 == req_r_addr[13:5] | valid_265; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_798 = 9'h10a == req_r_addr[13:5] | valid_266; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_799 = 9'h10b == req_r_addr[13:5] | valid_267; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_800 = 9'h10c == req_r_addr[13:5] | valid_268; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_801 = 9'h10d == req_r_addr[13:5] | valid_269; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_802 = 9'h10e == req_r_addr[13:5] | valid_270; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_803 = 9'h10f == req_r_addr[13:5] | valid_271; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_804 = 9'h110 == req_r_addr[13:5] | valid_272; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_805 = 9'h111 == req_r_addr[13:5] | valid_273; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_806 = 9'h112 == req_r_addr[13:5] | valid_274; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_807 = 9'h113 == req_r_addr[13:5] | valid_275; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_808 = 9'h114 == req_r_addr[13:5] | valid_276; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_809 = 9'h115 == req_r_addr[13:5] | valid_277; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_810 = 9'h116 == req_r_addr[13:5] | valid_278; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_811 = 9'h117 == req_r_addr[13:5] | valid_279; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_812 = 9'h118 == req_r_addr[13:5] | valid_280; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_813 = 9'h119 == req_r_addr[13:5] | valid_281; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_814 = 9'h11a == req_r_addr[13:5] | valid_282; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_815 = 9'h11b == req_r_addr[13:5] | valid_283; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_816 = 9'h11c == req_r_addr[13:5] | valid_284; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_817 = 9'h11d == req_r_addr[13:5] | valid_285; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_818 = 9'h11e == req_r_addr[13:5] | valid_286; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_819 = 9'h11f == req_r_addr[13:5] | valid_287; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_820 = 9'h120 == req_r_addr[13:5] | valid_288; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_821 = 9'h121 == req_r_addr[13:5] | valid_289; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_822 = 9'h122 == req_r_addr[13:5] | valid_290; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_823 = 9'h123 == req_r_addr[13:5] | valid_291; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_824 = 9'h124 == req_r_addr[13:5] | valid_292; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_825 = 9'h125 == req_r_addr[13:5] | valid_293; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_826 = 9'h126 == req_r_addr[13:5] | valid_294; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_827 = 9'h127 == req_r_addr[13:5] | valid_295; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_828 = 9'h128 == req_r_addr[13:5] | valid_296; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_829 = 9'h129 == req_r_addr[13:5] | valid_297; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_830 = 9'h12a == req_r_addr[13:5] | valid_298; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_831 = 9'h12b == req_r_addr[13:5] | valid_299; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_832 = 9'h12c == req_r_addr[13:5] | valid_300; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_833 = 9'h12d == req_r_addr[13:5] | valid_301; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_834 = 9'h12e == req_r_addr[13:5] | valid_302; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_835 = 9'h12f == req_r_addr[13:5] | valid_303; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_836 = 9'h130 == req_r_addr[13:5] | valid_304; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_837 = 9'h131 == req_r_addr[13:5] | valid_305; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_838 = 9'h132 == req_r_addr[13:5] | valid_306; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_839 = 9'h133 == req_r_addr[13:5] | valid_307; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_840 = 9'h134 == req_r_addr[13:5] | valid_308; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_841 = 9'h135 == req_r_addr[13:5] | valid_309; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_842 = 9'h136 == req_r_addr[13:5] | valid_310; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_843 = 9'h137 == req_r_addr[13:5] | valid_311; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_844 = 9'h138 == req_r_addr[13:5] | valid_312; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_845 = 9'h139 == req_r_addr[13:5] | valid_313; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_846 = 9'h13a == req_r_addr[13:5] | valid_314; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_847 = 9'h13b == req_r_addr[13:5] | valid_315; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_848 = 9'h13c == req_r_addr[13:5] | valid_316; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_849 = 9'h13d == req_r_addr[13:5] | valid_317; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_850 = 9'h13e == req_r_addr[13:5] | valid_318; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_851 = 9'h13f == req_r_addr[13:5] | valid_319; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_852 = 9'h140 == req_r_addr[13:5] | valid_320; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_853 = 9'h141 == req_r_addr[13:5] | valid_321; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_854 = 9'h142 == req_r_addr[13:5] | valid_322; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_855 = 9'h143 == req_r_addr[13:5] | valid_323; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_856 = 9'h144 == req_r_addr[13:5] | valid_324; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_857 = 9'h145 == req_r_addr[13:5] | valid_325; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_858 = 9'h146 == req_r_addr[13:5] | valid_326; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_859 = 9'h147 == req_r_addr[13:5] | valid_327; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_860 = 9'h148 == req_r_addr[13:5] | valid_328; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_861 = 9'h149 == req_r_addr[13:5] | valid_329; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_862 = 9'h14a == req_r_addr[13:5] | valid_330; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_863 = 9'h14b == req_r_addr[13:5] | valid_331; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_864 = 9'h14c == req_r_addr[13:5] | valid_332; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_865 = 9'h14d == req_r_addr[13:5] | valid_333; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_866 = 9'h14e == req_r_addr[13:5] | valid_334; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_867 = 9'h14f == req_r_addr[13:5] | valid_335; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_868 = 9'h150 == req_r_addr[13:5] | valid_336; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_869 = 9'h151 == req_r_addr[13:5] | valid_337; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_870 = 9'h152 == req_r_addr[13:5] | valid_338; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_871 = 9'h153 == req_r_addr[13:5] | valid_339; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_872 = 9'h154 == req_r_addr[13:5] | valid_340; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_873 = 9'h155 == req_r_addr[13:5] | valid_341; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_874 = 9'h156 == req_r_addr[13:5] | valid_342; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_875 = 9'h157 == req_r_addr[13:5] | valid_343; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_876 = 9'h158 == req_r_addr[13:5] | valid_344; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_877 = 9'h159 == req_r_addr[13:5] | valid_345; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_878 = 9'h15a == req_r_addr[13:5] | valid_346; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_879 = 9'h15b == req_r_addr[13:5] | valid_347; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_880 = 9'h15c == req_r_addr[13:5] | valid_348; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_881 = 9'h15d == req_r_addr[13:5] | valid_349; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_882 = 9'h15e == req_r_addr[13:5] | valid_350; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_883 = 9'h15f == req_r_addr[13:5] | valid_351; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_884 = 9'h160 == req_r_addr[13:5] | valid_352; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_885 = 9'h161 == req_r_addr[13:5] | valid_353; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_886 = 9'h162 == req_r_addr[13:5] | valid_354; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_887 = 9'h163 == req_r_addr[13:5] | valid_355; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_888 = 9'h164 == req_r_addr[13:5] | valid_356; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_889 = 9'h165 == req_r_addr[13:5] | valid_357; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_890 = 9'h166 == req_r_addr[13:5] | valid_358; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_891 = 9'h167 == req_r_addr[13:5] | valid_359; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_892 = 9'h168 == req_r_addr[13:5] | valid_360; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_893 = 9'h169 == req_r_addr[13:5] | valid_361; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_894 = 9'h16a == req_r_addr[13:5] | valid_362; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_895 = 9'h16b == req_r_addr[13:5] | valid_363; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_896 = 9'h16c == req_r_addr[13:5] | valid_364; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_897 = 9'h16d == req_r_addr[13:5] | valid_365; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_898 = 9'h16e == req_r_addr[13:5] | valid_366; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_899 = 9'h16f == req_r_addr[13:5] | valid_367; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_900 = 9'h170 == req_r_addr[13:5] | valid_368; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_901 = 9'h171 == req_r_addr[13:5] | valid_369; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_902 = 9'h172 == req_r_addr[13:5] | valid_370; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_903 = 9'h173 == req_r_addr[13:5] | valid_371; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_904 = 9'h174 == req_r_addr[13:5] | valid_372; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_905 = 9'h175 == req_r_addr[13:5] | valid_373; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_906 = 9'h176 == req_r_addr[13:5] | valid_374; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_907 = 9'h177 == req_r_addr[13:5] | valid_375; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_908 = 9'h178 == req_r_addr[13:5] | valid_376; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_909 = 9'h179 == req_r_addr[13:5] | valid_377; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_910 = 9'h17a == req_r_addr[13:5] | valid_378; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_911 = 9'h17b == req_r_addr[13:5] | valid_379; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_912 = 9'h17c == req_r_addr[13:5] | valid_380; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_913 = 9'h17d == req_r_addr[13:5] | valid_381; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_914 = 9'h17e == req_r_addr[13:5] | valid_382; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_915 = 9'h17f == req_r_addr[13:5] | valid_383; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_916 = 9'h180 == req_r_addr[13:5] | valid_384; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_917 = 9'h181 == req_r_addr[13:5] | valid_385; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_918 = 9'h182 == req_r_addr[13:5] | valid_386; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_919 = 9'h183 == req_r_addr[13:5] | valid_387; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_920 = 9'h184 == req_r_addr[13:5] | valid_388; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_921 = 9'h185 == req_r_addr[13:5] | valid_389; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_922 = 9'h186 == req_r_addr[13:5] | valid_390; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_923 = 9'h187 == req_r_addr[13:5] | valid_391; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_924 = 9'h188 == req_r_addr[13:5] | valid_392; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_925 = 9'h189 == req_r_addr[13:5] | valid_393; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_926 = 9'h18a == req_r_addr[13:5] | valid_394; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_927 = 9'h18b == req_r_addr[13:5] | valid_395; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_928 = 9'h18c == req_r_addr[13:5] | valid_396; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_929 = 9'h18d == req_r_addr[13:5] | valid_397; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_930 = 9'h18e == req_r_addr[13:5] | valid_398; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_931 = 9'h18f == req_r_addr[13:5] | valid_399; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_932 = 9'h190 == req_r_addr[13:5] | valid_400; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_933 = 9'h191 == req_r_addr[13:5] | valid_401; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_934 = 9'h192 == req_r_addr[13:5] | valid_402; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_935 = 9'h193 == req_r_addr[13:5] | valid_403; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_936 = 9'h194 == req_r_addr[13:5] | valid_404; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_937 = 9'h195 == req_r_addr[13:5] | valid_405; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_938 = 9'h196 == req_r_addr[13:5] | valid_406; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_939 = 9'h197 == req_r_addr[13:5] | valid_407; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_940 = 9'h198 == req_r_addr[13:5] | valid_408; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_941 = 9'h199 == req_r_addr[13:5] | valid_409; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_942 = 9'h19a == req_r_addr[13:5] | valid_410; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_943 = 9'h19b == req_r_addr[13:5] | valid_411; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_944 = 9'h19c == req_r_addr[13:5] | valid_412; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_945 = 9'h19d == req_r_addr[13:5] | valid_413; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_946 = 9'h19e == req_r_addr[13:5] | valid_414; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_947 = 9'h19f == req_r_addr[13:5] | valid_415; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_948 = 9'h1a0 == req_r_addr[13:5] | valid_416; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_949 = 9'h1a1 == req_r_addr[13:5] | valid_417; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_950 = 9'h1a2 == req_r_addr[13:5] | valid_418; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_951 = 9'h1a3 == req_r_addr[13:5] | valid_419; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_952 = 9'h1a4 == req_r_addr[13:5] | valid_420; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_953 = 9'h1a5 == req_r_addr[13:5] | valid_421; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_954 = 9'h1a6 == req_r_addr[13:5] | valid_422; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_955 = 9'h1a7 == req_r_addr[13:5] | valid_423; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_956 = 9'h1a8 == req_r_addr[13:5] | valid_424; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_957 = 9'h1a9 == req_r_addr[13:5] | valid_425; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_958 = 9'h1aa == req_r_addr[13:5] | valid_426; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_959 = 9'h1ab == req_r_addr[13:5] | valid_427; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_960 = 9'h1ac == req_r_addr[13:5] | valid_428; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_961 = 9'h1ad == req_r_addr[13:5] | valid_429; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_962 = 9'h1ae == req_r_addr[13:5] | valid_430; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_963 = 9'h1af == req_r_addr[13:5] | valid_431; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_964 = 9'h1b0 == req_r_addr[13:5] | valid_432; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_965 = 9'h1b1 == req_r_addr[13:5] | valid_433; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_966 = 9'h1b2 == req_r_addr[13:5] | valid_434; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_967 = 9'h1b3 == req_r_addr[13:5] | valid_435; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_968 = 9'h1b4 == req_r_addr[13:5] | valid_436; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_969 = 9'h1b5 == req_r_addr[13:5] | valid_437; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_970 = 9'h1b6 == req_r_addr[13:5] | valid_438; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_971 = 9'h1b7 == req_r_addr[13:5] | valid_439; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_972 = 9'h1b8 == req_r_addr[13:5] | valid_440; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_973 = 9'h1b9 == req_r_addr[13:5] | valid_441; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_974 = 9'h1ba == req_r_addr[13:5] | valid_442; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_975 = 9'h1bb == req_r_addr[13:5] | valid_443; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_976 = 9'h1bc == req_r_addr[13:5] | valid_444; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_977 = 9'h1bd == req_r_addr[13:5] | valid_445; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_978 = 9'h1be == req_r_addr[13:5] | valid_446; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_979 = 9'h1bf == req_r_addr[13:5] | valid_447; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_980 = 9'h1c0 == req_r_addr[13:5] | valid_448; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_981 = 9'h1c1 == req_r_addr[13:5] | valid_449; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_982 = 9'h1c2 == req_r_addr[13:5] | valid_450; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_983 = 9'h1c3 == req_r_addr[13:5] | valid_451; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_984 = 9'h1c4 == req_r_addr[13:5] | valid_452; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_985 = 9'h1c5 == req_r_addr[13:5] | valid_453; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_986 = 9'h1c6 == req_r_addr[13:5] | valid_454; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_987 = 9'h1c7 == req_r_addr[13:5] | valid_455; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_988 = 9'h1c8 == req_r_addr[13:5] | valid_456; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_989 = 9'h1c9 == req_r_addr[13:5] | valid_457; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_990 = 9'h1ca == req_r_addr[13:5] | valid_458; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_991 = 9'h1cb == req_r_addr[13:5] | valid_459; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_992 = 9'h1cc == req_r_addr[13:5] | valid_460; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_993 = 9'h1cd == req_r_addr[13:5] | valid_461; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_994 = 9'h1ce == req_r_addr[13:5] | valid_462; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_995 = 9'h1cf == req_r_addr[13:5] | valid_463; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_996 = 9'h1d0 == req_r_addr[13:5] | valid_464; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_997 = 9'h1d1 == req_r_addr[13:5] | valid_465; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_998 = 9'h1d2 == req_r_addr[13:5] | valid_466; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_999 = 9'h1d3 == req_r_addr[13:5] | valid_467; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1000 = 9'h1d4 == req_r_addr[13:5] | valid_468; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1001 = 9'h1d5 == req_r_addr[13:5] | valid_469; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1002 = 9'h1d6 == req_r_addr[13:5] | valid_470; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1003 = 9'h1d7 == req_r_addr[13:5] | valid_471; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1004 = 9'h1d8 == req_r_addr[13:5] | valid_472; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1005 = 9'h1d9 == req_r_addr[13:5] | valid_473; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1006 = 9'h1da == req_r_addr[13:5] | valid_474; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1007 = 9'h1db == req_r_addr[13:5] | valid_475; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1008 = 9'h1dc == req_r_addr[13:5] | valid_476; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1009 = 9'h1dd == req_r_addr[13:5] | valid_477; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1010 = 9'h1de == req_r_addr[13:5] | valid_478; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1011 = 9'h1df == req_r_addr[13:5] | valid_479; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1012 = 9'h1e0 == req_r_addr[13:5] | valid_480; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1013 = 9'h1e1 == req_r_addr[13:5] | valid_481; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1014 = 9'h1e2 == req_r_addr[13:5] | valid_482; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1015 = 9'h1e3 == req_r_addr[13:5] | valid_483; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1016 = 9'h1e4 == req_r_addr[13:5] | valid_484; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1017 = 9'h1e5 == req_r_addr[13:5] | valid_485; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1018 = 9'h1e6 == req_r_addr[13:5] | valid_486; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1019 = 9'h1e7 == req_r_addr[13:5] | valid_487; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1020 = 9'h1e8 == req_r_addr[13:5] | valid_488; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1021 = 9'h1e9 == req_r_addr[13:5] | valid_489; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1022 = 9'h1ea == req_r_addr[13:5] | valid_490; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1023 = 9'h1eb == req_r_addr[13:5] | valid_491; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1024 = 9'h1ec == req_r_addr[13:5] | valid_492; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1025 = 9'h1ed == req_r_addr[13:5] | valid_493; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1026 = 9'h1ee == req_r_addr[13:5] | valid_494; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1027 = 9'h1ef == req_r_addr[13:5] | valid_495; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1028 = 9'h1f0 == req_r_addr[13:5] | valid_496; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1029 = 9'h1f1 == req_r_addr[13:5] | valid_497; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1030 = 9'h1f2 == req_r_addr[13:5] | valid_498; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1031 = 9'h1f3 == req_r_addr[13:5] | valid_499; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1032 = 9'h1f4 == req_r_addr[13:5] | valid_500; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1033 = 9'h1f5 == req_r_addr[13:5] | valid_501; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1034 = 9'h1f6 == req_r_addr[13:5] | valid_502; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1035 = 9'h1f7 == req_r_addr[13:5] | valid_503; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1036 = 9'h1f8 == req_r_addr[13:5] | valid_504; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1037 = 9'h1f9 == req_r_addr[13:5] | valid_505; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1038 = 9'h1fa == req_r_addr[13:5] | valid_506; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1039 = 9'h1fb == req_r_addr[13:5] | valid_507; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1040 = 9'h1fc == req_r_addr[13:5] | valid_508; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1041 = 9'h1fd == req_r_addr[13:5] | valid_509; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1042 = 9'h1fe == req_r_addr[13:5] | valid_510; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1043 = 9'h1ff == req_r_addr[13:5] | valid_511; // @[ICache.scala 128:{33,33} 51:22]
  wire [63:0] _refill_data_T_6 = 2'h1 == req_r_addr[4:3] ? wdata[127:64] : wdata[63:0]; // @[Mux.scala 81:58]
  wire [63:0] _refill_data_T_8 = 2'h2 == req_r_addr[4:3] ? wdata[191:128] : _refill_data_T_6; // @[Mux.scala 81:58]
  wire [63:0] refill_data = 2'h3 == req_r_addr[4:3] ? wdata[255:192] : _refill_data_T_8; // @[Mux.scala 81:58]
  reg [1:0] source; // @[Counter.scala 61:40]
  wire [1:0] _source_wrap_value_T_1 = source + 2'h1; // @[Counter.scala 77:24]
  SRAM array ( // @[ICache.scala 50:21]
    .clock(array_clock),
    .io_en(array_io_en),
    .io_addr(array_io_addr),
    .io_wdata(array_io_wdata),
    .io_wen(array_io_wen),
    .io_rdata(array_io_rdata)
  );
  assign auto_out_a_valid = state == 3'h1; // @[ICache.scala 150:24]
  assign auto_out_a_bits_source = source; // @[Edges.scala 447:17 451:15]
  assign auto_out_a_bits_address = {req_r_addr[31:5],5'h0}; // @[Cat.scala 33:92]
  assign auto_out_d_ready = state == 3'h2; // @[ICache.scala 152:24]
  assign io_cache_req_ready = (state == 3'h0 & array_hit | state == 3'h3 | state == 3'h4) & io_cache_resp_ready; // @[ICache.scala 143:92]
  assign io_cache_resp_valid = _s2_ready_T_1 | _s2_ready_T_2; // @[ICache.scala 156:55]
  assign io_cache_resp_bits_rdata = _s2_ready_T_2 ? refill_data : _GEN_530; // @[ICache.scala 158:25]
  assign array_clock = clock;
  assign array_io_en = fire | _array_io_en_T; // @[ICache.scala 59:26]
  assign array_io_addr = _array_io_en_T ? req_r_addr[13:5] : _GEN_513; // @[ICache.scala 124:19 125:33]
  assign array_io_wdata = _array_io_en_T ? _array_io_wdata_T_1 : 274'h0; // @[ICache.scala 124:19 126:33 61:18]
  assign array_io_wen = tl_d_ready & auto_out_d_valid; // @[Decoupled.scala 51:35]
  always @(posedge clock) begin
    if (reset) begin // @[ICache.scala 48:22]
      req_r_addr <= 39'h0; // @[ICache.scala 48:22]
    end else if (fire) begin // @[ICache.scala 71:14]
      req_r_addr <= io_cache_req_bits_addr; // @[ICache.scala 73:19]
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_0 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_0 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_0 <= _GEN_532;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_1 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_1 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_1 <= _GEN_533;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_2 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_2 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_2 <= _GEN_534;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_3 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_3 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_3 <= _GEN_535;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_4 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_4 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_4 <= _GEN_536;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_5 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_5 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_5 <= _GEN_537;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_6 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_6 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_6 <= _GEN_538;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_7 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_7 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_7 <= _GEN_539;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_8 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_8 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_8 <= _GEN_540;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_9 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_9 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_9 <= _GEN_541;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_10 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_10 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_10 <= _GEN_542;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_11 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_11 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_11 <= _GEN_543;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_12 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_12 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_12 <= _GEN_544;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_13 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_13 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_13 <= _GEN_545;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_14 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_14 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_14 <= _GEN_546;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_15 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_15 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_15 <= _GEN_547;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_16 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_16 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_16 <= _GEN_548;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_17 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_17 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_17 <= _GEN_549;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_18 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_18 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_18 <= _GEN_550;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_19 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_19 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_19 <= _GEN_551;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_20 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_20 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_20 <= _GEN_552;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_21 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_21 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_21 <= _GEN_553;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_22 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_22 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_22 <= _GEN_554;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_23 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_23 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_23 <= _GEN_555;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_24 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_24 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_24 <= _GEN_556;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_25 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_25 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_25 <= _GEN_557;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_26 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_26 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_26 <= _GEN_558;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_27 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_27 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_27 <= _GEN_559;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_28 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_28 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_28 <= _GEN_560;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_29 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_29 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_29 <= _GEN_561;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_30 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_30 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_30 <= _GEN_562;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_31 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_31 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_31 <= _GEN_563;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_32 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_32 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_32 <= _GEN_564;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_33 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_33 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_33 <= _GEN_565;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_34 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_34 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_34 <= _GEN_566;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_35 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_35 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_35 <= _GEN_567;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_36 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_36 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_36 <= _GEN_568;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_37 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_37 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_37 <= _GEN_569;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_38 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_38 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_38 <= _GEN_570;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_39 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_39 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_39 <= _GEN_571;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_40 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_40 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_40 <= _GEN_572;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_41 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_41 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_41 <= _GEN_573;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_42 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_42 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_42 <= _GEN_574;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_43 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_43 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_43 <= _GEN_575;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_44 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_44 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_44 <= _GEN_576;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_45 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_45 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_45 <= _GEN_577;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_46 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_46 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_46 <= _GEN_578;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_47 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_47 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_47 <= _GEN_579;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_48 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_48 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_48 <= _GEN_580;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_49 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_49 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_49 <= _GEN_581;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_50 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_50 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_50 <= _GEN_582;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_51 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_51 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_51 <= _GEN_583;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_52 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_52 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_52 <= _GEN_584;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_53 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_53 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_53 <= _GEN_585;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_54 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_54 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_54 <= _GEN_586;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_55 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_55 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_55 <= _GEN_587;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_56 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_56 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_56 <= _GEN_588;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_57 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_57 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_57 <= _GEN_589;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_58 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_58 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_58 <= _GEN_590;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_59 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_59 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_59 <= _GEN_591;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_60 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_60 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_60 <= _GEN_592;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_61 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_61 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_61 <= _GEN_593;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_62 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_62 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_62 <= _GEN_594;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_63 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_63 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_63 <= _GEN_595;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_64 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_64 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_64 <= _GEN_596;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_65 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_65 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_65 <= _GEN_597;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_66 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_66 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_66 <= _GEN_598;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_67 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_67 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_67 <= _GEN_599;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_68 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_68 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_68 <= _GEN_600;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_69 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_69 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_69 <= _GEN_601;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_70 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_70 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_70 <= _GEN_602;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_71 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_71 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_71 <= _GEN_603;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_72 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_72 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_72 <= _GEN_604;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_73 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_73 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_73 <= _GEN_605;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_74 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_74 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_74 <= _GEN_606;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_75 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_75 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_75 <= _GEN_607;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_76 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_76 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_76 <= _GEN_608;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_77 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_77 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_77 <= _GEN_609;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_78 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_78 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_78 <= _GEN_610;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_79 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_79 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_79 <= _GEN_611;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_80 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_80 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_80 <= _GEN_612;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_81 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_81 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_81 <= _GEN_613;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_82 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_82 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_82 <= _GEN_614;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_83 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_83 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_83 <= _GEN_615;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_84 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_84 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_84 <= _GEN_616;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_85 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_85 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_85 <= _GEN_617;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_86 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_86 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_86 <= _GEN_618;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_87 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_87 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_87 <= _GEN_619;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_88 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_88 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_88 <= _GEN_620;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_89 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_89 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_89 <= _GEN_621;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_90 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_90 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_90 <= _GEN_622;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_91 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_91 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_91 <= _GEN_623;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_92 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_92 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_92 <= _GEN_624;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_93 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_93 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_93 <= _GEN_625;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_94 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_94 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_94 <= _GEN_626;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_95 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_95 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_95 <= _GEN_627;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_96 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_96 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_96 <= _GEN_628;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_97 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_97 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_97 <= _GEN_629;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_98 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_98 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_98 <= _GEN_630;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_99 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_99 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_99 <= _GEN_631;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_100 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_100 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_100 <= _GEN_632;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_101 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_101 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_101 <= _GEN_633;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_102 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_102 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_102 <= _GEN_634;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_103 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_103 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_103 <= _GEN_635;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_104 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_104 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_104 <= _GEN_636;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_105 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_105 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_105 <= _GEN_637;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_106 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_106 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_106 <= _GEN_638;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_107 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_107 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_107 <= _GEN_639;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_108 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_108 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_108 <= _GEN_640;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_109 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_109 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_109 <= _GEN_641;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_110 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_110 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_110 <= _GEN_642;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_111 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_111 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_111 <= _GEN_643;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_112 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_112 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_112 <= _GEN_644;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_113 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_113 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_113 <= _GEN_645;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_114 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_114 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_114 <= _GEN_646;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_115 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_115 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_115 <= _GEN_647;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_116 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_116 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_116 <= _GEN_648;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_117 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_117 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_117 <= _GEN_649;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_118 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_118 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_118 <= _GEN_650;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_119 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_119 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_119 <= _GEN_651;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_120 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_120 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_120 <= _GEN_652;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_121 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_121 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_121 <= _GEN_653;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_122 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_122 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_122 <= _GEN_654;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_123 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_123 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_123 <= _GEN_655;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_124 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_124 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_124 <= _GEN_656;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_125 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_125 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_125 <= _GEN_657;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_126 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_126 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_126 <= _GEN_658;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_127 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_127 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_127 <= _GEN_659;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_128 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_128 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_128 <= _GEN_660;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_129 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_129 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_129 <= _GEN_661;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_130 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_130 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_130 <= _GEN_662;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_131 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_131 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_131 <= _GEN_663;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_132 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_132 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_132 <= _GEN_664;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_133 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_133 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_133 <= _GEN_665;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_134 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_134 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_134 <= _GEN_666;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_135 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_135 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_135 <= _GEN_667;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_136 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_136 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_136 <= _GEN_668;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_137 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_137 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_137 <= _GEN_669;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_138 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_138 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_138 <= _GEN_670;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_139 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_139 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_139 <= _GEN_671;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_140 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_140 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_140 <= _GEN_672;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_141 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_141 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_141 <= _GEN_673;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_142 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_142 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_142 <= _GEN_674;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_143 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_143 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_143 <= _GEN_675;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_144 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_144 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_144 <= _GEN_676;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_145 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_145 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_145 <= _GEN_677;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_146 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_146 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_146 <= _GEN_678;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_147 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_147 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_147 <= _GEN_679;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_148 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_148 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_148 <= _GEN_680;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_149 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_149 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_149 <= _GEN_681;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_150 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_150 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_150 <= _GEN_682;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_151 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_151 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_151 <= _GEN_683;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_152 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_152 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_152 <= _GEN_684;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_153 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_153 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_153 <= _GEN_685;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_154 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_154 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_154 <= _GEN_686;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_155 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_155 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_155 <= _GEN_687;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_156 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_156 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_156 <= _GEN_688;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_157 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_157 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_157 <= _GEN_689;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_158 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_158 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_158 <= _GEN_690;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_159 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_159 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_159 <= _GEN_691;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_160 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_160 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_160 <= _GEN_692;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_161 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_161 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_161 <= _GEN_693;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_162 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_162 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_162 <= _GEN_694;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_163 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_163 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_163 <= _GEN_695;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_164 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_164 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_164 <= _GEN_696;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_165 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_165 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_165 <= _GEN_697;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_166 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_166 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_166 <= _GEN_698;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_167 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_167 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_167 <= _GEN_699;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_168 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_168 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_168 <= _GEN_700;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_169 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_169 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_169 <= _GEN_701;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_170 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_170 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_170 <= _GEN_702;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_171 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_171 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_171 <= _GEN_703;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_172 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_172 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_172 <= _GEN_704;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_173 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_173 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_173 <= _GEN_705;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_174 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_174 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_174 <= _GEN_706;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_175 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_175 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_175 <= _GEN_707;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_176 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_176 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_176 <= _GEN_708;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_177 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_177 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_177 <= _GEN_709;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_178 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_178 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_178 <= _GEN_710;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_179 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_179 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_179 <= _GEN_711;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_180 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_180 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_180 <= _GEN_712;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_181 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_181 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_181 <= _GEN_713;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_182 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_182 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_182 <= _GEN_714;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_183 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_183 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_183 <= _GEN_715;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_184 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_184 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_184 <= _GEN_716;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_185 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_185 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_185 <= _GEN_717;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_186 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_186 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_186 <= _GEN_718;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_187 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_187 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_187 <= _GEN_719;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_188 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_188 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_188 <= _GEN_720;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_189 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_189 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_189 <= _GEN_721;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_190 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_190 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_190 <= _GEN_722;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_191 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_191 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_191 <= _GEN_723;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_192 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_192 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_192 <= _GEN_724;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_193 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_193 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_193 <= _GEN_725;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_194 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_194 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_194 <= _GEN_726;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_195 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_195 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_195 <= _GEN_727;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_196 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_196 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_196 <= _GEN_728;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_197 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_197 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_197 <= _GEN_729;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_198 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_198 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_198 <= _GEN_730;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_199 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_199 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_199 <= _GEN_731;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_200 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_200 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_200 <= _GEN_732;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_201 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_201 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_201 <= _GEN_733;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_202 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_202 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_202 <= _GEN_734;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_203 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_203 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_203 <= _GEN_735;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_204 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_204 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_204 <= _GEN_736;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_205 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_205 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_205 <= _GEN_737;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_206 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_206 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_206 <= _GEN_738;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_207 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_207 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_207 <= _GEN_739;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_208 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_208 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_208 <= _GEN_740;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_209 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_209 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_209 <= _GEN_741;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_210 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_210 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_210 <= _GEN_742;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_211 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_211 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_211 <= _GEN_743;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_212 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_212 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_212 <= _GEN_744;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_213 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_213 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_213 <= _GEN_745;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_214 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_214 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_214 <= _GEN_746;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_215 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_215 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_215 <= _GEN_747;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_216 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_216 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_216 <= _GEN_748;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_217 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_217 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_217 <= _GEN_749;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_218 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_218 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_218 <= _GEN_750;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_219 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_219 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_219 <= _GEN_751;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_220 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_220 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_220 <= _GEN_752;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_221 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_221 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_221 <= _GEN_753;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_222 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_222 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_222 <= _GEN_754;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_223 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_223 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_223 <= _GEN_755;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_224 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_224 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_224 <= _GEN_756;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_225 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_225 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_225 <= _GEN_757;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_226 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_226 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_226 <= _GEN_758;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_227 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_227 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_227 <= _GEN_759;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_228 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_228 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_228 <= _GEN_760;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_229 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_229 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_229 <= _GEN_761;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_230 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_230 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_230 <= _GEN_762;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_231 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_231 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_231 <= _GEN_763;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_232 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_232 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_232 <= _GEN_764;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_233 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_233 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_233 <= _GEN_765;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_234 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_234 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_234 <= _GEN_766;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_235 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_235 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_235 <= _GEN_767;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_236 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_236 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_236 <= _GEN_768;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_237 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_237 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_237 <= _GEN_769;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_238 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_238 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_238 <= _GEN_770;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_239 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_239 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_239 <= _GEN_771;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_240 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_240 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_240 <= _GEN_772;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_241 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_241 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_241 <= _GEN_773;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_242 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_242 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_242 <= _GEN_774;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_243 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_243 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_243 <= _GEN_775;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_244 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_244 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_244 <= _GEN_776;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_245 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_245 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_245 <= _GEN_777;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_246 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_246 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_246 <= _GEN_778;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_247 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_247 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_247 <= _GEN_779;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_248 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_248 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_248 <= _GEN_780;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_249 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_249 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_249 <= _GEN_781;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_250 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_250 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_250 <= _GEN_782;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_251 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_251 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_251 <= _GEN_783;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_252 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_252 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_252 <= _GEN_784;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_253 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_253 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_253 <= _GEN_785;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_254 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_254 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_254 <= _GEN_786;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_255 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_255 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_255 <= _GEN_787;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_256 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_256 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_256 <= _GEN_788;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_257 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_257 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_257 <= _GEN_789;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_258 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_258 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_258 <= _GEN_790;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_259 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_259 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_259 <= _GEN_791;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_260 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_260 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_260 <= _GEN_792;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_261 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_261 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_261 <= _GEN_793;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_262 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_262 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_262 <= _GEN_794;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_263 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_263 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_263 <= _GEN_795;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_264 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_264 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_264 <= _GEN_796;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_265 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_265 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_265 <= _GEN_797;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_266 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_266 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_266 <= _GEN_798;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_267 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_267 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_267 <= _GEN_799;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_268 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_268 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_268 <= _GEN_800;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_269 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_269 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_269 <= _GEN_801;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_270 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_270 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_270 <= _GEN_802;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_271 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_271 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_271 <= _GEN_803;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_272 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_272 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_272 <= _GEN_804;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_273 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_273 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_273 <= _GEN_805;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_274 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_274 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_274 <= _GEN_806;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_275 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_275 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_275 <= _GEN_807;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_276 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_276 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_276 <= _GEN_808;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_277 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_277 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_277 <= _GEN_809;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_278 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_278 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_278 <= _GEN_810;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_279 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_279 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_279 <= _GEN_811;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_280 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_280 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_280 <= _GEN_812;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_281 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_281 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_281 <= _GEN_813;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_282 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_282 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_282 <= _GEN_814;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_283 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_283 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_283 <= _GEN_815;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_284 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_284 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_284 <= _GEN_816;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_285 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_285 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_285 <= _GEN_817;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_286 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_286 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_286 <= _GEN_818;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_287 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_287 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_287 <= _GEN_819;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_288 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_288 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_288 <= _GEN_820;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_289 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_289 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_289 <= _GEN_821;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_290 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_290 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_290 <= _GEN_822;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_291 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_291 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_291 <= _GEN_823;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_292 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_292 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_292 <= _GEN_824;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_293 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_293 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_293 <= _GEN_825;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_294 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_294 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_294 <= _GEN_826;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_295 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_295 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_295 <= _GEN_827;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_296 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_296 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_296 <= _GEN_828;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_297 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_297 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_297 <= _GEN_829;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_298 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_298 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_298 <= _GEN_830;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_299 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_299 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_299 <= _GEN_831;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_300 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_300 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_300 <= _GEN_832;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_301 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_301 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_301 <= _GEN_833;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_302 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_302 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_302 <= _GEN_834;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_303 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_303 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_303 <= _GEN_835;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_304 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_304 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_304 <= _GEN_836;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_305 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_305 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_305 <= _GEN_837;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_306 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_306 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_306 <= _GEN_838;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_307 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_307 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_307 <= _GEN_839;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_308 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_308 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_308 <= _GEN_840;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_309 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_309 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_309 <= _GEN_841;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_310 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_310 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_310 <= _GEN_842;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_311 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_311 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_311 <= _GEN_843;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_312 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_312 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_312 <= _GEN_844;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_313 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_313 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_313 <= _GEN_845;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_314 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_314 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_314 <= _GEN_846;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_315 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_315 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_315 <= _GEN_847;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_316 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_316 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_316 <= _GEN_848;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_317 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_317 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_317 <= _GEN_849;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_318 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_318 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_318 <= _GEN_850;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_319 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_319 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_319 <= _GEN_851;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_320 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_320 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_320 <= _GEN_852;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_321 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_321 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_321 <= _GEN_853;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_322 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_322 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_322 <= _GEN_854;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_323 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_323 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_323 <= _GEN_855;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_324 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_324 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_324 <= _GEN_856;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_325 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_325 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_325 <= _GEN_857;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_326 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_326 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_326 <= _GEN_858;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_327 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_327 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_327 <= _GEN_859;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_328 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_328 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_328 <= _GEN_860;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_329 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_329 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_329 <= _GEN_861;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_330 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_330 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_330 <= _GEN_862;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_331 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_331 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_331 <= _GEN_863;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_332 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_332 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_332 <= _GEN_864;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_333 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_333 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_333 <= _GEN_865;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_334 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_334 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_334 <= _GEN_866;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_335 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_335 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_335 <= _GEN_867;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_336 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_336 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_336 <= _GEN_868;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_337 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_337 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_337 <= _GEN_869;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_338 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_338 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_338 <= _GEN_870;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_339 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_339 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_339 <= _GEN_871;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_340 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_340 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_340 <= _GEN_872;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_341 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_341 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_341 <= _GEN_873;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_342 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_342 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_342 <= _GEN_874;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_343 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_343 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_343 <= _GEN_875;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_344 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_344 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_344 <= _GEN_876;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_345 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_345 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_345 <= _GEN_877;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_346 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_346 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_346 <= _GEN_878;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_347 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_347 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_347 <= _GEN_879;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_348 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_348 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_348 <= _GEN_880;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_349 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_349 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_349 <= _GEN_881;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_350 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_350 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_350 <= _GEN_882;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_351 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_351 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_351 <= _GEN_883;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_352 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_352 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_352 <= _GEN_884;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_353 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_353 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_353 <= _GEN_885;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_354 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_354 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_354 <= _GEN_886;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_355 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_355 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_355 <= _GEN_887;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_356 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_356 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_356 <= _GEN_888;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_357 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_357 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_357 <= _GEN_889;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_358 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_358 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_358 <= _GEN_890;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_359 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_359 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_359 <= _GEN_891;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_360 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_360 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_360 <= _GEN_892;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_361 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_361 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_361 <= _GEN_893;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_362 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_362 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_362 <= _GEN_894;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_363 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_363 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_363 <= _GEN_895;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_364 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_364 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_364 <= _GEN_896;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_365 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_365 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_365 <= _GEN_897;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_366 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_366 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_366 <= _GEN_898;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_367 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_367 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_367 <= _GEN_899;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_368 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_368 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_368 <= _GEN_900;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_369 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_369 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_369 <= _GEN_901;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_370 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_370 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_370 <= _GEN_902;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_371 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_371 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_371 <= _GEN_903;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_372 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_372 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_372 <= _GEN_904;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_373 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_373 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_373 <= _GEN_905;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_374 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_374 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_374 <= _GEN_906;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_375 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_375 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_375 <= _GEN_907;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_376 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_376 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_376 <= _GEN_908;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_377 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_377 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_377 <= _GEN_909;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_378 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_378 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_378 <= _GEN_910;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_379 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_379 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_379 <= _GEN_911;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_380 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_380 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_380 <= _GEN_912;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_381 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_381 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_381 <= _GEN_913;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_382 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_382 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_382 <= _GEN_914;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_383 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_383 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_383 <= _GEN_915;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_384 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_384 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_384 <= _GEN_916;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_385 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_385 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_385 <= _GEN_917;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_386 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_386 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_386 <= _GEN_918;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_387 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_387 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_387 <= _GEN_919;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_388 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_388 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_388 <= _GEN_920;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_389 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_389 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_389 <= _GEN_921;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_390 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_390 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_390 <= _GEN_922;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_391 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_391 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_391 <= _GEN_923;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_392 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_392 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_392 <= _GEN_924;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_393 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_393 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_393 <= _GEN_925;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_394 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_394 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_394 <= _GEN_926;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_395 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_395 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_395 <= _GEN_927;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_396 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_396 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_396 <= _GEN_928;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_397 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_397 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_397 <= _GEN_929;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_398 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_398 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_398 <= _GEN_930;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_399 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_399 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_399 <= _GEN_931;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_400 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_400 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_400 <= _GEN_932;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_401 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_401 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_401 <= _GEN_933;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_402 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_402 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_402 <= _GEN_934;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_403 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_403 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_403 <= _GEN_935;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_404 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_404 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_404 <= _GEN_936;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_405 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_405 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_405 <= _GEN_937;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_406 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_406 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_406 <= _GEN_938;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_407 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_407 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_407 <= _GEN_939;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_408 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_408 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_408 <= _GEN_940;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_409 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_409 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_409 <= _GEN_941;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_410 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_410 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_410 <= _GEN_942;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_411 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_411 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_411 <= _GEN_943;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_412 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_412 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_412 <= _GEN_944;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_413 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_413 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_413 <= _GEN_945;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_414 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_414 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_414 <= _GEN_946;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_415 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_415 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_415 <= _GEN_947;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_416 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_416 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_416 <= _GEN_948;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_417 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_417 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_417 <= _GEN_949;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_418 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_418 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_418 <= _GEN_950;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_419 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_419 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_419 <= _GEN_951;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_420 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_420 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_420 <= _GEN_952;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_421 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_421 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_421 <= _GEN_953;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_422 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_422 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_422 <= _GEN_954;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_423 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_423 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_423 <= _GEN_955;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_424 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_424 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_424 <= _GEN_956;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_425 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_425 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_425 <= _GEN_957;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_426 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_426 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_426 <= _GEN_958;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_427 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_427 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_427 <= _GEN_959;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_428 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_428 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_428 <= _GEN_960;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_429 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_429 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_429 <= _GEN_961;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_430 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_430 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_430 <= _GEN_962;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_431 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_431 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_431 <= _GEN_963;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_432 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_432 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_432 <= _GEN_964;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_433 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_433 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_433 <= _GEN_965;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_434 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_434 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_434 <= _GEN_966;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_435 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_435 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_435 <= _GEN_967;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_436 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_436 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_436 <= _GEN_968;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_437 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_437 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_437 <= _GEN_969;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_438 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_438 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_438 <= _GEN_970;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_439 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_439 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_439 <= _GEN_971;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_440 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_440 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_440 <= _GEN_972;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_441 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_441 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_441 <= _GEN_973;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_442 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_442 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_442 <= _GEN_974;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_443 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_443 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_443 <= _GEN_975;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_444 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_444 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_444 <= _GEN_976;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_445 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_445 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_445 <= _GEN_977;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_446 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_446 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_446 <= _GEN_978;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_447 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_447 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_447 <= _GEN_979;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_448 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_448 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_448 <= _GEN_980;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_449 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_449 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_449 <= _GEN_981;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_450 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_450 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_450 <= _GEN_982;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_451 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_451 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_451 <= _GEN_983;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_452 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_452 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_452 <= _GEN_984;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_453 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_453 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_453 <= _GEN_985;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_454 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_454 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_454 <= _GEN_986;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_455 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_455 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_455 <= _GEN_987;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_456 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_456 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_456 <= _GEN_988;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_457 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_457 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_457 <= _GEN_989;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_458 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_458 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_458 <= _GEN_990;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_459 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_459 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_459 <= _GEN_991;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_460 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_460 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_460 <= _GEN_992;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_461 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_461 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_461 <= _GEN_993;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_462 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_462 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_462 <= _GEN_994;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_463 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_463 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_463 <= _GEN_995;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_464 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_464 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_464 <= _GEN_996;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_465 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_465 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_465 <= _GEN_997;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_466 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_466 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_466 <= _GEN_998;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_467 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_467 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_467 <= _GEN_999;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_468 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_468 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_468 <= _GEN_1000;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_469 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_469 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_469 <= _GEN_1001;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_470 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_470 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_470 <= _GEN_1002;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_471 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_471 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_471 <= _GEN_1003;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_472 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_472 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_472 <= _GEN_1004;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_473 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_473 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_473 <= _GEN_1005;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_474 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_474 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_474 <= _GEN_1006;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_475 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_475 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_475 <= _GEN_1007;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_476 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_476 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_476 <= _GEN_1008;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_477 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_477 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_477 <= _GEN_1009;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_478 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_478 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_478 <= _GEN_1010;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_479 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_479 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_479 <= _GEN_1011;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_480 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_480 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_480 <= _GEN_1012;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_481 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_481 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_481 <= _GEN_1013;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_482 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_482 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_482 <= _GEN_1014;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_483 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_483 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_483 <= _GEN_1015;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_484 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_484 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_484 <= _GEN_1016;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_485 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_485 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_485 <= _GEN_1017;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_486 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_486 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_486 <= _GEN_1018;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_487 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_487 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_487 <= _GEN_1019;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_488 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_488 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_488 <= _GEN_1020;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_489 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_489 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_489 <= _GEN_1021;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_490 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_490 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_490 <= _GEN_1022;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_491 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_491 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_491 <= _GEN_1023;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_492 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_492 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_492 <= _GEN_1024;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_493 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_493 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_493 <= _GEN_1025;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_494 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_494 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_494 <= _GEN_1026;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_495 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_495 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_495 <= _GEN_1027;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_496 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_496 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_496 <= _GEN_1028;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_497 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_497 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_497 <= _GEN_1029;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_498 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_498 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_498 <= _GEN_1030;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_499 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_499 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_499 <= _GEN_1031;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_500 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_500 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_500 <= _GEN_1032;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_501 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_501 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_501 <= _GEN_1033;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_502 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_502 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_502 <= _GEN_1034;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_503 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_503 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_503 <= _GEN_1035;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_504 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_504 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_504 <= _GEN_1036;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_505 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_505 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_505 <= _GEN_1037;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_506 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_506 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_506 <= _GEN_1038;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_507 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_507 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_507 <= _GEN_1039;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_508 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_508 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_508 <= _GEN_1040;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_509 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_509 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_509 <= _GEN_1041;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_510 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_510 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_510 <= _GEN_1042;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_511 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_511 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_511 <= _GEN_1043;
    end
    if (reset) begin // @[ICache.scala 78:68]
      state <= 3'h4; // @[ICache.scala 78:68]
    end else if (3'h0 == state) begin // @[ICache.scala 80:17]
      if (_state_T & ~_state_T_1) begin // @[ICache.scala 82:19]
        state <= 3'h4;
      end else if (array_hit) begin // @[ICache.scala 82:55]
        state <= 3'h0;
      end else begin
        state <= 3'h1;
      end
    end else if (3'h1 == state) begin // @[ICache.scala 80:17]
      if (_T_2) begin // @[ICache.scala 85:23]
        state <= 3'h2; // @[ICache.scala 86:15]
      end
    end else if (3'h2 == state) begin // @[ICache.scala 80:17]
      state <= _GEN_522;
    end else begin
      state <= _GEN_526;
    end
    array_out_REG <= io_cache_req_valid & s2_ready; // @[ICache.scala 56:27]
    if (reset) begin // @[Reg.scala 35:20]
      array_out_r <= 274'h0; // @[Reg.scala 35:20]
    end else if (array_out_REG) begin // @[Utils.scala 50:8]
      array_out_r <= array_io_rdata;
    end
    array_data_REG <= io_cache_req_ready & io_cache_req_valid; // @[Decoupled.scala 51:35]
    if (reset) begin // @[Reg.scala 35:20]
      array_data_r <= 64'h0; // @[Reg.scala 35:20]
    end else if (array_data_REG) begin // @[Reg.scala 36:18]
      if (2'h3 == req_r_addr[4:3]) begin // @[Mux.scala 81:58]
        array_data_r <= array_out_data[255:192];
      end else if (2'h2 == req_r_addr[4:3]) begin // @[Mux.scala 81:58]
        array_data_r <= array_out_data[191:128];
      end else begin
        array_data_r <= _array_data_T_6;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      wdata <= 256'h0; // @[Reg.scala 35:20]
    end else if (_array_io_en_T) begin // @[Reg.scala 36:18]
      wdata <= auto_out_d_bits_data; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Counter.scala 61:40]
      source <= 2'h0; // @[Counter.scala 61:40]
    end else if (_T_2) begin // @[Counter.scala 118:16]
      source <= _source_wrap_value_T_1; // @[Counter.scala 77:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  req_r_addr = _RAND_0[38:0];
  _RAND_1 = {1{`RANDOM}};
  valid_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  valid_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  valid_2 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  valid_3 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  valid_4 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  valid_5 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  valid_6 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  valid_7 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  valid_8 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  valid_9 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  valid_10 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  valid_11 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  valid_12 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  valid_13 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  valid_14 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  valid_15 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  valid_16 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  valid_17 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  valid_18 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  valid_19 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  valid_20 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  valid_21 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  valid_22 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  valid_23 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  valid_24 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  valid_25 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  valid_26 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  valid_27 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  valid_28 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  valid_29 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  valid_30 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  valid_31 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  valid_32 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  valid_33 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  valid_34 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  valid_35 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  valid_36 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  valid_37 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  valid_38 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  valid_39 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  valid_40 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  valid_41 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  valid_42 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  valid_43 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  valid_44 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  valid_45 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  valid_46 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  valid_47 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  valid_48 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  valid_49 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  valid_50 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  valid_51 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  valid_52 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  valid_53 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  valid_54 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  valid_55 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  valid_56 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  valid_57 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  valid_58 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  valid_59 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  valid_60 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  valid_61 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  valid_62 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  valid_63 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  valid_64 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  valid_65 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  valid_66 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  valid_67 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  valid_68 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  valid_69 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  valid_70 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  valid_71 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  valid_72 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  valid_73 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  valid_74 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  valid_75 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  valid_76 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  valid_77 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  valid_78 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  valid_79 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  valid_80 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  valid_81 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  valid_82 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  valid_83 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  valid_84 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  valid_85 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  valid_86 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  valid_87 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  valid_88 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  valid_89 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  valid_90 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  valid_91 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  valid_92 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  valid_93 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  valid_94 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  valid_95 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  valid_96 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  valid_97 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  valid_98 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  valid_99 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  valid_100 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  valid_101 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  valid_102 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  valid_103 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  valid_104 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  valid_105 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  valid_106 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  valid_107 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  valid_108 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  valid_109 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  valid_110 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  valid_111 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  valid_112 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  valid_113 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  valid_114 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  valid_115 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  valid_116 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  valid_117 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  valid_118 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  valid_119 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  valid_120 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  valid_121 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  valid_122 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  valid_123 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  valid_124 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  valid_125 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  valid_126 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  valid_127 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  valid_128 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  valid_129 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  valid_130 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  valid_131 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  valid_132 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  valid_133 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  valid_134 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  valid_135 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  valid_136 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  valid_137 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  valid_138 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  valid_139 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  valid_140 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  valid_141 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  valid_142 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  valid_143 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  valid_144 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  valid_145 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  valid_146 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  valid_147 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  valid_148 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  valid_149 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  valid_150 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  valid_151 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  valid_152 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  valid_153 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  valid_154 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  valid_155 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  valid_156 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  valid_157 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  valid_158 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  valid_159 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  valid_160 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  valid_161 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  valid_162 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  valid_163 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  valid_164 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  valid_165 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  valid_166 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  valid_167 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  valid_168 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  valid_169 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  valid_170 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  valid_171 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  valid_172 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  valid_173 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  valid_174 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  valid_175 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  valid_176 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  valid_177 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  valid_178 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  valid_179 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  valid_180 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  valid_181 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  valid_182 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  valid_183 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  valid_184 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  valid_185 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  valid_186 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  valid_187 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  valid_188 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  valid_189 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  valid_190 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  valid_191 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  valid_192 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  valid_193 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  valid_194 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  valid_195 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  valid_196 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  valid_197 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  valid_198 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  valid_199 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  valid_200 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  valid_201 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  valid_202 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  valid_203 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  valid_204 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  valid_205 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  valid_206 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  valid_207 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  valid_208 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  valid_209 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  valid_210 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  valid_211 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  valid_212 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  valid_213 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  valid_214 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  valid_215 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  valid_216 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  valid_217 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  valid_218 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  valid_219 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  valid_220 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  valid_221 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  valid_222 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  valid_223 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  valid_224 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  valid_225 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  valid_226 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  valid_227 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  valid_228 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  valid_229 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  valid_230 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  valid_231 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  valid_232 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  valid_233 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  valid_234 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  valid_235 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  valid_236 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  valid_237 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  valid_238 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  valid_239 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  valid_240 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  valid_241 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  valid_242 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  valid_243 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  valid_244 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  valid_245 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  valid_246 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  valid_247 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  valid_248 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  valid_249 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  valid_250 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  valid_251 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  valid_252 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  valid_253 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  valid_254 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  valid_255 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  valid_256 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  valid_257 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  valid_258 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  valid_259 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  valid_260 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  valid_261 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  valid_262 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  valid_263 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  valid_264 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  valid_265 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  valid_266 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  valid_267 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  valid_268 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  valid_269 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  valid_270 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  valid_271 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  valid_272 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  valid_273 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  valid_274 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  valid_275 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  valid_276 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  valid_277 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  valid_278 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  valid_279 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  valid_280 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  valid_281 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  valid_282 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  valid_283 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  valid_284 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  valid_285 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  valid_286 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  valid_287 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  valid_288 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  valid_289 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  valid_290 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  valid_291 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  valid_292 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  valid_293 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  valid_294 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  valid_295 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  valid_296 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  valid_297 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  valid_298 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  valid_299 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  valid_300 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  valid_301 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  valid_302 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  valid_303 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  valid_304 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  valid_305 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  valid_306 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  valid_307 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  valid_308 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  valid_309 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  valid_310 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  valid_311 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  valid_312 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  valid_313 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  valid_314 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  valid_315 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  valid_316 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  valid_317 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  valid_318 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  valid_319 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  valid_320 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  valid_321 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  valid_322 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  valid_323 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  valid_324 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  valid_325 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  valid_326 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  valid_327 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  valid_328 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  valid_329 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  valid_330 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  valid_331 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  valid_332 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  valid_333 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  valid_334 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  valid_335 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  valid_336 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  valid_337 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  valid_338 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  valid_339 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  valid_340 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  valid_341 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  valid_342 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  valid_343 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  valid_344 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  valid_345 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  valid_346 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  valid_347 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  valid_348 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  valid_349 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  valid_350 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  valid_351 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  valid_352 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  valid_353 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  valid_354 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  valid_355 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  valid_356 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  valid_357 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  valid_358 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  valid_359 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  valid_360 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  valid_361 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  valid_362 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  valid_363 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  valid_364 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  valid_365 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  valid_366 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  valid_367 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  valid_368 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  valid_369 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  valid_370 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  valid_371 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  valid_372 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  valid_373 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  valid_374 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  valid_375 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  valid_376 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  valid_377 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  valid_378 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  valid_379 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  valid_380 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  valid_381 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  valid_382 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  valid_383 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  valid_384 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  valid_385 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  valid_386 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  valid_387 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  valid_388 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  valid_389 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  valid_390 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  valid_391 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  valid_392 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  valid_393 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  valid_394 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  valid_395 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  valid_396 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  valid_397 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  valid_398 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  valid_399 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  valid_400 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  valid_401 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  valid_402 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  valid_403 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  valid_404 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  valid_405 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  valid_406 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  valid_407 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  valid_408 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  valid_409 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  valid_410 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  valid_411 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  valid_412 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  valid_413 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  valid_414 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  valid_415 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  valid_416 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  valid_417 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  valid_418 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  valid_419 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  valid_420 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  valid_421 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  valid_422 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  valid_423 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  valid_424 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  valid_425 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  valid_426 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  valid_427 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  valid_428 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  valid_429 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  valid_430 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  valid_431 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  valid_432 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  valid_433 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  valid_434 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  valid_435 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  valid_436 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  valid_437 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  valid_438 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  valid_439 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  valid_440 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  valid_441 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  valid_442 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  valid_443 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  valid_444 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  valid_445 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  valid_446 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  valid_447 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  valid_448 = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  valid_449 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  valid_450 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  valid_451 = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  valid_452 = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  valid_453 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  valid_454 = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  valid_455 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  valid_456 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  valid_457 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  valid_458 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  valid_459 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  valid_460 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  valid_461 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  valid_462 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  valid_463 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  valid_464 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  valid_465 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  valid_466 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  valid_467 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  valid_468 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  valid_469 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  valid_470 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  valid_471 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  valid_472 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  valid_473 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  valid_474 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  valid_475 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  valid_476 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  valid_477 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  valid_478 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  valid_479 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  valid_480 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  valid_481 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  valid_482 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  valid_483 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  valid_484 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  valid_485 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  valid_486 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  valid_487 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  valid_488 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  valid_489 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  valid_490 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  valid_491 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  valid_492 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  valid_493 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  valid_494 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  valid_495 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  valid_496 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  valid_497 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  valid_498 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  valid_499 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  valid_500 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  valid_501 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  valid_502 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  valid_503 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  valid_504 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  valid_505 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  valid_506 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  valid_507 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  valid_508 = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  valid_509 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  valid_510 = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  valid_511 = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  state = _RAND_513[2:0];
  _RAND_514 = {1{`RANDOM}};
  array_out_REG = _RAND_514[0:0];
  _RAND_515 = {9{`RANDOM}};
  array_out_r = _RAND_515[273:0];
  _RAND_516 = {1{`RANDOM}};
  array_data_REG = _RAND_516[0:0];
  _RAND_517 = {2{`RANDOM}};
  array_data_r = _RAND_517[63:0];
  _RAND_518 = {8{`RANDOM}};
  wdata = _RAND_518[255:0];
  _RAND_519 = {1{`RANDOM}};
  source = _RAND_519[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DCache(
  input          clock,
  input          reset,
  input          auto_out_a_ready,
  output         auto_out_a_valid,
  output [1:0]   auto_out_a_bits_source,
  output [31:0]  auto_out_a_bits_address,
  output         auto_out_b_ready,
  input          auto_out_b_valid,
  input  [2:0]   auto_out_b_bits_size,
  input  [1:0]   auto_out_b_bits_source,
  input  [31:0]  auto_out_b_bits_address,
  input          auto_out_c_ready,
  output         auto_out_c_valid,
  output [2:0]   auto_out_c_bits_opcode,
  output [2:0]   auto_out_c_bits_param,
  output [2:0]   auto_out_c_bits_size,
  output [1:0]   auto_out_c_bits_source,
  output [31:0]  auto_out_c_bits_address,
  output [255:0] auto_out_c_bits_data,
  output         auto_out_d_ready,
  input          auto_out_d_valid,
  input  [5:0]   auto_out_d_bits_sink,
  input  [255:0] auto_out_d_bits_data,
  input          auto_out_e_ready,
  output         auto_out_e_valid,
  output [5:0]   auto_out_e_bits_sink,
  output         io_cache_req_ready,
  input          io_cache_req_valid,
  input  [38:0]  io_cache_req_bits_addr,
  input  [63:0]  io_cache_req_bits_wdata,
  input  [7:0]   io_cache_req_bits_wmask,
  input          io_cache_req_bits_wen,
  input  [1:0]   io_cache_req_bits_len,
  input          io_cache_req_bits_lrsc,
  input  [4:0]   io_cache_req_bits_amo,
  input          io_cache_resp_ready,
  output         io_cache_resp_valid,
  output [63:0]  io_cache_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [255:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [287:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [287:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
`endif // RANDOMIZE_REG_INIT
  wire  array_clock; // @[DCache.scala 55:21]
  wire  array_io_en; // @[DCache.scala 55:21]
  wire [8:0] array_io_addr; // @[DCache.scala 55:21]
  wire [273:0] array_io_wdata; // @[DCache.scala 55:21]
  wire  array_io_wen; // @[DCache.scala 55:21]
  wire [273:0] array_io_rdata; // @[DCache.scala 55:21]
  reg  probing; // @[Utils.scala 36:20]
  wire  _x1_b_ready_T = ~probing; // @[DCache.scala 258:17]
  reg  lrsc_reserved; // @[DCache.scala 127:30]
  wire  _x1_b_ready_T_1 = ~lrsc_reserved; // @[DCache.scala 258:30]
  reg [4:0] lrsc_counter; // @[DCache.scala 129:30]
  wire  lrsc_backoff = lrsc_counter[4]; // @[DCache.scala 130:35]
  wire  tl_b_ready = ~probing & (~lrsc_reserved | lrsc_backoff); // @[DCache.scala 258:26]
  wire  _tl_b_bits_r_T = tl_b_ready & auto_out_b_valid; // @[Decoupled.scala 51:35]
  reg [2:0] tl_b_bits_r_size; // @[Reg.scala 35:20]
  reg [1:0] tl_b_bits_r_source; // @[Reg.scala 35:20]
  reg [31:0] tl_b_bits_r_address; // @[Reg.scala 35:20]
  wire [31:0] _GEN_4 = _tl_b_bits_r_T ? auto_out_b_bits_address : tl_b_bits_r_address; // @[Reg.scala 36:18 35:20 36:22]
  reg [2:0] state; // @[DCache.scala 60:118]
  wire  tl_d_ready = state == 3'h3 | state == 3'h5; // @[DCache.scala 261:43]
  wire  _tl_d_bits_r_T = tl_d_ready & auto_out_d_valid; // @[Decoupled.scala 51:35]
  reg [5:0] tl_d_bits_r_sink; // @[Reg.scala 35:20]
  reg [255:0] tl_d_bits_r_data; // @[Reg.scala 35:20]
  wire  _req_r_T = io_cache_req_ready & io_cache_req_valid; // @[Decoupled.scala 51:35]
  reg [38:0] req_r_addr; // @[Reg.scala 35:20]
  reg [63:0] req_r_wdata; // @[Reg.scala 35:20]
  reg [7:0] req_r_wmask; // @[Reg.scala 35:20]
  reg  req_r_wen; // @[Reg.scala 35:20]
  reg [1:0] req_r_len; // @[Reg.scala 35:20]
  reg  req_r_lrsc; // @[Reg.scala 35:20]
  reg [4:0] req_r_amo; // @[Reg.scala 35:20]
  wire [38:0] _GEN_16 = _req_r_T ? io_cache_req_bits_addr : req_r_addr; // @[Reg.scala 36:18 35:20 36:22]
  reg  valid_0; // @[DCache.scala 56:22]
  reg  valid_1; // @[DCache.scala 56:22]
  reg  valid_2; // @[DCache.scala 56:22]
  reg  valid_3; // @[DCache.scala 56:22]
  reg  valid_4; // @[DCache.scala 56:22]
  reg  valid_5; // @[DCache.scala 56:22]
  reg  valid_6; // @[DCache.scala 56:22]
  reg  valid_7; // @[DCache.scala 56:22]
  reg  valid_8; // @[DCache.scala 56:22]
  reg  valid_9; // @[DCache.scala 56:22]
  reg  valid_10; // @[DCache.scala 56:22]
  reg  valid_11; // @[DCache.scala 56:22]
  reg  valid_12; // @[DCache.scala 56:22]
  reg  valid_13; // @[DCache.scala 56:22]
  reg  valid_14; // @[DCache.scala 56:22]
  reg  valid_15; // @[DCache.scala 56:22]
  reg  valid_16; // @[DCache.scala 56:22]
  reg  valid_17; // @[DCache.scala 56:22]
  reg  valid_18; // @[DCache.scala 56:22]
  reg  valid_19; // @[DCache.scala 56:22]
  reg  valid_20; // @[DCache.scala 56:22]
  reg  valid_21; // @[DCache.scala 56:22]
  reg  valid_22; // @[DCache.scala 56:22]
  reg  valid_23; // @[DCache.scala 56:22]
  reg  valid_24; // @[DCache.scala 56:22]
  reg  valid_25; // @[DCache.scala 56:22]
  reg  valid_26; // @[DCache.scala 56:22]
  reg  valid_27; // @[DCache.scala 56:22]
  reg  valid_28; // @[DCache.scala 56:22]
  reg  valid_29; // @[DCache.scala 56:22]
  reg  valid_30; // @[DCache.scala 56:22]
  reg  valid_31; // @[DCache.scala 56:22]
  reg  valid_32; // @[DCache.scala 56:22]
  reg  valid_33; // @[DCache.scala 56:22]
  reg  valid_34; // @[DCache.scala 56:22]
  reg  valid_35; // @[DCache.scala 56:22]
  reg  valid_36; // @[DCache.scala 56:22]
  reg  valid_37; // @[DCache.scala 56:22]
  reg  valid_38; // @[DCache.scala 56:22]
  reg  valid_39; // @[DCache.scala 56:22]
  reg  valid_40; // @[DCache.scala 56:22]
  reg  valid_41; // @[DCache.scala 56:22]
  reg  valid_42; // @[DCache.scala 56:22]
  reg  valid_43; // @[DCache.scala 56:22]
  reg  valid_44; // @[DCache.scala 56:22]
  reg  valid_45; // @[DCache.scala 56:22]
  reg  valid_46; // @[DCache.scala 56:22]
  reg  valid_47; // @[DCache.scala 56:22]
  reg  valid_48; // @[DCache.scala 56:22]
  reg  valid_49; // @[DCache.scala 56:22]
  reg  valid_50; // @[DCache.scala 56:22]
  reg  valid_51; // @[DCache.scala 56:22]
  reg  valid_52; // @[DCache.scala 56:22]
  reg  valid_53; // @[DCache.scala 56:22]
  reg  valid_54; // @[DCache.scala 56:22]
  reg  valid_55; // @[DCache.scala 56:22]
  reg  valid_56; // @[DCache.scala 56:22]
  reg  valid_57; // @[DCache.scala 56:22]
  reg  valid_58; // @[DCache.scala 56:22]
  reg  valid_59; // @[DCache.scala 56:22]
  reg  valid_60; // @[DCache.scala 56:22]
  reg  valid_61; // @[DCache.scala 56:22]
  reg  valid_62; // @[DCache.scala 56:22]
  reg  valid_63; // @[DCache.scala 56:22]
  reg  valid_64; // @[DCache.scala 56:22]
  reg  valid_65; // @[DCache.scala 56:22]
  reg  valid_66; // @[DCache.scala 56:22]
  reg  valid_67; // @[DCache.scala 56:22]
  reg  valid_68; // @[DCache.scala 56:22]
  reg  valid_69; // @[DCache.scala 56:22]
  reg  valid_70; // @[DCache.scala 56:22]
  reg  valid_71; // @[DCache.scala 56:22]
  reg  valid_72; // @[DCache.scala 56:22]
  reg  valid_73; // @[DCache.scala 56:22]
  reg  valid_74; // @[DCache.scala 56:22]
  reg  valid_75; // @[DCache.scala 56:22]
  reg  valid_76; // @[DCache.scala 56:22]
  reg  valid_77; // @[DCache.scala 56:22]
  reg  valid_78; // @[DCache.scala 56:22]
  reg  valid_79; // @[DCache.scala 56:22]
  reg  valid_80; // @[DCache.scala 56:22]
  reg  valid_81; // @[DCache.scala 56:22]
  reg  valid_82; // @[DCache.scala 56:22]
  reg  valid_83; // @[DCache.scala 56:22]
  reg  valid_84; // @[DCache.scala 56:22]
  reg  valid_85; // @[DCache.scala 56:22]
  reg  valid_86; // @[DCache.scala 56:22]
  reg  valid_87; // @[DCache.scala 56:22]
  reg  valid_88; // @[DCache.scala 56:22]
  reg  valid_89; // @[DCache.scala 56:22]
  reg  valid_90; // @[DCache.scala 56:22]
  reg  valid_91; // @[DCache.scala 56:22]
  reg  valid_92; // @[DCache.scala 56:22]
  reg  valid_93; // @[DCache.scala 56:22]
  reg  valid_94; // @[DCache.scala 56:22]
  reg  valid_95; // @[DCache.scala 56:22]
  reg  valid_96; // @[DCache.scala 56:22]
  reg  valid_97; // @[DCache.scala 56:22]
  reg  valid_98; // @[DCache.scala 56:22]
  reg  valid_99; // @[DCache.scala 56:22]
  reg  valid_100; // @[DCache.scala 56:22]
  reg  valid_101; // @[DCache.scala 56:22]
  reg  valid_102; // @[DCache.scala 56:22]
  reg  valid_103; // @[DCache.scala 56:22]
  reg  valid_104; // @[DCache.scala 56:22]
  reg  valid_105; // @[DCache.scala 56:22]
  reg  valid_106; // @[DCache.scala 56:22]
  reg  valid_107; // @[DCache.scala 56:22]
  reg  valid_108; // @[DCache.scala 56:22]
  reg  valid_109; // @[DCache.scala 56:22]
  reg  valid_110; // @[DCache.scala 56:22]
  reg  valid_111; // @[DCache.scala 56:22]
  reg  valid_112; // @[DCache.scala 56:22]
  reg  valid_113; // @[DCache.scala 56:22]
  reg  valid_114; // @[DCache.scala 56:22]
  reg  valid_115; // @[DCache.scala 56:22]
  reg  valid_116; // @[DCache.scala 56:22]
  reg  valid_117; // @[DCache.scala 56:22]
  reg  valid_118; // @[DCache.scala 56:22]
  reg  valid_119; // @[DCache.scala 56:22]
  reg  valid_120; // @[DCache.scala 56:22]
  reg  valid_121; // @[DCache.scala 56:22]
  reg  valid_122; // @[DCache.scala 56:22]
  reg  valid_123; // @[DCache.scala 56:22]
  reg  valid_124; // @[DCache.scala 56:22]
  reg  valid_125; // @[DCache.scala 56:22]
  reg  valid_126; // @[DCache.scala 56:22]
  reg  valid_127; // @[DCache.scala 56:22]
  reg  valid_128; // @[DCache.scala 56:22]
  reg  valid_129; // @[DCache.scala 56:22]
  reg  valid_130; // @[DCache.scala 56:22]
  reg  valid_131; // @[DCache.scala 56:22]
  reg  valid_132; // @[DCache.scala 56:22]
  reg  valid_133; // @[DCache.scala 56:22]
  reg  valid_134; // @[DCache.scala 56:22]
  reg  valid_135; // @[DCache.scala 56:22]
  reg  valid_136; // @[DCache.scala 56:22]
  reg  valid_137; // @[DCache.scala 56:22]
  reg  valid_138; // @[DCache.scala 56:22]
  reg  valid_139; // @[DCache.scala 56:22]
  reg  valid_140; // @[DCache.scala 56:22]
  reg  valid_141; // @[DCache.scala 56:22]
  reg  valid_142; // @[DCache.scala 56:22]
  reg  valid_143; // @[DCache.scala 56:22]
  reg  valid_144; // @[DCache.scala 56:22]
  reg  valid_145; // @[DCache.scala 56:22]
  reg  valid_146; // @[DCache.scala 56:22]
  reg  valid_147; // @[DCache.scala 56:22]
  reg  valid_148; // @[DCache.scala 56:22]
  reg  valid_149; // @[DCache.scala 56:22]
  reg  valid_150; // @[DCache.scala 56:22]
  reg  valid_151; // @[DCache.scala 56:22]
  reg  valid_152; // @[DCache.scala 56:22]
  reg  valid_153; // @[DCache.scala 56:22]
  reg  valid_154; // @[DCache.scala 56:22]
  reg  valid_155; // @[DCache.scala 56:22]
  reg  valid_156; // @[DCache.scala 56:22]
  reg  valid_157; // @[DCache.scala 56:22]
  reg  valid_158; // @[DCache.scala 56:22]
  reg  valid_159; // @[DCache.scala 56:22]
  reg  valid_160; // @[DCache.scala 56:22]
  reg  valid_161; // @[DCache.scala 56:22]
  reg  valid_162; // @[DCache.scala 56:22]
  reg  valid_163; // @[DCache.scala 56:22]
  reg  valid_164; // @[DCache.scala 56:22]
  reg  valid_165; // @[DCache.scala 56:22]
  reg  valid_166; // @[DCache.scala 56:22]
  reg  valid_167; // @[DCache.scala 56:22]
  reg  valid_168; // @[DCache.scala 56:22]
  reg  valid_169; // @[DCache.scala 56:22]
  reg  valid_170; // @[DCache.scala 56:22]
  reg  valid_171; // @[DCache.scala 56:22]
  reg  valid_172; // @[DCache.scala 56:22]
  reg  valid_173; // @[DCache.scala 56:22]
  reg  valid_174; // @[DCache.scala 56:22]
  reg  valid_175; // @[DCache.scala 56:22]
  reg  valid_176; // @[DCache.scala 56:22]
  reg  valid_177; // @[DCache.scala 56:22]
  reg  valid_178; // @[DCache.scala 56:22]
  reg  valid_179; // @[DCache.scala 56:22]
  reg  valid_180; // @[DCache.scala 56:22]
  reg  valid_181; // @[DCache.scala 56:22]
  reg  valid_182; // @[DCache.scala 56:22]
  reg  valid_183; // @[DCache.scala 56:22]
  reg  valid_184; // @[DCache.scala 56:22]
  reg  valid_185; // @[DCache.scala 56:22]
  reg  valid_186; // @[DCache.scala 56:22]
  reg  valid_187; // @[DCache.scala 56:22]
  reg  valid_188; // @[DCache.scala 56:22]
  reg  valid_189; // @[DCache.scala 56:22]
  reg  valid_190; // @[DCache.scala 56:22]
  reg  valid_191; // @[DCache.scala 56:22]
  reg  valid_192; // @[DCache.scala 56:22]
  reg  valid_193; // @[DCache.scala 56:22]
  reg  valid_194; // @[DCache.scala 56:22]
  reg  valid_195; // @[DCache.scala 56:22]
  reg  valid_196; // @[DCache.scala 56:22]
  reg  valid_197; // @[DCache.scala 56:22]
  reg  valid_198; // @[DCache.scala 56:22]
  reg  valid_199; // @[DCache.scala 56:22]
  reg  valid_200; // @[DCache.scala 56:22]
  reg  valid_201; // @[DCache.scala 56:22]
  reg  valid_202; // @[DCache.scala 56:22]
  reg  valid_203; // @[DCache.scala 56:22]
  reg  valid_204; // @[DCache.scala 56:22]
  reg  valid_205; // @[DCache.scala 56:22]
  reg  valid_206; // @[DCache.scala 56:22]
  reg  valid_207; // @[DCache.scala 56:22]
  reg  valid_208; // @[DCache.scala 56:22]
  reg  valid_209; // @[DCache.scala 56:22]
  reg  valid_210; // @[DCache.scala 56:22]
  reg  valid_211; // @[DCache.scala 56:22]
  reg  valid_212; // @[DCache.scala 56:22]
  reg  valid_213; // @[DCache.scala 56:22]
  reg  valid_214; // @[DCache.scala 56:22]
  reg  valid_215; // @[DCache.scala 56:22]
  reg  valid_216; // @[DCache.scala 56:22]
  reg  valid_217; // @[DCache.scala 56:22]
  reg  valid_218; // @[DCache.scala 56:22]
  reg  valid_219; // @[DCache.scala 56:22]
  reg  valid_220; // @[DCache.scala 56:22]
  reg  valid_221; // @[DCache.scala 56:22]
  reg  valid_222; // @[DCache.scala 56:22]
  reg  valid_223; // @[DCache.scala 56:22]
  reg  valid_224; // @[DCache.scala 56:22]
  reg  valid_225; // @[DCache.scala 56:22]
  reg  valid_226; // @[DCache.scala 56:22]
  reg  valid_227; // @[DCache.scala 56:22]
  reg  valid_228; // @[DCache.scala 56:22]
  reg  valid_229; // @[DCache.scala 56:22]
  reg  valid_230; // @[DCache.scala 56:22]
  reg  valid_231; // @[DCache.scala 56:22]
  reg  valid_232; // @[DCache.scala 56:22]
  reg  valid_233; // @[DCache.scala 56:22]
  reg  valid_234; // @[DCache.scala 56:22]
  reg  valid_235; // @[DCache.scala 56:22]
  reg  valid_236; // @[DCache.scala 56:22]
  reg  valid_237; // @[DCache.scala 56:22]
  reg  valid_238; // @[DCache.scala 56:22]
  reg  valid_239; // @[DCache.scala 56:22]
  reg  valid_240; // @[DCache.scala 56:22]
  reg  valid_241; // @[DCache.scala 56:22]
  reg  valid_242; // @[DCache.scala 56:22]
  reg  valid_243; // @[DCache.scala 56:22]
  reg  valid_244; // @[DCache.scala 56:22]
  reg  valid_245; // @[DCache.scala 56:22]
  reg  valid_246; // @[DCache.scala 56:22]
  reg  valid_247; // @[DCache.scala 56:22]
  reg  valid_248; // @[DCache.scala 56:22]
  reg  valid_249; // @[DCache.scala 56:22]
  reg  valid_250; // @[DCache.scala 56:22]
  reg  valid_251; // @[DCache.scala 56:22]
  reg  valid_252; // @[DCache.scala 56:22]
  reg  valid_253; // @[DCache.scala 56:22]
  reg  valid_254; // @[DCache.scala 56:22]
  reg  valid_255; // @[DCache.scala 56:22]
  reg  valid_256; // @[DCache.scala 56:22]
  reg  valid_257; // @[DCache.scala 56:22]
  reg  valid_258; // @[DCache.scala 56:22]
  reg  valid_259; // @[DCache.scala 56:22]
  reg  valid_260; // @[DCache.scala 56:22]
  reg  valid_261; // @[DCache.scala 56:22]
  reg  valid_262; // @[DCache.scala 56:22]
  reg  valid_263; // @[DCache.scala 56:22]
  reg  valid_264; // @[DCache.scala 56:22]
  reg  valid_265; // @[DCache.scala 56:22]
  reg  valid_266; // @[DCache.scala 56:22]
  reg  valid_267; // @[DCache.scala 56:22]
  reg  valid_268; // @[DCache.scala 56:22]
  reg  valid_269; // @[DCache.scala 56:22]
  reg  valid_270; // @[DCache.scala 56:22]
  reg  valid_271; // @[DCache.scala 56:22]
  reg  valid_272; // @[DCache.scala 56:22]
  reg  valid_273; // @[DCache.scala 56:22]
  reg  valid_274; // @[DCache.scala 56:22]
  reg  valid_275; // @[DCache.scala 56:22]
  reg  valid_276; // @[DCache.scala 56:22]
  reg  valid_277; // @[DCache.scala 56:22]
  reg  valid_278; // @[DCache.scala 56:22]
  reg  valid_279; // @[DCache.scala 56:22]
  reg  valid_280; // @[DCache.scala 56:22]
  reg  valid_281; // @[DCache.scala 56:22]
  reg  valid_282; // @[DCache.scala 56:22]
  reg  valid_283; // @[DCache.scala 56:22]
  reg  valid_284; // @[DCache.scala 56:22]
  reg  valid_285; // @[DCache.scala 56:22]
  reg  valid_286; // @[DCache.scala 56:22]
  reg  valid_287; // @[DCache.scala 56:22]
  reg  valid_288; // @[DCache.scala 56:22]
  reg  valid_289; // @[DCache.scala 56:22]
  reg  valid_290; // @[DCache.scala 56:22]
  reg  valid_291; // @[DCache.scala 56:22]
  reg  valid_292; // @[DCache.scala 56:22]
  reg  valid_293; // @[DCache.scala 56:22]
  reg  valid_294; // @[DCache.scala 56:22]
  reg  valid_295; // @[DCache.scala 56:22]
  reg  valid_296; // @[DCache.scala 56:22]
  reg  valid_297; // @[DCache.scala 56:22]
  reg  valid_298; // @[DCache.scala 56:22]
  reg  valid_299; // @[DCache.scala 56:22]
  reg  valid_300; // @[DCache.scala 56:22]
  reg  valid_301; // @[DCache.scala 56:22]
  reg  valid_302; // @[DCache.scala 56:22]
  reg  valid_303; // @[DCache.scala 56:22]
  reg  valid_304; // @[DCache.scala 56:22]
  reg  valid_305; // @[DCache.scala 56:22]
  reg  valid_306; // @[DCache.scala 56:22]
  reg  valid_307; // @[DCache.scala 56:22]
  reg  valid_308; // @[DCache.scala 56:22]
  reg  valid_309; // @[DCache.scala 56:22]
  reg  valid_310; // @[DCache.scala 56:22]
  reg  valid_311; // @[DCache.scala 56:22]
  reg  valid_312; // @[DCache.scala 56:22]
  reg  valid_313; // @[DCache.scala 56:22]
  reg  valid_314; // @[DCache.scala 56:22]
  reg  valid_315; // @[DCache.scala 56:22]
  reg  valid_316; // @[DCache.scala 56:22]
  reg  valid_317; // @[DCache.scala 56:22]
  reg  valid_318; // @[DCache.scala 56:22]
  reg  valid_319; // @[DCache.scala 56:22]
  reg  valid_320; // @[DCache.scala 56:22]
  reg  valid_321; // @[DCache.scala 56:22]
  reg  valid_322; // @[DCache.scala 56:22]
  reg  valid_323; // @[DCache.scala 56:22]
  reg  valid_324; // @[DCache.scala 56:22]
  reg  valid_325; // @[DCache.scala 56:22]
  reg  valid_326; // @[DCache.scala 56:22]
  reg  valid_327; // @[DCache.scala 56:22]
  reg  valid_328; // @[DCache.scala 56:22]
  reg  valid_329; // @[DCache.scala 56:22]
  reg  valid_330; // @[DCache.scala 56:22]
  reg  valid_331; // @[DCache.scala 56:22]
  reg  valid_332; // @[DCache.scala 56:22]
  reg  valid_333; // @[DCache.scala 56:22]
  reg  valid_334; // @[DCache.scala 56:22]
  reg  valid_335; // @[DCache.scala 56:22]
  reg  valid_336; // @[DCache.scala 56:22]
  reg  valid_337; // @[DCache.scala 56:22]
  reg  valid_338; // @[DCache.scala 56:22]
  reg  valid_339; // @[DCache.scala 56:22]
  reg  valid_340; // @[DCache.scala 56:22]
  reg  valid_341; // @[DCache.scala 56:22]
  reg  valid_342; // @[DCache.scala 56:22]
  reg  valid_343; // @[DCache.scala 56:22]
  reg  valid_344; // @[DCache.scala 56:22]
  reg  valid_345; // @[DCache.scala 56:22]
  reg  valid_346; // @[DCache.scala 56:22]
  reg  valid_347; // @[DCache.scala 56:22]
  reg  valid_348; // @[DCache.scala 56:22]
  reg  valid_349; // @[DCache.scala 56:22]
  reg  valid_350; // @[DCache.scala 56:22]
  reg  valid_351; // @[DCache.scala 56:22]
  reg  valid_352; // @[DCache.scala 56:22]
  reg  valid_353; // @[DCache.scala 56:22]
  reg  valid_354; // @[DCache.scala 56:22]
  reg  valid_355; // @[DCache.scala 56:22]
  reg  valid_356; // @[DCache.scala 56:22]
  reg  valid_357; // @[DCache.scala 56:22]
  reg  valid_358; // @[DCache.scala 56:22]
  reg  valid_359; // @[DCache.scala 56:22]
  reg  valid_360; // @[DCache.scala 56:22]
  reg  valid_361; // @[DCache.scala 56:22]
  reg  valid_362; // @[DCache.scala 56:22]
  reg  valid_363; // @[DCache.scala 56:22]
  reg  valid_364; // @[DCache.scala 56:22]
  reg  valid_365; // @[DCache.scala 56:22]
  reg  valid_366; // @[DCache.scala 56:22]
  reg  valid_367; // @[DCache.scala 56:22]
  reg  valid_368; // @[DCache.scala 56:22]
  reg  valid_369; // @[DCache.scala 56:22]
  reg  valid_370; // @[DCache.scala 56:22]
  reg  valid_371; // @[DCache.scala 56:22]
  reg  valid_372; // @[DCache.scala 56:22]
  reg  valid_373; // @[DCache.scala 56:22]
  reg  valid_374; // @[DCache.scala 56:22]
  reg  valid_375; // @[DCache.scala 56:22]
  reg  valid_376; // @[DCache.scala 56:22]
  reg  valid_377; // @[DCache.scala 56:22]
  reg  valid_378; // @[DCache.scala 56:22]
  reg  valid_379; // @[DCache.scala 56:22]
  reg  valid_380; // @[DCache.scala 56:22]
  reg  valid_381; // @[DCache.scala 56:22]
  reg  valid_382; // @[DCache.scala 56:22]
  reg  valid_383; // @[DCache.scala 56:22]
  reg  valid_384; // @[DCache.scala 56:22]
  reg  valid_385; // @[DCache.scala 56:22]
  reg  valid_386; // @[DCache.scala 56:22]
  reg  valid_387; // @[DCache.scala 56:22]
  reg  valid_388; // @[DCache.scala 56:22]
  reg  valid_389; // @[DCache.scala 56:22]
  reg  valid_390; // @[DCache.scala 56:22]
  reg  valid_391; // @[DCache.scala 56:22]
  reg  valid_392; // @[DCache.scala 56:22]
  reg  valid_393; // @[DCache.scala 56:22]
  reg  valid_394; // @[DCache.scala 56:22]
  reg  valid_395; // @[DCache.scala 56:22]
  reg  valid_396; // @[DCache.scala 56:22]
  reg  valid_397; // @[DCache.scala 56:22]
  reg  valid_398; // @[DCache.scala 56:22]
  reg  valid_399; // @[DCache.scala 56:22]
  reg  valid_400; // @[DCache.scala 56:22]
  reg  valid_401; // @[DCache.scala 56:22]
  reg  valid_402; // @[DCache.scala 56:22]
  reg  valid_403; // @[DCache.scala 56:22]
  reg  valid_404; // @[DCache.scala 56:22]
  reg  valid_405; // @[DCache.scala 56:22]
  reg  valid_406; // @[DCache.scala 56:22]
  reg  valid_407; // @[DCache.scala 56:22]
  reg  valid_408; // @[DCache.scala 56:22]
  reg  valid_409; // @[DCache.scala 56:22]
  reg  valid_410; // @[DCache.scala 56:22]
  reg  valid_411; // @[DCache.scala 56:22]
  reg  valid_412; // @[DCache.scala 56:22]
  reg  valid_413; // @[DCache.scala 56:22]
  reg  valid_414; // @[DCache.scala 56:22]
  reg  valid_415; // @[DCache.scala 56:22]
  reg  valid_416; // @[DCache.scala 56:22]
  reg  valid_417; // @[DCache.scala 56:22]
  reg  valid_418; // @[DCache.scala 56:22]
  reg  valid_419; // @[DCache.scala 56:22]
  reg  valid_420; // @[DCache.scala 56:22]
  reg  valid_421; // @[DCache.scala 56:22]
  reg  valid_422; // @[DCache.scala 56:22]
  reg  valid_423; // @[DCache.scala 56:22]
  reg  valid_424; // @[DCache.scala 56:22]
  reg  valid_425; // @[DCache.scala 56:22]
  reg  valid_426; // @[DCache.scala 56:22]
  reg  valid_427; // @[DCache.scala 56:22]
  reg  valid_428; // @[DCache.scala 56:22]
  reg  valid_429; // @[DCache.scala 56:22]
  reg  valid_430; // @[DCache.scala 56:22]
  reg  valid_431; // @[DCache.scala 56:22]
  reg  valid_432; // @[DCache.scala 56:22]
  reg  valid_433; // @[DCache.scala 56:22]
  reg  valid_434; // @[DCache.scala 56:22]
  reg  valid_435; // @[DCache.scala 56:22]
  reg  valid_436; // @[DCache.scala 56:22]
  reg  valid_437; // @[DCache.scala 56:22]
  reg  valid_438; // @[DCache.scala 56:22]
  reg  valid_439; // @[DCache.scala 56:22]
  reg  valid_440; // @[DCache.scala 56:22]
  reg  valid_441; // @[DCache.scala 56:22]
  reg  valid_442; // @[DCache.scala 56:22]
  reg  valid_443; // @[DCache.scala 56:22]
  reg  valid_444; // @[DCache.scala 56:22]
  reg  valid_445; // @[DCache.scala 56:22]
  reg  valid_446; // @[DCache.scala 56:22]
  reg  valid_447; // @[DCache.scala 56:22]
  reg  valid_448; // @[DCache.scala 56:22]
  reg  valid_449; // @[DCache.scala 56:22]
  reg  valid_450; // @[DCache.scala 56:22]
  reg  valid_451; // @[DCache.scala 56:22]
  reg  valid_452; // @[DCache.scala 56:22]
  reg  valid_453; // @[DCache.scala 56:22]
  reg  valid_454; // @[DCache.scala 56:22]
  reg  valid_455; // @[DCache.scala 56:22]
  reg  valid_456; // @[DCache.scala 56:22]
  reg  valid_457; // @[DCache.scala 56:22]
  reg  valid_458; // @[DCache.scala 56:22]
  reg  valid_459; // @[DCache.scala 56:22]
  reg  valid_460; // @[DCache.scala 56:22]
  reg  valid_461; // @[DCache.scala 56:22]
  reg  valid_462; // @[DCache.scala 56:22]
  reg  valid_463; // @[DCache.scala 56:22]
  reg  valid_464; // @[DCache.scala 56:22]
  reg  valid_465; // @[DCache.scala 56:22]
  reg  valid_466; // @[DCache.scala 56:22]
  reg  valid_467; // @[DCache.scala 56:22]
  reg  valid_468; // @[DCache.scala 56:22]
  reg  valid_469; // @[DCache.scala 56:22]
  reg  valid_470; // @[DCache.scala 56:22]
  reg  valid_471; // @[DCache.scala 56:22]
  reg  valid_472; // @[DCache.scala 56:22]
  reg  valid_473; // @[DCache.scala 56:22]
  reg  valid_474; // @[DCache.scala 56:22]
  reg  valid_475; // @[DCache.scala 56:22]
  reg  valid_476; // @[DCache.scala 56:22]
  reg  valid_477; // @[DCache.scala 56:22]
  reg  valid_478; // @[DCache.scala 56:22]
  reg  valid_479; // @[DCache.scala 56:22]
  reg  valid_480; // @[DCache.scala 56:22]
  reg  valid_481; // @[DCache.scala 56:22]
  reg  valid_482; // @[DCache.scala 56:22]
  reg  valid_483; // @[DCache.scala 56:22]
  reg  valid_484; // @[DCache.scala 56:22]
  reg  valid_485; // @[DCache.scala 56:22]
  reg  valid_486; // @[DCache.scala 56:22]
  reg  valid_487; // @[DCache.scala 56:22]
  reg  valid_488; // @[DCache.scala 56:22]
  reg  valid_489; // @[DCache.scala 56:22]
  reg  valid_490; // @[DCache.scala 56:22]
  reg  valid_491; // @[DCache.scala 56:22]
  reg  valid_492; // @[DCache.scala 56:22]
  reg  valid_493; // @[DCache.scala 56:22]
  reg  valid_494; // @[DCache.scala 56:22]
  reg  valid_495; // @[DCache.scala 56:22]
  reg  valid_496; // @[DCache.scala 56:22]
  reg  valid_497; // @[DCache.scala 56:22]
  reg  valid_498; // @[DCache.scala 56:22]
  reg  valid_499; // @[DCache.scala 56:22]
  reg  valid_500; // @[DCache.scala 56:22]
  reg  valid_501; // @[DCache.scala 56:22]
  reg  valid_502; // @[DCache.scala 56:22]
  reg  valid_503; // @[DCache.scala 56:22]
  reg  valid_504; // @[DCache.scala 56:22]
  reg  valid_505; // @[DCache.scala 56:22]
  reg  valid_506; // @[DCache.scala 56:22]
  reg  valid_507; // @[DCache.scala 56:22]
  reg  valid_508; // @[DCache.scala 56:22]
  reg  valid_509; // @[DCache.scala 56:22]
  reg  valid_510; // @[DCache.scala 56:22]
  reg  valid_511; // @[DCache.scala 56:22]
  wire [31:0] array_addr = _GEN_16[31:0]; // @[DCache.scala 63:24 64:14]
  wire [17:0] array_wdata_tag = array_addr[31:14]; // @[DCache.scala 53:29]
  wire  _array_io_en_T_1 = io_cache_resp_ready & io_cache_resp_valid; // @[Decoupled.scala 51:35]
  wire  _T_11 = state == 3'h7; // @[DCache.scala 165:16]
  wire  amo_w = req_r_len == 2'h2; // @[DCache.scala 98:37]
  wire [31:0] _amo_wdata_raw_64_T_4 = req_r_addr[2] ? req_r_wdata[63:32] : req_r_wdata[31:0]; // @[DCache.scala 106:21]
  wire [31:0] _amo_wdata_raw_64_T_7 = _amo_wdata_raw_64_T_4[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _amo_wdata_raw_64_T_8 = {_amo_wdata_raw_64_T_7,_amo_wdata_raw_64_T_4}; // @[Cat.scala 33:92]
  wire [63:0] amo_wdata_raw_64 = amo_w ? _amo_wdata_raw_64_T_8 : req_r_wdata; // @[DCache.scala 104:26]
  reg  array_out_REG; // @[DCache.scala 76:55]
  reg [273:0] array_out_r; // @[Reg.scala 35:20]
  wire [273:0] _array_out_T_1 = array_out_REG ? array_io_rdata : array_out_r; // @[Utils.scala 50:8]
  wire [255:0] array_out_data = _array_out_T_1[255:0]; // @[DCache.scala 76:75]
  wire [255:0] rdata_256 = _T_11 ? tl_d_bits_r_data : array_out_data; // @[DCache.scala 81:22]
  wire [63:0] _rdata_64_T_6 = 2'h1 == array_addr[4:3] ? rdata_256[127:64] : rdata_256[63:0]; // @[Mux.scala 81:58]
  wire [63:0] _rdata_64_T_8 = 2'h2 == array_addr[4:3] ? rdata_256[191:128] : _rdata_64_T_6; // @[Mux.scala 81:58]
  wire [63:0] rdata_64 = 2'h3 == array_addr[4:3] ? rdata_256[255:192] : _rdata_64_T_8; // @[Mux.scala 81:58]
  wire [31:0] _amo_rdata_raw_64_T_4 = req_r_addr[2] ? rdata_64[63:32] : rdata_64[31:0]; // @[DCache.scala 101:21]
  wire [31:0] _amo_rdata_raw_64_T_7 = _amo_rdata_raw_64_T_4[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _amo_rdata_raw_64_T_8 = {_amo_rdata_raw_64_T_7,_amo_rdata_raw_64_T_4}; // @[Cat.scala 33:92]
  wire [63:0] amo_rdata_raw_64 = amo_w ? _amo_rdata_raw_64_T_8 : rdata_64; // @[DCache.scala 99:26]
  wire [63:0] _amo_result_64_T_16 = amo_wdata_raw_64 < amo_rdata_raw_64 ? amo_wdata_raw_64 : amo_rdata_raw_64; // @[DCache.scala 121:32]
  wire [63:0] _amo_result_64_T_11 = amo_w ? _amo_wdata_raw_64_T_8 : req_r_wdata; // @[DCache.scala 120:50]
  wire [63:0] _amo_result_64_T_12 = amo_w ? _amo_rdata_raw_64_T_8 : rdata_64; // @[DCache.scala 120:76]
  wire [63:0] _amo_result_64_T_14 = $signed(_amo_result_64_T_11) < $signed(_amo_result_64_T_12) ? amo_wdata_raw_64 :
    amo_rdata_raw_64; // @[DCache.scala 120:32]
  wire [63:0] _amo_result_64_T_10 = amo_wdata_raw_64 > amo_rdata_raw_64 ? amo_wdata_raw_64 : amo_rdata_raw_64; // @[DCache.scala 119:32]
  wire [63:0] _amo_result_64_T_8 = $signed(_amo_result_64_T_11) > $signed(_amo_result_64_T_12) ? amo_wdata_raw_64 :
    amo_rdata_raw_64; // @[DCache.scala 118:32]
  wire [63:0] _amo_result_64_T_4 = amo_wdata_raw_64 ^ amo_rdata_raw_64; // @[DCache.scala 117:47]
  wire [63:0] _amo_result_64_T_3 = amo_wdata_raw_64 | amo_rdata_raw_64; // @[DCache.scala 116:47]
  wire [63:0] _amo_result_64_T_2 = amo_wdata_raw_64 & amo_rdata_raw_64; // @[DCache.scala 115:47]
  wire [63:0] _amo_result_64_T_1 = amo_wdata_raw_64 + amo_rdata_raw_64; // @[DCache.scala 114:47]
  wire [63:0] _amo_result_64_T_18 = 5'h1b == req_r_amo ? amo_wdata_raw_64 : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _amo_result_64_T_20 = 5'h14 == req_r_amo ? _amo_result_64_T_1 : _amo_result_64_T_18; // @[Mux.scala 81:58]
  wire [63:0] _amo_result_64_T_22 = 5'h1a == req_r_amo ? _amo_result_64_T_2 : _amo_result_64_T_20; // @[Mux.scala 81:58]
  wire [63:0] _amo_result_64_T_24 = 5'h19 == req_r_amo ? _amo_result_64_T_3 : _amo_result_64_T_22; // @[Mux.scala 81:58]
  wire [63:0] _amo_result_64_T_26 = 5'h18 == req_r_amo ? _amo_result_64_T_4 : _amo_result_64_T_24; // @[Mux.scala 81:58]
  wire [63:0] _amo_result_64_T_28 = 5'h11 == req_r_amo ? _amo_result_64_T_8 : _amo_result_64_T_26; // @[Mux.scala 81:58]
  wire [63:0] _amo_result_64_T_30 = 5'h13 == req_r_amo ? _amo_result_64_T_10 : _amo_result_64_T_28; // @[Mux.scala 81:58]
  wire [63:0] _amo_result_64_T_32 = 5'h10 == req_r_amo ? _amo_result_64_T_14 : _amo_result_64_T_30; // @[Mux.scala 81:58]
  wire [63:0] amo_result_64 = 5'h12 == req_r_amo ? _amo_result_64_T_16 : _amo_result_64_T_32; // @[Mux.scala 81:58]
  wire [63:0] _amo_wdata_64_T_4 = {amo_result_64[31:0],32'h0}; // @[Cat.scala 33:92]
  wire [63:0] amo_wdata_64 = amo_w & req_r_addr[2] ? _amo_wdata_64_T_4 : amo_result_64; // @[DCache.scala 124:22]
  wire [63:0] wdata_64 = req_r_amo[4] ? amo_wdata_64 : req_r_wdata; // @[DCache.scala 157:22]
  wire [7:0] _wdata_256_T_1 = {req_r_addr[4:3], 6'h0}; // @[DCache.scala 160:51]
  wire [318:0] _GEN_0 = {{255'd0}, wdata_64}; // @[DCache.scala 160:25]
  wire [318:0] _wdata_256_T_2 = _GEN_0 << _wdata_256_T_1; // @[DCache.scala 160:25]
  wire [255:0] wdata_256 = _wdata_256_T_2[255:0]; // @[DCache.scala 158:23 160:13]
  wire [7:0] _wmask_256_T_23 = req_r_wmask[7] ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _wmask_256_T_21 = req_r_wmask[6] ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _wmask_256_T_19 = req_r_wmask[5] ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _wmask_256_T_17 = req_r_wmask[4] ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _wmask_256_T_15 = req_r_wmask[3] ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _wmask_256_T_13 = req_r_wmask[2] ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _wmask_256_T_11 = req_r_wmask[1] ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _wmask_256_T_9 = req_r_wmask[0] ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _wmask_256_T_24 = {_wmask_256_T_23,_wmask_256_T_21,_wmask_256_T_19,_wmask_256_T_17,_wmask_256_T_15,
    _wmask_256_T_13,_wmask_256_T_11,_wmask_256_T_9}; // @[Cat.scala 33:92]
  wire [318:0] _GEN_1 = {{255'd0}, _wmask_256_T_24}; // @[DCache.scala 161:40]
  wire [318:0] _wmask_256_T_27 = _GEN_1 << _wdata_256_T_1; // @[DCache.scala 161:40]
  wire [255:0] wmask_256 = _wmask_256_T_27[255:0]; // @[DCache.scala 159:23 161:13]
  wire [255:0] _array_wdata_data_T = wdata_256 & wmask_256; // @[Utils.scala 18:15]
  wire [255:0] _array_wdata_data_T_1 = ~wmask_256; // @[Utils.scala 18:38]
  wire [255:0] _array_wdata_data_T_2 = tl_d_bits_r_data & _array_wdata_data_T_1; // @[Utils.scala 18:35]
  wire [255:0] _array_wdata_data_T_3 = _array_wdata_data_T | _array_wdata_data_T_2; // @[Utils.scala 18:23]
  wire [255:0] _array_wdata_data_T_4 = req_r_wen ? _array_wdata_data_T_3 : tl_d_bits_r_data; // @[DCache.scala 166:30]
  wire [255:0] _array_wdata_data_T_7 = array_out_data & _array_wdata_data_T_1; // @[Utils.scala 18:35]
  wire [255:0] _array_wdata_data_T_8 = _array_wdata_data_T | _array_wdata_data_T_7; // @[Utils.scala 18:23]
  wire [255:0] _GEN_1570 = state == 3'h7 ? _array_wdata_data_T_4 : _array_wdata_data_T_8; // @[DCache.scala 165:26 166:24 176:24]
  wire [255:0] array_wdata_data = _array_io_en_T_1 ? _GEN_1570 : 256'h0; // @[DCache.scala 164:19 69:20]
  wire [17:0] array_out_tag = _array_out_T_1[273:256]; // @[DCache.scala 76:75]
  wire  _GEN_25 = 9'h1 == array_addr[13:5] ? valid_1 : valid_0; // @[DCache.scala 78:{33,33}]
  wire  _GEN_26 = 9'h2 == array_addr[13:5] ? valid_2 : _GEN_25; // @[DCache.scala 78:{33,33}]
  wire  _GEN_27 = 9'h3 == array_addr[13:5] ? valid_3 : _GEN_26; // @[DCache.scala 78:{33,33}]
  wire  _GEN_28 = 9'h4 == array_addr[13:5] ? valid_4 : _GEN_27; // @[DCache.scala 78:{33,33}]
  wire  _GEN_29 = 9'h5 == array_addr[13:5] ? valid_5 : _GEN_28; // @[DCache.scala 78:{33,33}]
  wire  _GEN_30 = 9'h6 == array_addr[13:5] ? valid_6 : _GEN_29; // @[DCache.scala 78:{33,33}]
  wire  _GEN_31 = 9'h7 == array_addr[13:5] ? valid_7 : _GEN_30; // @[DCache.scala 78:{33,33}]
  wire  _GEN_32 = 9'h8 == array_addr[13:5] ? valid_8 : _GEN_31; // @[DCache.scala 78:{33,33}]
  wire  _GEN_33 = 9'h9 == array_addr[13:5] ? valid_9 : _GEN_32; // @[DCache.scala 78:{33,33}]
  wire  _GEN_34 = 9'ha == array_addr[13:5] ? valid_10 : _GEN_33; // @[DCache.scala 78:{33,33}]
  wire  _GEN_35 = 9'hb == array_addr[13:5] ? valid_11 : _GEN_34; // @[DCache.scala 78:{33,33}]
  wire  _GEN_36 = 9'hc == array_addr[13:5] ? valid_12 : _GEN_35; // @[DCache.scala 78:{33,33}]
  wire  _GEN_37 = 9'hd == array_addr[13:5] ? valid_13 : _GEN_36; // @[DCache.scala 78:{33,33}]
  wire  _GEN_38 = 9'he == array_addr[13:5] ? valid_14 : _GEN_37; // @[DCache.scala 78:{33,33}]
  wire  _GEN_39 = 9'hf == array_addr[13:5] ? valid_15 : _GEN_38; // @[DCache.scala 78:{33,33}]
  wire  _GEN_40 = 9'h10 == array_addr[13:5] ? valid_16 : _GEN_39; // @[DCache.scala 78:{33,33}]
  wire  _GEN_41 = 9'h11 == array_addr[13:5] ? valid_17 : _GEN_40; // @[DCache.scala 78:{33,33}]
  wire  _GEN_42 = 9'h12 == array_addr[13:5] ? valid_18 : _GEN_41; // @[DCache.scala 78:{33,33}]
  wire  _GEN_43 = 9'h13 == array_addr[13:5] ? valid_19 : _GEN_42; // @[DCache.scala 78:{33,33}]
  wire  _GEN_44 = 9'h14 == array_addr[13:5] ? valid_20 : _GEN_43; // @[DCache.scala 78:{33,33}]
  wire  _GEN_45 = 9'h15 == array_addr[13:5] ? valid_21 : _GEN_44; // @[DCache.scala 78:{33,33}]
  wire  _GEN_46 = 9'h16 == array_addr[13:5] ? valid_22 : _GEN_45; // @[DCache.scala 78:{33,33}]
  wire  _GEN_47 = 9'h17 == array_addr[13:5] ? valid_23 : _GEN_46; // @[DCache.scala 78:{33,33}]
  wire  _GEN_48 = 9'h18 == array_addr[13:5] ? valid_24 : _GEN_47; // @[DCache.scala 78:{33,33}]
  wire  _GEN_49 = 9'h19 == array_addr[13:5] ? valid_25 : _GEN_48; // @[DCache.scala 78:{33,33}]
  wire  _GEN_50 = 9'h1a == array_addr[13:5] ? valid_26 : _GEN_49; // @[DCache.scala 78:{33,33}]
  wire  _GEN_51 = 9'h1b == array_addr[13:5] ? valid_27 : _GEN_50; // @[DCache.scala 78:{33,33}]
  wire  _GEN_52 = 9'h1c == array_addr[13:5] ? valid_28 : _GEN_51; // @[DCache.scala 78:{33,33}]
  wire  _GEN_53 = 9'h1d == array_addr[13:5] ? valid_29 : _GEN_52; // @[DCache.scala 78:{33,33}]
  wire  _GEN_54 = 9'h1e == array_addr[13:5] ? valid_30 : _GEN_53; // @[DCache.scala 78:{33,33}]
  wire  _GEN_55 = 9'h1f == array_addr[13:5] ? valid_31 : _GEN_54; // @[DCache.scala 78:{33,33}]
  wire  _GEN_56 = 9'h20 == array_addr[13:5] ? valid_32 : _GEN_55; // @[DCache.scala 78:{33,33}]
  wire  _GEN_57 = 9'h21 == array_addr[13:5] ? valid_33 : _GEN_56; // @[DCache.scala 78:{33,33}]
  wire  _GEN_58 = 9'h22 == array_addr[13:5] ? valid_34 : _GEN_57; // @[DCache.scala 78:{33,33}]
  wire  _GEN_59 = 9'h23 == array_addr[13:5] ? valid_35 : _GEN_58; // @[DCache.scala 78:{33,33}]
  wire  _GEN_60 = 9'h24 == array_addr[13:5] ? valid_36 : _GEN_59; // @[DCache.scala 78:{33,33}]
  wire  _GEN_61 = 9'h25 == array_addr[13:5] ? valid_37 : _GEN_60; // @[DCache.scala 78:{33,33}]
  wire  _GEN_62 = 9'h26 == array_addr[13:5] ? valid_38 : _GEN_61; // @[DCache.scala 78:{33,33}]
  wire  _GEN_63 = 9'h27 == array_addr[13:5] ? valid_39 : _GEN_62; // @[DCache.scala 78:{33,33}]
  wire  _GEN_64 = 9'h28 == array_addr[13:5] ? valid_40 : _GEN_63; // @[DCache.scala 78:{33,33}]
  wire  _GEN_65 = 9'h29 == array_addr[13:5] ? valid_41 : _GEN_64; // @[DCache.scala 78:{33,33}]
  wire  _GEN_66 = 9'h2a == array_addr[13:5] ? valid_42 : _GEN_65; // @[DCache.scala 78:{33,33}]
  wire  _GEN_67 = 9'h2b == array_addr[13:5] ? valid_43 : _GEN_66; // @[DCache.scala 78:{33,33}]
  wire  _GEN_68 = 9'h2c == array_addr[13:5] ? valid_44 : _GEN_67; // @[DCache.scala 78:{33,33}]
  wire  _GEN_69 = 9'h2d == array_addr[13:5] ? valid_45 : _GEN_68; // @[DCache.scala 78:{33,33}]
  wire  _GEN_70 = 9'h2e == array_addr[13:5] ? valid_46 : _GEN_69; // @[DCache.scala 78:{33,33}]
  wire  _GEN_71 = 9'h2f == array_addr[13:5] ? valid_47 : _GEN_70; // @[DCache.scala 78:{33,33}]
  wire  _GEN_72 = 9'h30 == array_addr[13:5] ? valid_48 : _GEN_71; // @[DCache.scala 78:{33,33}]
  wire  _GEN_73 = 9'h31 == array_addr[13:5] ? valid_49 : _GEN_72; // @[DCache.scala 78:{33,33}]
  wire  _GEN_74 = 9'h32 == array_addr[13:5] ? valid_50 : _GEN_73; // @[DCache.scala 78:{33,33}]
  wire  _GEN_75 = 9'h33 == array_addr[13:5] ? valid_51 : _GEN_74; // @[DCache.scala 78:{33,33}]
  wire  _GEN_76 = 9'h34 == array_addr[13:5] ? valid_52 : _GEN_75; // @[DCache.scala 78:{33,33}]
  wire  _GEN_77 = 9'h35 == array_addr[13:5] ? valid_53 : _GEN_76; // @[DCache.scala 78:{33,33}]
  wire  _GEN_78 = 9'h36 == array_addr[13:5] ? valid_54 : _GEN_77; // @[DCache.scala 78:{33,33}]
  wire  _GEN_79 = 9'h37 == array_addr[13:5] ? valid_55 : _GEN_78; // @[DCache.scala 78:{33,33}]
  wire  _GEN_80 = 9'h38 == array_addr[13:5] ? valid_56 : _GEN_79; // @[DCache.scala 78:{33,33}]
  wire  _GEN_81 = 9'h39 == array_addr[13:5] ? valid_57 : _GEN_80; // @[DCache.scala 78:{33,33}]
  wire  _GEN_82 = 9'h3a == array_addr[13:5] ? valid_58 : _GEN_81; // @[DCache.scala 78:{33,33}]
  wire  _GEN_83 = 9'h3b == array_addr[13:5] ? valid_59 : _GEN_82; // @[DCache.scala 78:{33,33}]
  wire  _GEN_84 = 9'h3c == array_addr[13:5] ? valid_60 : _GEN_83; // @[DCache.scala 78:{33,33}]
  wire  _GEN_85 = 9'h3d == array_addr[13:5] ? valid_61 : _GEN_84; // @[DCache.scala 78:{33,33}]
  wire  _GEN_86 = 9'h3e == array_addr[13:5] ? valid_62 : _GEN_85; // @[DCache.scala 78:{33,33}]
  wire  _GEN_87 = 9'h3f == array_addr[13:5] ? valid_63 : _GEN_86; // @[DCache.scala 78:{33,33}]
  wire  _GEN_88 = 9'h40 == array_addr[13:5] ? valid_64 : _GEN_87; // @[DCache.scala 78:{33,33}]
  wire  _GEN_89 = 9'h41 == array_addr[13:5] ? valid_65 : _GEN_88; // @[DCache.scala 78:{33,33}]
  wire  _GEN_90 = 9'h42 == array_addr[13:5] ? valid_66 : _GEN_89; // @[DCache.scala 78:{33,33}]
  wire  _GEN_91 = 9'h43 == array_addr[13:5] ? valid_67 : _GEN_90; // @[DCache.scala 78:{33,33}]
  wire  _GEN_92 = 9'h44 == array_addr[13:5] ? valid_68 : _GEN_91; // @[DCache.scala 78:{33,33}]
  wire  _GEN_93 = 9'h45 == array_addr[13:5] ? valid_69 : _GEN_92; // @[DCache.scala 78:{33,33}]
  wire  _GEN_94 = 9'h46 == array_addr[13:5] ? valid_70 : _GEN_93; // @[DCache.scala 78:{33,33}]
  wire  _GEN_95 = 9'h47 == array_addr[13:5] ? valid_71 : _GEN_94; // @[DCache.scala 78:{33,33}]
  wire  _GEN_96 = 9'h48 == array_addr[13:5] ? valid_72 : _GEN_95; // @[DCache.scala 78:{33,33}]
  wire  _GEN_97 = 9'h49 == array_addr[13:5] ? valid_73 : _GEN_96; // @[DCache.scala 78:{33,33}]
  wire  _GEN_98 = 9'h4a == array_addr[13:5] ? valid_74 : _GEN_97; // @[DCache.scala 78:{33,33}]
  wire  _GEN_99 = 9'h4b == array_addr[13:5] ? valid_75 : _GEN_98; // @[DCache.scala 78:{33,33}]
  wire  _GEN_100 = 9'h4c == array_addr[13:5] ? valid_76 : _GEN_99; // @[DCache.scala 78:{33,33}]
  wire  _GEN_101 = 9'h4d == array_addr[13:5] ? valid_77 : _GEN_100; // @[DCache.scala 78:{33,33}]
  wire  _GEN_102 = 9'h4e == array_addr[13:5] ? valid_78 : _GEN_101; // @[DCache.scala 78:{33,33}]
  wire  _GEN_103 = 9'h4f == array_addr[13:5] ? valid_79 : _GEN_102; // @[DCache.scala 78:{33,33}]
  wire  _GEN_104 = 9'h50 == array_addr[13:5] ? valid_80 : _GEN_103; // @[DCache.scala 78:{33,33}]
  wire  _GEN_105 = 9'h51 == array_addr[13:5] ? valid_81 : _GEN_104; // @[DCache.scala 78:{33,33}]
  wire  _GEN_106 = 9'h52 == array_addr[13:5] ? valid_82 : _GEN_105; // @[DCache.scala 78:{33,33}]
  wire  _GEN_107 = 9'h53 == array_addr[13:5] ? valid_83 : _GEN_106; // @[DCache.scala 78:{33,33}]
  wire  _GEN_108 = 9'h54 == array_addr[13:5] ? valid_84 : _GEN_107; // @[DCache.scala 78:{33,33}]
  wire  _GEN_109 = 9'h55 == array_addr[13:5] ? valid_85 : _GEN_108; // @[DCache.scala 78:{33,33}]
  wire  _GEN_110 = 9'h56 == array_addr[13:5] ? valid_86 : _GEN_109; // @[DCache.scala 78:{33,33}]
  wire  _GEN_111 = 9'h57 == array_addr[13:5] ? valid_87 : _GEN_110; // @[DCache.scala 78:{33,33}]
  wire  _GEN_112 = 9'h58 == array_addr[13:5] ? valid_88 : _GEN_111; // @[DCache.scala 78:{33,33}]
  wire  _GEN_113 = 9'h59 == array_addr[13:5] ? valid_89 : _GEN_112; // @[DCache.scala 78:{33,33}]
  wire  _GEN_114 = 9'h5a == array_addr[13:5] ? valid_90 : _GEN_113; // @[DCache.scala 78:{33,33}]
  wire  _GEN_115 = 9'h5b == array_addr[13:5] ? valid_91 : _GEN_114; // @[DCache.scala 78:{33,33}]
  wire  _GEN_116 = 9'h5c == array_addr[13:5] ? valid_92 : _GEN_115; // @[DCache.scala 78:{33,33}]
  wire  _GEN_117 = 9'h5d == array_addr[13:5] ? valid_93 : _GEN_116; // @[DCache.scala 78:{33,33}]
  wire  _GEN_118 = 9'h5e == array_addr[13:5] ? valid_94 : _GEN_117; // @[DCache.scala 78:{33,33}]
  wire  _GEN_119 = 9'h5f == array_addr[13:5] ? valid_95 : _GEN_118; // @[DCache.scala 78:{33,33}]
  wire  _GEN_120 = 9'h60 == array_addr[13:5] ? valid_96 : _GEN_119; // @[DCache.scala 78:{33,33}]
  wire  _GEN_121 = 9'h61 == array_addr[13:5] ? valid_97 : _GEN_120; // @[DCache.scala 78:{33,33}]
  wire  _GEN_122 = 9'h62 == array_addr[13:5] ? valid_98 : _GEN_121; // @[DCache.scala 78:{33,33}]
  wire  _GEN_123 = 9'h63 == array_addr[13:5] ? valid_99 : _GEN_122; // @[DCache.scala 78:{33,33}]
  wire  _GEN_124 = 9'h64 == array_addr[13:5] ? valid_100 : _GEN_123; // @[DCache.scala 78:{33,33}]
  wire  _GEN_125 = 9'h65 == array_addr[13:5] ? valid_101 : _GEN_124; // @[DCache.scala 78:{33,33}]
  wire  _GEN_126 = 9'h66 == array_addr[13:5] ? valid_102 : _GEN_125; // @[DCache.scala 78:{33,33}]
  wire  _GEN_127 = 9'h67 == array_addr[13:5] ? valid_103 : _GEN_126; // @[DCache.scala 78:{33,33}]
  wire  _GEN_128 = 9'h68 == array_addr[13:5] ? valid_104 : _GEN_127; // @[DCache.scala 78:{33,33}]
  wire  _GEN_129 = 9'h69 == array_addr[13:5] ? valid_105 : _GEN_128; // @[DCache.scala 78:{33,33}]
  wire  _GEN_130 = 9'h6a == array_addr[13:5] ? valid_106 : _GEN_129; // @[DCache.scala 78:{33,33}]
  wire  _GEN_131 = 9'h6b == array_addr[13:5] ? valid_107 : _GEN_130; // @[DCache.scala 78:{33,33}]
  wire  _GEN_132 = 9'h6c == array_addr[13:5] ? valid_108 : _GEN_131; // @[DCache.scala 78:{33,33}]
  wire  _GEN_133 = 9'h6d == array_addr[13:5] ? valid_109 : _GEN_132; // @[DCache.scala 78:{33,33}]
  wire  _GEN_134 = 9'h6e == array_addr[13:5] ? valid_110 : _GEN_133; // @[DCache.scala 78:{33,33}]
  wire  _GEN_135 = 9'h6f == array_addr[13:5] ? valid_111 : _GEN_134; // @[DCache.scala 78:{33,33}]
  wire  _GEN_136 = 9'h70 == array_addr[13:5] ? valid_112 : _GEN_135; // @[DCache.scala 78:{33,33}]
  wire  _GEN_137 = 9'h71 == array_addr[13:5] ? valid_113 : _GEN_136; // @[DCache.scala 78:{33,33}]
  wire  _GEN_138 = 9'h72 == array_addr[13:5] ? valid_114 : _GEN_137; // @[DCache.scala 78:{33,33}]
  wire  _GEN_139 = 9'h73 == array_addr[13:5] ? valid_115 : _GEN_138; // @[DCache.scala 78:{33,33}]
  wire  _GEN_140 = 9'h74 == array_addr[13:5] ? valid_116 : _GEN_139; // @[DCache.scala 78:{33,33}]
  wire  _GEN_141 = 9'h75 == array_addr[13:5] ? valid_117 : _GEN_140; // @[DCache.scala 78:{33,33}]
  wire  _GEN_142 = 9'h76 == array_addr[13:5] ? valid_118 : _GEN_141; // @[DCache.scala 78:{33,33}]
  wire  _GEN_143 = 9'h77 == array_addr[13:5] ? valid_119 : _GEN_142; // @[DCache.scala 78:{33,33}]
  wire  _GEN_144 = 9'h78 == array_addr[13:5] ? valid_120 : _GEN_143; // @[DCache.scala 78:{33,33}]
  wire  _GEN_145 = 9'h79 == array_addr[13:5] ? valid_121 : _GEN_144; // @[DCache.scala 78:{33,33}]
  wire  _GEN_146 = 9'h7a == array_addr[13:5] ? valid_122 : _GEN_145; // @[DCache.scala 78:{33,33}]
  wire  _GEN_147 = 9'h7b == array_addr[13:5] ? valid_123 : _GEN_146; // @[DCache.scala 78:{33,33}]
  wire  _GEN_148 = 9'h7c == array_addr[13:5] ? valid_124 : _GEN_147; // @[DCache.scala 78:{33,33}]
  wire  _GEN_149 = 9'h7d == array_addr[13:5] ? valid_125 : _GEN_148; // @[DCache.scala 78:{33,33}]
  wire  _GEN_150 = 9'h7e == array_addr[13:5] ? valid_126 : _GEN_149; // @[DCache.scala 78:{33,33}]
  wire  _GEN_151 = 9'h7f == array_addr[13:5] ? valid_127 : _GEN_150; // @[DCache.scala 78:{33,33}]
  wire  _GEN_152 = 9'h80 == array_addr[13:5] ? valid_128 : _GEN_151; // @[DCache.scala 78:{33,33}]
  wire  _GEN_153 = 9'h81 == array_addr[13:5] ? valid_129 : _GEN_152; // @[DCache.scala 78:{33,33}]
  wire  _GEN_154 = 9'h82 == array_addr[13:5] ? valid_130 : _GEN_153; // @[DCache.scala 78:{33,33}]
  wire  _GEN_155 = 9'h83 == array_addr[13:5] ? valid_131 : _GEN_154; // @[DCache.scala 78:{33,33}]
  wire  _GEN_156 = 9'h84 == array_addr[13:5] ? valid_132 : _GEN_155; // @[DCache.scala 78:{33,33}]
  wire  _GEN_157 = 9'h85 == array_addr[13:5] ? valid_133 : _GEN_156; // @[DCache.scala 78:{33,33}]
  wire  _GEN_158 = 9'h86 == array_addr[13:5] ? valid_134 : _GEN_157; // @[DCache.scala 78:{33,33}]
  wire  _GEN_159 = 9'h87 == array_addr[13:5] ? valid_135 : _GEN_158; // @[DCache.scala 78:{33,33}]
  wire  _GEN_160 = 9'h88 == array_addr[13:5] ? valid_136 : _GEN_159; // @[DCache.scala 78:{33,33}]
  wire  _GEN_161 = 9'h89 == array_addr[13:5] ? valid_137 : _GEN_160; // @[DCache.scala 78:{33,33}]
  wire  _GEN_162 = 9'h8a == array_addr[13:5] ? valid_138 : _GEN_161; // @[DCache.scala 78:{33,33}]
  wire  _GEN_163 = 9'h8b == array_addr[13:5] ? valid_139 : _GEN_162; // @[DCache.scala 78:{33,33}]
  wire  _GEN_164 = 9'h8c == array_addr[13:5] ? valid_140 : _GEN_163; // @[DCache.scala 78:{33,33}]
  wire  _GEN_165 = 9'h8d == array_addr[13:5] ? valid_141 : _GEN_164; // @[DCache.scala 78:{33,33}]
  wire  _GEN_166 = 9'h8e == array_addr[13:5] ? valid_142 : _GEN_165; // @[DCache.scala 78:{33,33}]
  wire  _GEN_167 = 9'h8f == array_addr[13:5] ? valid_143 : _GEN_166; // @[DCache.scala 78:{33,33}]
  wire  _GEN_168 = 9'h90 == array_addr[13:5] ? valid_144 : _GEN_167; // @[DCache.scala 78:{33,33}]
  wire  _GEN_169 = 9'h91 == array_addr[13:5] ? valid_145 : _GEN_168; // @[DCache.scala 78:{33,33}]
  wire  _GEN_170 = 9'h92 == array_addr[13:5] ? valid_146 : _GEN_169; // @[DCache.scala 78:{33,33}]
  wire  _GEN_171 = 9'h93 == array_addr[13:5] ? valid_147 : _GEN_170; // @[DCache.scala 78:{33,33}]
  wire  _GEN_172 = 9'h94 == array_addr[13:5] ? valid_148 : _GEN_171; // @[DCache.scala 78:{33,33}]
  wire  _GEN_173 = 9'h95 == array_addr[13:5] ? valid_149 : _GEN_172; // @[DCache.scala 78:{33,33}]
  wire  _GEN_174 = 9'h96 == array_addr[13:5] ? valid_150 : _GEN_173; // @[DCache.scala 78:{33,33}]
  wire  _GEN_175 = 9'h97 == array_addr[13:5] ? valid_151 : _GEN_174; // @[DCache.scala 78:{33,33}]
  wire  _GEN_176 = 9'h98 == array_addr[13:5] ? valid_152 : _GEN_175; // @[DCache.scala 78:{33,33}]
  wire  _GEN_177 = 9'h99 == array_addr[13:5] ? valid_153 : _GEN_176; // @[DCache.scala 78:{33,33}]
  wire  _GEN_178 = 9'h9a == array_addr[13:5] ? valid_154 : _GEN_177; // @[DCache.scala 78:{33,33}]
  wire  _GEN_179 = 9'h9b == array_addr[13:5] ? valid_155 : _GEN_178; // @[DCache.scala 78:{33,33}]
  wire  _GEN_180 = 9'h9c == array_addr[13:5] ? valid_156 : _GEN_179; // @[DCache.scala 78:{33,33}]
  wire  _GEN_181 = 9'h9d == array_addr[13:5] ? valid_157 : _GEN_180; // @[DCache.scala 78:{33,33}]
  wire  _GEN_182 = 9'h9e == array_addr[13:5] ? valid_158 : _GEN_181; // @[DCache.scala 78:{33,33}]
  wire  _GEN_183 = 9'h9f == array_addr[13:5] ? valid_159 : _GEN_182; // @[DCache.scala 78:{33,33}]
  wire  _GEN_184 = 9'ha0 == array_addr[13:5] ? valid_160 : _GEN_183; // @[DCache.scala 78:{33,33}]
  wire  _GEN_185 = 9'ha1 == array_addr[13:5] ? valid_161 : _GEN_184; // @[DCache.scala 78:{33,33}]
  wire  _GEN_186 = 9'ha2 == array_addr[13:5] ? valid_162 : _GEN_185; // @[DCache.scala 78:{33,33}]
  wire  _GEN_187 = 9'ha3 == array_addr[13:5] ? valid_163 : _GEN_186; // @[DCache.scala 78:{33,33}]
  wire  _GEN_188 = 9'ha4 == array_addr[13:5] ? valid_164 : _GEN_187; // @[DCache.scala 78:{33,33}]
  wire  _GEN_189 = 9'ha5 == array_addr[13:5] ? valid_165 : _GEN_188; // @[DCache.scala 78:{33,33}]
  wire  _GEN_190 = 9'ha6 == array_addr[13:5] ? valid_166 : _GEN_189; // @[DCache.scala 78:{33,33}]
  wire  _GEN_191 = 9'ha7 == array_addr[13:5] ? valid_167 : _GEN_190; // @[DCache.scala 78:{33,33}]
  wire  _GEN_192 = 9'ha8 == array_addr[13:5] ? valid_168 : _GEN_191; // @[DCache.scala 78:{33,33}]
  wire  _GEN_193 = 9'ha9 == array_addr[13:5] ? valid_169 : _GEN_192; // @[DCache.scala 78:{33,33}]
  wire  _GEN_194 = 9'haa == array_addr[13:5] ? valid_170 : _GEN_193; // @[DCache.scala 78:{33,33}]
  wire  _GEN_195 = 9'hab == array_addr[13:5] ? valid_171 : _GEN_194; // @[DCache.scala 78:{33,33}]
  wire  _GEN_196 = 9'hac == array_addr[13:5] ? valid_172 : _GEN_195; // @[DCache.scala 78:{33,33}]
  wire  _GEN_197 = 9'had == array_addr[13:5] ? valid_173 : _GEN_196; // @[DCache.scala 78:{33,33}]
  wire  _GEN_198 = 9'hae == array_addr[13:5] ? valid_174 : _GEN_197; // @[DCache.scala 78:{33,33}]
  wire  _GEN_199 = 9'haf == array_addr[13:5] ? valid_175 : _GEN_198; // @[DCache.scala 78:{33,33}]
  wire  _GEN_200 = 9'hb0 == array_addr[13:5] ? valid_176 : _GEN_199; // @[DCache.scala 78:{33,33}]
  wire  _GEN_201 = 9'hb1 == array_addr[13:5] ? valid_177 : _GEN_200; // @[DCache.scala 78:{33,33}]
  wire  _GEN_202 = 9'hb2 == array_addr[13:5] ? valid_178 : _GEN_201; // @[DCache.scala 78:{33,33}]
  wire  _GEN_203 = 9'hb3 == array_addr[13:5] ? valid_179 : _GEN_202; // @[DCache.scala 78:{33,33}]
  wire  _GEN_204 = 9'hb4 == array_addr[13:5] ? valid_180 : _GEN_203; // @[DCache.scala 78:{33,33}]
  wire  _GEN_205 = 9'hb5 == array_addr[13:5] ? valid_181 : _GEN_204; // @[DCache.scala 78:{33,33}]
  wire  _GEN_206 = 9'hb6 == array_addr[13:5] ? valid_182 : _GEN_205; // @[DCache.scala 78:{33,33}]
  wire  _GEN_207 = 9'hb7 == array_addr[13:5] ? valid_183 : _GEN_206; // @[DCache.scala 78:{33,33}]
  wire  _GEN_208 = 9'hb8 == array_addr[13:5] ? valid_184 : _GEN_207; // @[DCache.scala 78:{33,33}]
  wire  _GEN_209 = 9'hb9 == array_addr[13:5] ? valid_185 : _GEN_208; // @[DCache.scala 78:{33,33}]
  wire  _GEN_210 = 9'hba == array_addr[13:5] ? valid_186 : _GEN_209; // @[DCache.scala 78:{33,33}]
  wire  _GEN_211 = 9'hbb == array_addr[13:5] ? valid_187 : _GEN_210; // @[DCache.scala 78:{33,33}]
  wire  _GEN_212 = 9'hbc == array_addr[13:5] ? valid_188 : _GEN_211; // @[DCache.scala 78:{33,33}]
  wire  _GEN_213 = 9'hbd == array_addr[13:5] ? valid_189 : _GEN_212; // @[DCache.scala 78:{33,33}]
  wire  _GEN_214 = 9'hbe == array_addr[13:5] ? valid_190 : _GEN_213; // @[DCache.scala 78:{33,33}]
  wire  _GEN_215 = 9'hbf == array_addr[13:5] ? valid_191 : _GEN_214; // @[DCache.scala 78:{33,33}]
  wire  _GEN_216 = 9'hc0 == array_addr[13:5] ? valid_192 : _GEN_215; // @[DCache.scala 78:{33,33}]
  wire  _GEN_217 = 9'hc1 == array_addr[13:5] ? valid_193 : _GEN_216; // @[DCache.scala 78:{33,33}]
  wire  _GEN_218 = 9'hc2 == array_addr[13:5] ? valid_194 : _GEN_217; // @[DCache.scala 78:{33,33}]
  wire  _GEN_219 = 9'hc3 == array_addr[13:5] ? valid_195 : _GEN_218; // @[DCache.scala 78:{33,33}]
  wire  _GEN_220 = 9'hc4 == array_addr[13:5] ? valid_196 : _GEN_219; // @[DCache.scala 78:{33,33}]
  wire  _GEN_221 = 9'hc5 == array_addr[13:5] ? valid_197 : _GEN_220; // @[DCache.scala 78:{33,33}]
  wire  _GEN_222 = 9'hc6 == array_addr[13:5] ? valid_198 : _GEN_221; // @[DCache.scala 78:{33,33}]
  wire  _GEN_223 = 9'hc7 == array_addr[13:5] ? valid_199 : _GEN_222; // @[DCache.scala 78:{33,33}]
  wire  _GEN_224 = 9'hc8 == array_addr[13:5] ? valid_200 : _GEN_223; // @[DCache.scala 78:{33,33}]
  wire  _GEN_225 = 9'hc9 == array_addr[13:5] ? valid_201 : _GEN_224; // @[DCache.scala 78:{33,33}]
  wire  _GEN_226 = 9'hca == array_addr[13:5] ? valid_202 : _GEN_225; // @[DCache.scala 78:{33,33}]
  wire  _GEN_227 = 9'hcb == array_addr[13:5] ? valid_203 : _GEN_226; // @[DCache.scala 78:{33,33}]
  wire  _GEN_228 = 9'hcc == array_addr[13:5] ? valid_204 : _GEN_227; // @[DCache.scala 78:{33,33}]
  wire  _GEN_229 = 9'hcd == array_addr[13:5] ? valid_205 : _GEN_228; // @[DCache.scala 78:{33,33}]
  wire  _GEN_230 = 9'hce == array_addr[13:5] ? valid_206 : _GEN_229; // @[DCache.scala 78:{33,33}]
  wire  _GEN_231 = 9'hcf == array_addr[13:5] ? valid_207 : _GEN_230; // @[DCache.scala 78:{33,33}]
  wire  _GEN_232 = 9'hd0 == array_addr[13:5] ? valid_208 : _GEN_231; // @[DCache.scala 78:{33,33}]
  wire  _GEN_233 = 9'hd1 == array_addr[13:5] ? valid_209 : _GEN_232; // @[DCache.scala 78:{33,33}]
  wire  _GEN_234 = 9'hd2 == array_addr[13:5] ? valid_210 : _GEN_233; // @[DCache.scala 78:{33,33}]
  wire  _GEN_235 = 9'hd3 == array_addr[13:5] ? valid_211 : _GEN_234; // @[DCache.scala 78:{33,33}]
  wire  _GEN_236 = 9'hd4 == array_addr[13:5] ? valid_212 : _GEN_235; // @[DCache.scala 78:{33,33}]
  wire  _GEN_237 = 9'hd5 == array_addr[13:5] ? valid_213 : _GEN_236; // @[DCache.scala 78:{33,33}]
  wire  _GEN_238 = 9'hd6 == array_addr[13:5] ? valid_214 : _GEN_237; // @[DCache.scala 78:{33,33}]
  wire  _GEN_239 = 9'hd7 == array_addr[13:5] ? valid_215 : _GEN_238; // @[DCache.scala 78:{33,33}]
  wire  _GEN_240 = 9'hd8 == array_addr[13:5] ? valid_216 : _GEN_239; // @[DCache.scala 78:{33,33}]
  wire  _GEN_241 = 9'hd9 == array_addr[13:5] ? valid_217 : _GEN_240; // @[DCache.scala 78:{33,33}]
  wire  _GEN_242 = 9'hda == array_addr[13:5] ? valid_218 : _GEN_241; // @[DCache.scala 78:{33,33}]
  wire  _GEN_243 = 9'hdb == array_addr[13:5] ? valid_219 : _GEN_242; // @[DCache.scala 78:{33,33}]
  wire  _GEN_244 = 9'hdc == array_addr[13:5] ? valid_220 : _GEN_243; // @[DCache.scala 78:{33,33}]
  wire  _GEN_245 = 9'hdd == array_addr[13:5] ? valid_221 : _GEN_244; // @[DCache.scala 78:{33,33}]
  wire  _GEN_246 = 9'hde == array_addr[13:5] ? valid_222 : _GEN_245; // @[DCache.scala 78:{33,33}]
  wire  _GEN_247 = 9'hdf == array_addr[13:5] ? valid_223 : _GEN_246; // @[DCache.scala 78:{33,33}]
  wire  _GEN_248 = 9'he0 == array_addr[13:5] ? valid_224 : _GEN_247; // @[DCache.scala 78:{33,33}]
  wire  _GEN_249 = 9'he1 == array_addr[13:5] ? valid_225 : _GEN_248; // @[DCache.scala 78:{33,33}]
  wire  _GEN_250 = 9'he2 == array_addr[13:5] ? valid_226 : _GEN_249; // @[DCache.scala 78:{33,33}]
  wire  _GEN_251 = 9'he3 == array_addr[13:5] ? valid_227 : _GEN_250; // @[DCache.scala 78:{33,33}]
  wire  _GEN_252 = 9'he4 == array_addr[13:5] ? valid_228 : _GEN_251; // @[DCache.scala 78:{33,33}]
  wire  _GEN_253 = 9'he5 == array_addr[13:5] ? valid_229 : _GEN_252; // @[DCache.scala 78:{33,33}]
  wire  _GEN_254 = 9'he6 == array_addr[13:5] ? valid_230 : _GEN_253; // @[DCache.scala 78:{33,33}]
  wire  _GEN_255 = 9'he7 == array_addr[13:5] ? valid_231 : _GEN_254; // @[DCache.scala 78:{33,33}]
  wire  _GEN_256 = 9'he8 == array_addr[13:5] ? valid_232 : _GEN_255; // @[DCache.scala 78:{33,33}]
  wire  _GEN_257 = 9'he9 == array_addr[13:5] ? valid_233 : _GEN_256; // @[DCache.scala 78:{33,33}]
  wire  _GEN_258 = 9'hea == array_addr[13:5] ? valid_234 : _GEN_257; // @[DCache.scala 78:{33,33}]
  wire  _GEN_259 = 9'heb == array_addr[13:5] ? valid_235 : _GEN_258; // @[DCache.scala 78:{33,33}]
  wire  _GEN_260 = 9'hec == array_addr[13:5] ? valid_236 : _GEN_259; // @[DCache.scala 78:{33,33}]
  wire  _GEN_261 = 9'hed == array_addr[13:5] ? valid_237 : _GEN_260; // @[DCache.scala 78:{33,33}]
  wire  _GEN_262 = 9'hee == array_addr[13:5] ? valid_238 : _GEN_261; // @[DCache.scala 78:{33,33}]
  wire  _GEN_263 = 9'hef == array_addr[13:5] ? valid_239 : _GEN_262; // @[DCache.scala 78:{33,33}]
  wire  _GEN_264 = 9'hf0 == array_addr[13:5] ? valid_240 : _GEN_263; // @[DCache.scala 78:{33,33}]
  wire  _GEN_265 = 9'hf1 == array_addr[13:5] ? valid_241 : _GEN_264; // @[DCache.scala 78:{33,33}]
  wire  _GEN_266 = 9'hf2 == array_addr[13:5] ? valid_242 : _GEN_265; // @[DCache.scala 78:{33,33}]
  wire  _GEN_267 = 9'hf3 == array_addr[13:5] ? valid_243 : _GEN_266; // @[DCache.scala 78:{33,33}]
  wire  _GEN_268 = 9'hf4 == array_addr[13:5] ? valid_244 : _GEN_267; // @[DCache.scala 78:{33,33}]
  wire  _GEN_269 = 9'hf5 == array_addr[13:5] ? valid_245 : _GEN_268; // @[DCache.scala 78:{33,33}]
  wire  _GEN_270 = 9'hf6 == array_addr[13:5] ? valid_246 : _GEN_269; // @[DCache.scala 78:{33,33}]
  wire  _GEN_271 = 9'hf7 == array_addr[13:5] ? valid_247 : _GEN_270; // @[DCache.scala 78:{33,33}]
  wire  _GEN_272 = 9'hf8 == array_addr[13:5] ? valid_248 : _GEN_271; // @[DCache.scala 78:{33,33}]
  wire  _GEN_273 = 9'hf9 == array_addr[13:5] ? valid_249 : _GEN_272; // @[DCache.scala 78:{33,33}]
  wire  _GEN_274 = 9'hfa == array_addr[13:5] ? valid_250 : _GEN_273; // @[DCache.scala 78:{33,33}]
  wire  _GEN_275 = 9'hfb == array_addr[13:5] ? valid_251 : _GEN_274; // @[DCache.scala 78:{33,33}]
  wire  _GEN_276 = 9'hfc == array_addr[13:5] ? valid_252 : _GEN_275; // @[DCache.scala 78:{33,33}]
  wire  _GEN_277 = 9'hfd == array_addr[13:5] ? valid_253 : _GEN_276; // @[DCache.scala 78:{33,33}]
  wire  _GEN_278 = 9'hfe == array_addr[13:5] ? valid_254 : _GEN_277; // @[DCache.scala 78:{33,33}]
  wire  _GEN_279 = 9'hff == array_addr[13:5] ? valid_255 : _GEN_278; // @[DCache.scala 78:{33,33}]
  wire  _GEN_280 = 9'h100 == array_addr[13:5] ? valid_256 : _GEN_279; // @[DCache.scala 78:{33,33}]
  wire  _GEN_281 = 9'h101 == array_addr[13:5] ? valid_257 : _GEN_280; // @[DCache.scala 78:{33,33}]
  wire  _GEN_282 = 9'h102 == array_addr[13:5] ? valid_258 : _GEN_281; // @[DCache.scala 78:{33,33}]
  wire  _GEN_283 = 9'h103 == array_addr[13:5] ? valid_259 : _GEN_282; // @[DCache.scala 78:{33,33}]
  wire  _GEN_284 = 9'h104 == array_addr[13:5] ? valid_260 : _GEN_283; // @[DCache.scala 78:{33,33}]
  wire  _GEN_285 = 9'h105 == array_addr[13:5] ? valid_261 : _GEN_284; // @[DCache.scala 78:{33,33}]
  wire  _GEN_286 = 9'h106 == array_addr[13:5] ? valid_262 : _GEN_285; // @[DCache.scala 78:{33,33}]
  wire  _GEN_287 = 9'h107 == array_addr[13:5] ? valid_263 : _GEN_286; // @[DCache.scala 78:{33,33}]
  wire  _GEN_288 = 9'h108 == array_addr[13:5] ? valid_264 : _GEN_287; // @[DCache.scala 78:{33,33}]
  wire  _GEN_289 = 9'h109 == array_addr[13:5] ? valid_265 : _GEN_288; // @[DCache.scala 78:{33,33}]
  wire  _GEN_290 = 9'h10a == array_addr[13:5] ? valid_266 : _GEN_289; // @[DCache.scala 78:{33,33}]
  wire  _GEN_291 = 9'h10b == array_addr[13:5] ? valid_267 : _GEN_290; // @[DCache.scala 78:{33,33}]
  wire  _GEN_292 = 9'h10c == array_addr[13:5] ? valid_268 : _GEN_291; // @[DCache.scala 78:{33,33}]
  wire  _GEN_293 = 9'h10d == array_addr[13:5] ? valid_269 : _GEN_292; // @[DCache.scala 78:{33,33}]
  wire  _GEN_294 = 9'h10e == array_addr[13:5] ? valid_270 : _GEN_293; // @[DCache.scala 78:{33,33}]
  wire  _GEN_295 = 9'h10f == array_addr[13:5] ? valid_271 : _GEN_294; // @[DCache.scala 78:{33,33}]
  wire  _GEN_296 = 9'h110 == array_addr[13:5] ? valid_272 : _GEN_295; // @[DCache.scala 78:{33,33}]
  wire  _GEN_297 = 9'h111 == array_addr[13:5] ? valid_273 : _GEN_296; // @[DCache.scala 78:{33,33}]
  wire  _GEN_298 = 9'h112 == array_addr[13:5] ? valid_274 : _GEN_297; // @[DCache.scala 78:{33,33}]
  wire  _GEN_299 = 9'h113 == array_addr[13:5] ? valid_275 : _GEN_298; // @[DCache.scala 78:{33,33}]
  wire  _GEN_300 = 9'h114 == array_addr[13:5] ? valid_276 : _GEN_299; // @[DCache.scala 78:{33,33}]
  wire  _GEN_301 = 9'h115 == array_addr[13:5] ? valid_277 : _GEN_300; // @[DCache.scala 78:{33,33}]
  wire  _GEN_302 = 9'h116 == array_addr[13:5] ? valid_278 : _GEN_301; // @[DCache.scala 78:{33,33}]
  wire  _GEN_303 = 9'h117 == array_addr[13:5] ? valid_279 : _GEN_302; // @[DCache.scala 78:{33,33}]
  wire  _GEN_304 = 9'h118 == array_addr[13:5] ? valid_280 : _GEN_303; // @[DCache.scala 78:{33,33}]
  wire  _GEN_305 = 9'h119 == array_addr[13:5] ? valid_281 : _GEN_304; // @[DCache.scala 78:{33,33}]
  wire  _GEN_306 = 9'h11a == array_addr[13:5] ? valid_282 : _GEN_305; // @[DCache.scala 78:{33,33}]
  wire  _GEN_307 = 9'h11b == array_addr[13:5] ? valid_283 : _GEN_306; // @[DCache.scala 78:{33,33}]
  wire  _GEN_308 = 9'h11c == array_addr[13:5] ? valid_284 : _GEN_307; // @[DCache.scala 78:{33,33}]
  wire  _GEN_309 = 9'h11d == array_addr[13:5] ? valid_285 : _GEN_308; // @[DCache.scala 78:{33,33}]
  wire  _GEN_310 = 9'h11e == array_addr[13:5] ? valid_286 : _GEN_309; // @[DCache.scala 78:{33,33}]
  wire  _GEN_311 = 9'h11f == array_addr[13:5] ? valid_287 : _GEN_310; // @[DCache.scala 78:{33,33}]
  wire  _GEN_312 = 9'h120 == array_addr[13:5] ? valid_288 : _GEN_311; // @[DCache.scala 78:{33,33}]
  wire  _GEN_313 = 9'h121 == array_addr[13:5] ? valid_289 : _GEN_312; // @[DCache.scala 78:{33,33}]
  wire  _GEN_314 = 9'h122 == array_addr[13:5] ? valid_290 : _GEN_313; // @[DCache.scala 78:{33,33}]
  wire  _GEN_315 = 9'h123 == array_addr[13:5] ? valid_291 : _GEN_314; // @[DCache.scala 78:{33,33}]
  wire  _GEN_316 = 9'h124 == array_addr[13:5] ? valid_292 : _GEN_315; // @[DCache.scala 78:{33,33}]
  wire  _GEN_317 = 9'h125 == array_addr[13:5] ? valid_293 : _GEN_316; // @[DCache.scala 78:{33,33}]
  wire  _GEN_318 = 9'h126 == array_addr[13:5] ? valid_294 : _GEN_317; // @[DCache.scala 78:{33,33}]
  wire  _GEN_319 = 9'h127 == array_addr[13:5] ? valid_295 : _GEN_318; // @[DCache.scala 78:{33,33}]
  wire  _GEN_320 = 9'h128 == array_addr[13:5] ? valid_296 : _GEN_319; // @[DCache.scala 78:{33,33}]
  wire  _GEN_321 = 9'h129 == array_addr[13:5] ? valid_297 : _GEN_320; // @[DCache.scala 78:{33,33}]
  wire  _GEN_322 = 9'h12a == array_addr[13:5] ? valid_298 : _GEN_321; // @[DCache.scala 78:{33,33}]
  wire  _GEN_323 = 9'h12b == array_addr[13:5] ? valid_299 : _GEN_322; // @[DCache.scala 78:{33,33}]
  wire  _GEN_324 = 9'h12c == array_addr[13:5] ? valid_300 : _GEN_323; // @[DCache.scala 78:{33,33}]
  wire  _GEN_325 = 9'h12d == array_addr[13:5] ? valid_301 : _GEN_324; // @[DCache.scala 78:{33,33}]
  wire  _GEN_326 = 9'h12e == array_addr[13:5] ? valid_302 : _GEN_325; // @[DCache.scala 78:{33,33}]
  wire  _GEN_327 = 9'h12f == array_addr[13:5] ? valid_303 : _GEN_326; // @[DCache.scala 78:{33,33}]
  wire  _GEN_328 = 9'h130 == array_addr[13:5] ? valid_304 : _GEN_327; // @[DCache.scala 78:{33,33}]
  wire  _GEN_329 = 9'h131 == array_addr[13:5] ? valid_305 : _GEN_328; // @[DCache.scala 78:{33,33}]
  wire  _GEN_330 = 9'h132 == array_addr[13:5] ? valid_306 : _GEN_329; // @[DCache.scala 78:{33,33}]
  wire  _GEN_331 = 9'h133 == array_addr[13:5] ? valid_307 : _GEN_330; // @[DCache.scala 78:{33,33}]
  wire  _GEN_332 = 9'h134 == array_addr[13:5] ? valid_308 : _GEN_331; // @[DCache.scala 78:{33,33}]
  wire  _GEN_333 = 9'h135 == array_addr[13:5] ? valid_309 : _GEN_332; // @[DCache.scala 78:{33,33}]
  wire  _GEN_334 = 9'h136 == array_addr[13:5] ? valid_310 : _GEN_333; // @[DCache.scala 78:{33,33}]
  wire  _GEN_335 = 9'h137 == array_addr[13:5] ? valid_311 : _GEN_334; // @[DCache.scala 78:{33,33}]
  wire  _GEN_336 = 9'h138 == array_addr[13:5] ? valid_312 : _GEN_335; // @[DCache.scala 78:{33,33}]
  wire  _GEN_337 = 9'h139 == array_addr[13:5] ? valid_313 : _GEN_336; // @[DCache.scala 78:{33,33}]
  wire  _GEN_338 = 9'h13a == array_addr[13:5] ? valid_314 : _GEN_337; // @[DCache.scala 78:{33,33}]
  wire  _GEN_339 = 9'h13b == array_addr[13:5] ? valid_315 : _GEN_338; // @[DCache.scala 78:{33,33}]
  wire  _GEN_340 = 9'h13c == array_addr[13:5] ? valid_316 : _GEN_339; // @[DCache.scala 78:{33,33}]
  wire  _GEN_341 = 9'h13d == array_addr[13:5] ? valid_317 : _GEN_340; // @[DCache.scala 78:{33,33}]
  wire  _GEN_342 = 9'h13e == array_addr[13:5] ? valid_318 : _GEN_341; // @[DCache.scala 78:{33,33}]
  wire  _GEN_343 = 9'h13f == array_addr[13:5] ? valid_319 : _GEN_342; // @[DCache.scala 78:{33,33}]
  wire  _GEN_344 = 9'h140 == array_addr[13:5] ? valid_320 : _GEN_343; // @[DCache.scala 78:{33,33}]
  wire  _GEN_345 = 9'h141 == array_addr[13:5] ? valid_321 : _GEN_344; // @[DCache.scala 78:{33,33}]
  wire  _GEN_346 = 9'h142 == array_addr[13:5] ? valid_322 : _GEN_345; // @[DCache.scala 78:{33,33}]
  wire  _GEN_347 = 9'h143 == array_addr[13:5] ? valid_323 : _GEN_346; // @[DCache.scala 78:{33,33}]
  wire  _GEN_348 = 9'h144 == array_addr[13:5] ? valid_324 : _GEN_347; // @[DCache.scala 78:{33,33}]
  wire  _GEN_349 = 9'h145 == array_addr[13:5] ? valid_325 : _GEN_348; // @[DCache.scala 78:{33,33}]
  wire  _GEN_350 = 9'h146 == array_addr[13:5] ? valid_326 : _GEN_349; // @[DCache.scala 78:{33,33}]
  wire  _GEN_351 = 9'h147 == array_addr[13:5] ? valid_327 : _GEN_350; // @[DCache.scala 78:{33,33}]
  wire  _GEN_352 = 9'h148 == array_addr[13:5] ? valid_328 : _GEN_351; // @[DCache.scala 78:{33,33}]
  wire  _GEN_353 = 9'h149 == array_addr[13:5] ? valid_329 : _GEN_352; // @[DCache.scala 78:{33,33}]
  wire  _GEN_354 = 9'h14a == array_addr[13:5] ? valid_330 : _GEN_353; // @[DCache.scala 78:{33,33}]
  wire  _GEN_355 = 9'h14b == array_addr[13:5] ? valid_331 : _GEN_354; // @[DCache.scala 78:{33,33}]
  wire  _GEN_356 = 9'h14c == array_addr[13:5] ? valid_332 : _GEN_355; // @[DCache.scala 78:{33,33}]
  wire  _GEN_357 = 9'h14d == array_addr[13:5] ? valid_333 : _GEN_356; // @[DCache.scala 78:{33,33}]
  wire  _GEN_358 = 9'h14e == array_addr[13:5] ? valid_334 : _GEN_357; // @[DCache.scala 78:{33,33}]
  wire  _GEN_359 = 9'h14f == array_addr[13:5] ? valid_335 : _GEN_358; // @[DCache.scala 78:{33,33}]
  wire  _GEN_360 = 9'h150 == array_addr[13:5] ? valid_336 : _GEN_359; // @[DCache.scala 78:{33,33}]
  wire  _GEN_361 = 9'h151 == array_addr[13:5] ? valid_337 : _GEN_360; // @[DCache.scala 78:{33,33}]
  wire  _GEN_362 = 9'h152 == array_addr[13:5] ? valid_338 : _GEN_361; // @[DCache.scala 78:{33,33}]
  wire  _GEN_363 = 9'h153 == array_addr[13:5] ? valid_339 : _GEN_362; // @[DCache.scala 78:{33,33}]
  wire  _GEN_364 = 9'h154 == array_addr[13:5] ? valid_340 : _GEN_363; // @[DCache.scala 78:{33,33}]
  wire  _GEN_365 = 9'h155 == array_addr[13:5] ? valid_341 : _GEN_364; // @[DCache.scala 78:{33,33}]
  wire  _GEN_366 = 9'h156 == array_addr[13:5] ? valid_342 : _GEN_365; // @[DCache.scala 78:{33,33}]
  wire  _GEN_367 = 9'h157 == array_addr[13:5] ? valid_343 : _GEN_366; // @[DCache.scala 78:{33,33}]
  wire  _GEN_368 = 9'h158 == array_addr[13:5] ? valid_344 : _GEN_367; // @[DCache.scala 78:{33,33}]
  wire  _GEN_369 = 9'h159 == array_addr[13:5] ? valid_345 : _GEN_368; // @[DCache.scala 78:{33,33}]
  wire  _GEN_370 = 9'h15a == array_addr[13:5] ? valid_346 : _GEN_369; // @[DCache.scala 78:{33,33}]
  wire  _GEN_371 = 9'h15b == array_addr[13:5] ? valid_347 : _GEN_370; // @[DCache.scala 78:{33,33}]
  wire  _GEN_372 = 9'h15c == array_addr[13:5] ? valid_348 : _GEN_371; // @[DCache.scala 78:{33,33}]
  wire  _GEN_373 = 9'h15d == array_addr[13:5] ? valid_349 : _GEN_372; // @[DCache.scala 78:{33,33}]
  wire  _GEN_374 = 9'h15e == array_addr[13:5] ? valid_350 : _GEN_373; // @[DCache.scala 78:{33,33}]
  wire  _GEN_375 = 9'h15f == array_addr[13:5] ? valid_351 : _GEN_374; // @[DCache.scala 78:{33,33}]
  wire  _GEN_376 = 9'h160 == array_addr[13:5] ? valid_352 : _GEN_375; // @[DCache.scala 78:{33,33}]
  wire  _GEN_377 = 9'h161 == array_addr[13:5] ? valid_353 : _GEN_376; // @[DCache.scala 78:{33,33}]
  wire  _GEN_378 = 9'h162 == array_addr[13:5] ? valid_354 : _GEN_377; // @[DCache.scala 78:{33,33}]
  wire  _GEN_379 = 9'h163 == array_addr[13:5] ? valid_355 : _GEN_378; // @[DCache.scala 78:{33,33}]
  wire  _GEN_380 = 9'h164 == array_addr[13:5] ? valid_356 : _GEN_379; // @[DCache.scala 78:{33,33}]
  wire  _GEN_381 = 9'h165 == array_addr[13:5] ? valid_357 : _GEN_380; // @[DCache.scala 78:{33,33}]
  wire  _GEN_382 = 9'h166 == array_addr[13:5] ? valid_358 : _GEN_381; // @[DCache.scala 78:{33,33}]
  wire  _GEN_383 = 9'h167 == array_addr[13:5] ? valid_359 : _GEN_382; // @[DCache.scala 78:{33,33}]
  wire  _GEN_384 = 9'h168 == array_addr[13:5] ? valid_360 : _GEN_383; // @[DCache.scala 78:{33,33}]
  wire  _GEN_385 = 9'h169 == array_addr[13:5] ? valid_361 : _GEN_384; // @[DCache.scala 78:{33,33}]
  wire  _GEN_386 = 9'h16a == array_addr[13:5] ? valid_362 : _GEN_385; // @[DCache.scala 78:{33,33}]
  wire  _GEN_387 = 9'h16b == array_addr[13:5] ? valid_363 : _GEN_386; // @[DCache.scala 78:{33,33}]
  wire  _GEN_388 = 9'h16c == array_addr[13:5] ? valid_364 : _GEN_387; // @[DCache.scala 78:{33,33}]
  wire  _GEN_389 = 9'h16d == array_addr[13:5] ? valid_365 : _GEN_388; // @[DCache.scala 78:{33,33}]
  wire  _GEN_390 = 9'h16e == array_addr[13:5] ? valid_366 : _GEN_389; // @[DCache.scala 78:{33,33}]
  wire  _GEN_391 = 9'h16f == array_addr[13:5] ? valid_367 : _GEN_390; // @[DCache.scala 78:{33,33}]
  wire  _GEN_392 = 9'h170 == array_addr[13:5] ? valid_368 : _GEN_391; // @[DCache.scala 78:{33,33}]
  wire  _GEN_393 = 9'h171 == array_addr[13:5] ? valid_369 : _GEN_392; // @[DCache.scala 78:{33,33}]
  wire  _GEN_394 = 9'h172 == array_addr[13:5] ? valid_370 : _GEN_393; // @[DCache.scala 78:{33,33}]
  wire  _GEN_395 = 9'h173 == array_addr[13:5] ? valid_371 : _GEN_394; // @[DCache.scala 78:{33,33}]
  wire  _GEN_396 = 9'h174 == array_addr[13:5] ? valid_372 : _GEN_395; // @[DCache.scala 78:{33,33}]
  wire  _GEN_397 = 9'h175 == array_addr[13:5] ? valid_373 : _GEN_396; // @[DCache.scala 78:{33,33}]
  wire  _GEN_398 = 9'h176 == array_addr[13:5] ? valid_374 : _GEN_397; // @[DCache.scala 78:{33,33}]
  wire  _GEN_399 = 9'h177 == array_addr[13:5] ? valid_375 : _GEN_398; // @[DCache.scala 78:{33,33}]
  wire  _GEN_400 = 9'h178 == array_addr[13:5] ? valid_376 : _GEN_399; // @[DCache.scala 78:{33,33}]
  wire  _GEN_401 = 9'h179 == array_addr[13:5] ? valid_377 : _GEN_400; // @[DCache.scala 78:{33,33}]
  wire  _GEN_402 = 9'h17a == array_addr[13:5] ? valid_378 : _GEN_401; // @[DCache.scala 78:{33,33}]
  wire  _GEN_403 = 9'h17b == array_addr[13:5] ? valid_379 : _GEN_402; // @[DCache.scala 78:{33,33}]
  wire  _GEN_404 = 9'h17c == array_addr[13:5] ? valid_380 : _GEN_403; // @[DCache.scala 78:{33,33}]
  wire  _GEN_405 = 9'h17d == array_addr[13:5] ? valid_381 : _GEN_404; // @[DCache.scala 78:{33,33}]
  wire  _GEN_406 = 9'h17e == array_addr[13:5] ? valid_382 : _GEN_405; // @[DCache.scala 78:{33,33}]
  wire  _GEN_407 = 9'h17f == array_addr[13:5] ? valid_383 : _GEN_406; // @[DCache.scala 78:{33,33}]
  wire  _GEN_408 = 9'h180 == array_addr[13:5] ? valid_384 : _GEN_407; // @[DCache.scala 78:{33,33}]
  wire  _GEN_409 = 9'h181 == array_addr[13:5] ? valid_385 : _GEN_408; // @[DCache.scala 78:{33,33}]
  wire  _GEN_410 = 9'h182 == array_addr[13:5] ? valid_386 : _GEN_409; // @[DCache.scala 78:{33,33}]
  wire  _GEN_411 = 9'h183 == array_addr[13:5] ? valid_387 : _GEN_410; // @[DCache.scala 78:{33,33}]
  wire  _GEN_412 = 9'h184 == array_addr[13:5] ? valid_388 : _GEN_411; // @[DCache.scala 78:{33,33}]
  wire  _GEN_413 = 9'h185 == array_addr[13:5] ? valid_389 : _GEN_412; // @[DCache.scala 78:{33,33}]
  wire  _GEN_414 = 9'h186 == array_addr[13:5] ? valid_390 : _GEN_413; // @[DCache.scala 78:{33,33}]
  wire  _GEN_415 = 9'h187 == array_addr[13:5] ? valid_391 : _GEN_414; // @[DCache.scala 78:{33,33}]
  wire  _GEN_416 = 9'h188 == array_addr[13:5] ? valid_392 : _GEN_415; // @[DCache.scala 78:{33,33}]
  wire  _GEN_417 = 9'h189 == array_addr[13:5] ? valid_393 : _GEN_416; // @[DCache.scala 78:{33,33}]
  wire  _GEN_418 = 9'h18a == array_addr[13:5] ? valid_394 : _GEN_417; // @[DCache.scala 78:{33,33}]
  wire  _GEN_419 = 9'h18b == array_addr[13:5] ? valid_395 : _GEN_418; // @[DCache.scala 78:{33,33}]
  wire  _GEN_420 = 9'h18c == array_addr[13:5] ? valid_396 : _GEN_419; // @[DCache.scala 78:{33,33}]
  wire  _GEN_421 = 9'h18d == array_addr[13:5] ? valid_397 : _GEN_420; // @[DCache.scala 78:{33,33}]
  wire  _GEN_422 = 9'h18e == array_addr[13:5] ? valid_398 : _GEN_421; // @[DCache.scala 78:{33,33}]
  wire  _GEN_423 = 9'h18f == array_addr[13:5] ? valid_399 : _GEN_422; // @[DCache.scala 78:{33,33}]
  wire  _GEN_424 = 9'h190 == array_addr[13:5] ? valid_400 : _GEN_423; // @[DCache.scala 78:{33,33}]
  wire  _GEN_425 = 9'h191 == array_addr[13:5] ? valid_401 : _GEN_424; // @[DCache.scala 78:{33,33}]
  wire  _GEN_426 = 9'h192 == array_addr[13:5] ? valid_402 : _GEN_425; // @[DCache.scala 78:{33,33}]
  wire  _GEN_427 = 9'h193 == array_addr[13:5] ? valid_403 : _GEN_426; // @[DCache.scala 78:{33,33}]
  wire  _GEN_428 = 9'h194 == array_addr[13:5] ? valid_404 : _GEN_427; // @[DCache.scala 78:{33,33}]
  wire  _GEN_429 = 9'h195 == array_addr[13:5] ? valid_405 : _GEN_428; // @[DCache.scala 78:{33,33}]
  wire  _GEN_430 = 9'h196 == array_addr[13:5] ? valid_406 : _GEN_429; // @[DCache.scala 78:{33,33}]
  wire  _GEN_431 = 9'h197 == array_addr[13:5] ? valid_407 : _GEN_430; // @[DCache.scala 78:{33,33}]
  wire  _GEN_432 = 9'h198 == array_addr[13:5] ? valid_408 : _GEN_431; // @[DCache.scala 78:{33,33}]
  wire  _GEN_433 = 9'h199 == array_addr[13:5] ? valid_409 : _GEN_432; // @[DCache.scala 78:{33,33}]
  wire  _GEN_434 = 9'h19a == array_addr[13:5] ? valid_410 : _GEN_433; // @[DCache.scala 78:{33,33}]
  wire  _GEN_435 = 9'h19b == array_addr[13:5] ? valid_411 : _GEN_434; // @[DCache.scala 78:{33,33}]
  wire  _GEN_436 = 9'h19c == array_addr[13:5] ? valid_412 : _GEN_435; // @[DCache.scala 78:{33,33}]
  wire  _GEN_437 = 9'h19d == array_addr[13:5] ? valid_413 : _GEN_436; // @[DCache.scala 78:{33,33}]
  wire  _GEN_438 = 9'h19e == array_addr[13:5] ? valid_414 : _GEN_437; // @[DCache.scala 78:{33,33}]
  wire  _GEN_439 = 9'h19f == array_addr[13:5] ? valid_415 : _GEN_438; // @[DCache.scala 78:{33,33}]
  wire  _GEN_440 = 9'h1a0 == array_addr[13:5] ? valid_416 : _GEN_439; // @[DCache.scala 78:{33,33}]
  wire  _GEN_441 = 9'h1a1 == array_addr[13:5] ? valid_417 : _GEN_440; // @[DCache.scala 78:{33,33}]
  wire  _GEN_442 = 9'h1a2 == array_addr[13:5] ? valid_418 : _GEN_441; // @[DCache.scala 78:{33,33}]
  wire  _GEN_443 = 9'h1a3 == array_addr[13:5] ? valid_419 : _GEN_442; // @[DCache.scala 78:{33,33}]
  wire  _GEN_444 = 9'h1a4 == array_addr[13:5] ? valid_420 : _GEN_443; // @[DCache.scala 78:{33,33}]
  wire  _GEN_445 = 9'h1a5 == array_addr[13:5] ? valid_421 : _GEN_444; // @[DCache.scala 78:{33,33}]
  wire  _GEN_446 = 9'h1a6 == array_addr[13:5] ? valid_422 : _GEN_445; // @[DCache.scala 78:{33,33}]
  wire  _GEN_447 = 9'h1a7 == array_addr[13:5] ? valid_423 : _GEN_446; // @[DCache.scala 78:{33,33}]
  wire  _GEN_448 = 9'h1a8 == array_addr[13:5] ? valid_424 : _GEN_447; // @[DCache.scala 78:{33,33}]
  wire  _GEN_449 = 9'h1a9 == array_addr[13:5] ? valid_425 : _GEN_448; // @[DCache.scala 78:{33,33}]
  wire  _GEN_450 = 9'h1aa == array_addr[13:5] ? valid_426 : _GEN_449; // @[DCache.scala 78:{33,33}]
  wire  _GEN_451 = 9'h1ab == array_addr[13:5] ? valid_427 : _GEN_450; // @[DCache.scala 78:{33,33}]
  wire  _GEN_452 = 9'h1ac == array_addr[13:5] ? valid_428 : _GEN_451; // @[DCache.scala 78:{33,33}]
  wire  _GEN_453 = 9'h1ad == array_addr[13:5] ? valid_429 : _GEN_452; // @[DCache.scala 78:{33,33}]
  wire  _GEN_454 = 9'h1ae == array_addr[13:5] ? valid_430 : _GEN_453; // @[DCache.scala 78:{33,33}]
  wire  _GEN_455 = 9'h1af == array_addr[13:5] ? valid_431 : _GEN_454; // @[DCache.scala 78:{33,33}]
  wire  _GEN_456 = 9'h1b0 == array_addr[13:5] ? valid_432 : _GEN_455; // @[DCache.scala 78:{33,33}]
  wire  _GEN_457 = 9'h1b1 == array_addr[13:5] ? valid_433 : _GEN_456; // @[DCache.scala 78:{33,33}]
  wire  _GEN_458 = 9'h1b2 == array_addr[13:5] ? valid_434 : _GEN_457; // @[DCache.scala 78:{33,33}]
  wire  _GEN_459 = 9'h1b3 == array_addr[13:5] ? valid_435 : _GEN_458; // @[DCache.scala 78:{33,33}]
  wire  _GEN_460 = 9'h1b4 == array_addr[13:5] ? valid_436 : _GEN_459; // @[DCache.scala 78:{33,33}]
  wire  _GEN_461 = 9'h1b5 == array_addr[13:5] ? valid_437 : _GEN_460; // @[DCache.scala 78:{33,33}]
  wire  _GEN_462 = 9'h1b6 == array_addr[13:5] ? valid_438 : _GEN_461; // @[DCache.scala 78:{33,33}]
  wire  _GEN_463 = 9'h1b7 == array_addr[13:5] ? valid_439 : _GEN_462; // @[DCache.scala 78:{33,33}]
  wire  _GEN_464 = 9'h1b8 == array_addr[13:5] ? valid_440 : _GEN_463; // @[DCache.scala 78:{33,33}]
  wire  _GEN_465 = 9'h1b9 == array_addr[13:5] ? valid_441 : _GEN_464; // @[DCache.scala 78:{33,33}]
  wire  _GEN_466 = 9'h1ba == array_addr[13:5] ? valid_442 : _GEN_465; // @[DCache.scala 78:{33,33}]
  wire  _GEN_467 = 9'h1bb == array_addr[13:5] ? valid_443 : _GEN_466; // @[DCache.scala 78:{33,33}]
  wire  _GEN_468 = 9'h1bc == array_addr[13:5] ? valid_444 : _GEN_467; // @[DCache.scala 78:{33,33}]
  wire  _GEN_469 = 9'h1bd == array_addr[13:5] ? valid_445 : _GEN_468; // @[DCache.scala 78:{33,33}]
  wire  _GEN_470 = 9'h1be == array_addr[13:5] ? valid_446 : _GEN_469; // @[DCache.scala 78:{33,33}]
  wire  _GEN_471 = 9'h1bf == array_addr[13:5] ? valid_447 : _GEN_470; // @[DCache.scala 78:{33,33}]
  wire  _GEN_472 = 9'h1c0 == array_addr[13:5] ? valid_448 : _GEN_471; // @[DCache.scala 78:{33,33}]
  wire  _GEN_473 = 9'h1c1 == array_addr[13:5] ? valid_449 : _GEN_472; // @[DCache.scala 78:{33,33}]
  wire  _GEN_474 = 9'h1c2 == array_addr[13:5] ? valid_450 : _GEN_473; // @[DCache.scala 78:{33,33}]
  wire  _GEN_475 = 9'h1c3 == array_addr[13:5] ? valid_451 : _GEN_474; // @[DCache.scala 78:{33,33}]
  wire  _GEN_476 = 9'h1c4 == array_addr[13:5] ? valid_452 : _GEN_475; // @[DCache.scala 78:{33,33}]
  wire  _GEN_477 = 9'h1c5 == array_addr[13:5] ? valid_453 : _GEN_476; // @[DCache.scala 78:{33,33}]
  wire  _GEN_478 = 9'h1c6 == array_addr[13:5] ? valid_454 : _GEN_477; // @[DCache.scala 78:{33,33}]
  wire  _GEN_479 = 9'h1c7 == array_addr[13:5] ? valid_455 : _GEN_478; // @[DCache.scala 78:{33,33}]
  wire  _GEN_480 = 9'h1c8 == array_addr[13:5] ? valid_456 : _GEN_479; // @[DCache.scala 78:{33,33}]
  wire  _GEN_481 = 9'h1c9 == array_addr[13:5] ? valid_457 : _GEN_480; // @[DCache.scala 78:{33,33}]
  wire  _GEN_482 = 9'h1ca == array_addr[13:5] ? valid_458 : _GEN_481; // @[DCache.scala 78:{33,33}]
  wire  _GEN_483 = 9'h1cb == array_addr[13:5] ? valid_459 : _GEN_482; // @[DCache.scala 78:{33,33}]
  wire  _GEN_484 = 9'h1cc == array_addr[13:5] ? valid_460 : _GEN_483; // @[DCache.scala 78:{33,33}]
  wire  _GEN_485 = 9'h1cd == array_addr[13:5] ? valid_461 : _GEN_484; // @[DCache.scala 78:{33,33}]
  wire  _GEN_486 = 9'h1ce == array_addr[13:5] ? valid_462 : _GEN_485; // @[DCache.scala 78:{33,33}]
  wire  _GEN_487 = 9'h1cf == array_addr[13:5] ? valid_463 : _GEN_486; // @[DCache.scala 78:{33,33}]
  wire  _GEN_488 = 9'h1d0 == array_addr[13:5] ? valid_464 : _GEN_487; // @[DCache.scala 78:{33,33}]
  wire  _GEN_489 = 9'h1d1 == array_addr[13:5] ? valid_465 : _GEN_488; // @[DCache.scala 78:{33,33}]
  wire  _GEN_490 = 9'h1d2 == array_addr[13:5] ? valid_466 : _GEN_489; // @[DCache.scala 78:{33,33}]
  wire  _GEN_491 = 9'h1d3 == array_addr[13:5] ? valid_467 : _GEN_490; // @[DCache.scala 78:{33,33}]
  wire  _GEN_492 = 9'h1d4 == array_addr[13:5] ? valid_468 : _GEN_491; // @[DCache.scala 78:{33,33}]
  wire  _GEN_493 = 9'h1d5 == array_addr[13:5] ? valid_469 : _GEN_492; // @[DCache.scala 78:{33,33}]
  wire  _GEN_494 = 9'h1d6 == array_addr[13:5] ? valid_470 : _GEN_493; // @[DCache.scala 78:{33,33}]
  wire  _GEN_495 = 9'h1d7 == array_addr[13:5] ? valid_471 : _GEN_494; // @[DCache.scala 78:{33,33}]
  wire  _GEN_496 = 9'h1d8 == array_addr[13:5] ? valid_472 : _GEN_495; // @[DCache.scala 78:{33,33}]
  wire  _GEN_497 = 9'h1d9 == array_addr[13:5] ? valid_473 : _GEN_496; // @[DCache.scala 78:{33,33}]
  wire  _GEN_498 = 9'h1da == array_addr[13:5] ? valid_474 : _GEN_497; // @[DCache.scala 78:{33,33}]
  wire  _GEN_499 = 9'h1db == array_addr[13:5] ? valid_475 : _GEN_498; // @[DCache.scala 78:{33,33}]
  wire  _GEN_500 = 9'h1dc == array_addr[13:5] ? valid_476 : _GEN_499; // @[DCache.scala 78:{33,33}]
  wire  _GEN_501 = 9'h1dd == array_addr[13:5] ? valid_477 : _GEN_500; // @[DCache.scala 78:{33,33}]
  wire  _GEN_502 = 9'h1de == array_addr[13:5] ? valid_478 : _GEN_501; // @[DCache.scala 78:{33,33}]
  wire  _GEN_503 = 9'h1df == array_addr[13:5] ? valid_479 : _GEN_502; // @[DCache.scala 78:{33,33}]
  wire  _GEN_504 = 9'h1e0 == array_addr[13:5] ? valid_480 : _GEN_503; // @[DCache.scala 78:{33,33}]
  wire  _GEN_505 = 9'h1e1 == array_addr[13:5] ? valid_481 : _GEN_504; // @[DCache.scala 78:{33,33}]
  wire  _GEN_506 = 9'h1e2 == array_addr[13:5] ? valid_482 : _GEN_505; // @[DCache.scala 78:{33,33}]
  wire  _GEN_507 = 9'h1e3 == array_addr[13:5] ? valid_483 : _GEN_506; // @[DCache.scala 78:{33,33}]
  wire  _GEN_508 = 9'h1e4 == array_addr[13:5] ? valid_484 : _GEN_507; // @[DCache.scala 78:{33,33}]
  wire  _GEN_509 = 9'h1e5 == array_addr[13:5] ? valid_485 : _GEN_508; // @[DCache.scala 78:{33,33}]
  wire  _GEN_510 = 9'h1e6 == array_addr[13:5] ? valid_486 : _GEN_509; // @[DCache.scala 78:{33,33}]
  wire  _GEN_511 = 9'h1e7 == array_addr[13:5] ? valid_487 : _GEN_510; // @[DCache.scala 78:{33,33}]
  wire  _GEN_512 = 9'h1e8 == array_addr[13:5] ? valid_488 : _GEN_511; // @[DCache.scala 78:{33,33}]
  wire  _GEN_513 = 9'h1e9 == array_addr[13:5] ? valid_489 : _GEN_512; // @[DCache.scala 78:{33,33}]
  wire  _GEN_514 = 9'h1ea == array_addr[13:5] ? valid_490 : _GEN_513; // @[DCache.scala 78:{33,33}]
  wire  _GEN_515 = 9'h1eb == array_addr[13:5] ? valid_491 : _GEN_514; // @[DCache.scala 78:{33,33}]
  wire  _GEN_516 = 9'h1ec == array_addr[13:5] ? valid_492 : _GEN_515; // @[DCache.scala 78:{33,33}]
  wire  _GEN_517 = 9'h1ed == array_addr[13:5] ? valid_493 : _GEN_516; // @[DCache.scala 78:{33,33}]
  wire  _GEN_518 = 9'h1ee == array_addr[13:5] ? valid_494 : _GEN_517; // @[DCache.scala 78:{33,33}]
  wire  _GEN_519 = 9'h1ef == array_addr[13:5] ? valid_495 : _GEN_518; // @[DCache.scala 78:{33,33}]
  wire  _GEN_520 = 9'h1f0 == array_addr[13:5] ? valid_496 : _GEN_519; // @[DCache.scala 78:{33,33}]
  wire  _GEN_521 = 9'h1f1 == array_addr[13:5] ? valid_497 : _GEN_520; // @[DCache.scala 78:{33,33}]
  wire  _GEN_522 = 9'h1f2 == array_addr[13:5] ? valid_498 : _GEN_521; // @[DCache.scala 78:{33,33}]
  wire  _GEN_523 = 9'h1f3 == array_addr[13:5] ? valid_499 : _GEN_522; // @[DCache.scala 78:{33,33}]
  wire  _GEN_524 = 9'h1f4 == array_addr[13:5] ? valid_500 : _GEN_523; // @[DCache.scala 78:{33,33}]
  wire  _GEN_525 = 9'h1f5 == array_addr[13:5] ? valid_501 : _GEN_524; // @[DCache.scala 78:{33,33}]
  wire  _GEN_526 = 9'h1f6 == array_addr[13:5] ? valid_502 : _GEN_525; // @[DCache.scala 78:{33,33}]
  wire  _GEN_527 = 9'h1f7 == array_addr[13:5] ? valid_503 : _GEN_526; // @[DCache.scala 78:{33,33}]
  wire  _GEN_528 = 9'h1f8 == array_addr[13:5] ? valid_504 : _GEN_527; // @[DCache.scala 78:{33,33}]
  wire  _GEN_529 = 9'h1f9 == array_addr[13:5] ? valid_505 : _GEN_528; // @[DCache.scala 78:{33,33}]
  wire  _GEN_530 = 9'h1fa == array_addr[13:5] ? valid_506 : _GEN_529; // @[DCache.scala 78:{33,33}]
  wire  _GEN_531 = 9'h1fb == array_addr[13:5] ? valid_507 : _GEN_530; // @[DCache.scala 78:{33,33}]
  wire  _GEN_532 = 9'h1fc == array_addr[13:5] ? valid_508 : _GEN_531; // @[DCache.scala 78:{33,33}]
  wire  _GEN_533 = 9'h1fd == array_addr[13:5] ? valid_509 : _GEN_532; // @[DCache.scala 78:{33,33}]
  wire  _GEN_534 = 9'h1fe == array_addr[13:5] ? valid_510 : _GEN_533; // @[DCache.scala 78:{33,33}]
  wire  _GEN_535 = 9'h1ff == array_addr[13:5] ? valid_511 : _GEN_534; // @[DCache.scala 78:{33,33}]
  wire  array_hit = _GEN_535 & array_wdata_tag == array_out_tag; // @[DCache.scala 78:33]
  reg [26:0] lrsc_addr; // @[DCache.scala 128:30]
  wire  is_lr_r = req_r_lrsc & ~req_r_wen; // @[DCache.scala 131:34]
  wire  _GEN_536 = _array_io_en_T_1 & is_lr_r | lrsc_reserved; // @[DCache.scala 132:30 133:19 127:30]
  wire [4:0] _lrsc_counter_T_1 = lrsc_counter + 5'h1; // @[DCache.scala 137:34]
  wire  is_sc = io_cache_req_bits_lrsc & io_cache_req_bits_wen; // @[DCache.scala 143:33]
  wire  sc_fail = is_sc & (_x1_b_ready_T_1 | io_cache_req_bits_addr[31:5] != lrsc_addr); // @[DCache.scala 144:25]
  wire  is_sc_r = req_r_lrsc & req_r_wen; // @[DCache.scala 145:30]
  reg  sc_fail_r; // @[Reg.scala 35:20]
  wire [5:0] _sc_rdata_64_T_1 = {req_r_addr[2], 5'h0}; // @[DCache.scala 153:42]
  wire [63:0] _sc_rdata_64_T_2 = 64'h1 << _sc_rdata_64_T_1; // @[DCache.scala 153:24]
  wire [63:0] sc_rdata_64 = sc_fail_r ? _sc_rdata_64_T_2 : 64'h0; // @[DCache.scala 152:19 153:17 151:32]
  wire  _T_12 = ~sc_fail_r; // @[DCache.scala 171:12]
  wire  _GEN_545 = 9'h0 == array_addr[13:5] | valid_0; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_546 = 9'h1 == array_addr[13:5] | valid_1; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_547 = 9'h2 == array_addr[13:5] | valid_2; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_548 = 9'h3 == array_addr[13:5] | valid_3; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_549 = 9'h4 == array_addr[13:5] | valid_4; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_550 = 9'h5 == array_addr[13:5] | valid_5; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_551 = 9'h6 == array_addr[13:5] | valid_6; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_552 = 9'h7 == array_addr[13:5] | valid_7; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_553 = 9'h8 == array_addr[13:5] | valid_8; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_554 = 9'h9 == array_addr[13:5] | valid_9; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_555 = 9'ha == array_addr[13:5] | valid_10; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_556 = 9'hb == array_addr[13:5] | valid_11; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_557 = 9'hc == array_addr[13:5] | valid_12; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_558 = 9'hd == array_addr[13:5] | valid_13; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_559 = 9'he == array_addr[13:5] | valid_14; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_560 = 9'hf == array_addr[13:5] | valid_15; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_561 = 9'h10 == array_addr[13:5] | valid_16; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_562 = 9'h11 == array_addr[13:5] | valid_17; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_563 = 9'h12 == array_addr[13:5] | valid_18; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_564 = 9'h13 == array_addr[13:5] | valid_19; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_565 = 9'h14 == array_addr[13:5] | valid_20; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_566 = 9'h15 == array_addr[13:5] | valid_21; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_567 = 9'h16 == array_addr[13:5] | valid_22; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_568 = 9'h17 == array_addr[13:5] | valid_23; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_569 = 9'h18 == array_addr[13:5] | valid_24; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_570 = 9'h19 == array_addr[13:5] | valid_25; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_571 = 9'h1a == array_addr[13:5] | valid_26; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_572 = 9'h1b == array_addr[13:5] | valid_27; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_573 = 9'h1c == array_addr[13:5] | valid_28; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_574 = 9'h1d == array_addr[13:5] | valid_29; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_575 = 9'h1e == array_addr[13:5] | valid_30; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_576 = 9'h1f == array_addr[13:5] | valid_31; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_577 = 9'h20 == array_addr[13:5] | valid_32; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_578 = 9'h21 == array_addr[13:5] | valid_33; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_579 = 9'h22 == array_addr[13:5] | valid_34; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_580 = 9'h23 == array_addr[13:5] | valid_35; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_581 = 9'h24 == array_addr[13:5] | valid_36; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_582 = 9'h25 == array_addr[13:5] | valid_37; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_583 = 9'h26 == array_addr[13:5] | valid_38; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_584 = 9'h27 == array_addr[13:5] | valid_39; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_585 = 9'h28 == array_addr[13:5] | valid_40; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_586 = 9'h29 == array_addr[13:5] | valid_41; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_587 = 9'h2a == array_addr[13:5] | valid_42; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_588 = 9'h2b == array_addr[13:5] | valid_43; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_589 = 9'h2c == array_addr[13:5] | valid_44; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_590 = 9'h2d == array_addr[13:5] | valid_45; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_591 = 9'h2e == array_addr[13:5] | valid_46; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_592 = 9'h2f == array_addr[13:5] | valid_47; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_593 = 9'h30 == array_addr[13:5] | valid_48; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_594 = 9'h31 == array_addr[13:5] | valid_49; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_595 = 9'h32 == array_addr[13:5] | valid_50; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_596 = 9'h33 == array_addr[13:5] | valid_51; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_597 = 9'h34 == array_addr[13:5] | valid_52; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_598 = 9'h35 == array_addr[13:5] | valid_53; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_599 = 9'h36 == array_addr[13:5] | valid_54; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_600 = 9'h37 == array_addr[13:5] | valid_55; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_601 = 9'h38 == array_addr[13:5] | valid_56; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_602 = 9'h39 == array_addr[13:5] | valid_57; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_603 = 9'h3a == array_addr[13:5] | valid_58; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_604 = 9'h3b == array_addr[13:5] | valid_59; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_605 = 9'h3c == array_addr[13:5] | valid_60; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_606 = 9'h3d == array_addr[13:5] | valid_61; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_607 = 9'h3e == array_addr[13:5] | valid_62; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_608 = 9'h3f == array_addr[13:5] | valid_63; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_609 = 9'h40 == array_addr[13:5] | valid_64; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_610 = 9'h41 == array_addr[13:5] | valid_65; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_611 = 9'h42 == array_addr[13:5] | valid_66; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_612 = 9'h43 == array_addr[13:5] | valid_67; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_613 = 9'h44 == array_addr[13:5] | valid_68; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_614 = 9'h45 == array_addr[13:5] | valid_69; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_615 = 9'h46 == array_addr[13:5] | valid_70; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_616 = 9'h47 == array_addr[13:5] | valid_71; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_617 = 9'h48 == array_addr[13:5] | valid_72; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_618 = 9'h49 == array_addr[13:5] | valid_73; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_619 = 9'h4a == array_addr[13:5] | valid_74; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_620 = 9'h4b == array_addr[13:5] | valid_75; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_621 = 9'h4c == array_addr[13:5] | valid_76; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_622 = 9'h4d == array_addr[13:5] | valid_77; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_623 = 9'h4e == array_addr[13:5] | valid_78; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_624 = 9'h4f == array_addr[13:5] | valid_79; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_625 = 9'h50 == array_addr[13:5] | valid_80; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_626 = 9'h51 == array_addr[13:5] | valid_81; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_627 = 9'h52 == array_addr[13:5] | valid_82; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_628 = 9'h53 == array_addr[13:5] | valid_83; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_629 = 9'h54 == array_addr[13:5] | valid_84; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_630 = 9'h55 == array_addr[13:5] | valid_85; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_631 = 9'h56 == array_addr[13:5] | valid_86; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_632 = 9'h57 == array_addr[13:5] | valid_87; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_633 = 9'h58 == array_addr[13:5] | valid_88; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_634 = 9'h59 == array_addr[13:5] | valid_89; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_635 = 9'h5a == array_addr[13:5] | valid_90; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_636 = 9'h5b == array_addr[13:5] | valid_91; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_637 = 9'h5c == array_addr[13:5] | valid_92; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_638 = 9'h5d == array_addr[13:5] | valid_93; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_639 = 9'h5e == array_addr[13:5] | valid_94; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_640 = 9'h5f == array_addr[13:5] | valid_95; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_641 = 9'h60 == array_addr[13:5] | valid_96; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_642 = 9'h61 == array_addr[13:5] | valid_97; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_643 = 9'h62 == array_addr[13:5] | valid_98; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_644 = 9'h63 == array_addr[13:5] | valid_99; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_645 = 9'h64 == array_addr[13:5] | valid_100; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_646 = 9'h65 == array_addr[13:5] | valid_101; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_647 = 9'h66 == array_addr[13:5] | valid_102; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_648 = 9'h67 == array_addr[13:5] | valid_103; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_649 = 9'h68 == array_addr[13:5] | valid_104; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_650 = 9'h69 == array_addr[13:5] | valid_105; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_651 = 9'h6a == array_addr[13:5] | valid_106; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_652 = 9'h6b == array_addr[13:5] | valid_107; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_653 = 9'h6c == array_addr[13:5] | valid_108; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_654 = 9'h6d == array_addr[13:5] | valid_109; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_655 = 9'h6e == array_addr[13:5] | valid_110; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_656 = 9'h6f == array_addr[13:5] | valid_111; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_657 = 9'h70 == array_addr[13:5] | valid_112; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_658 = 9'h71 == array_addr[13:5] | valid_113; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_659 = 9'h72 == array_addr[13:5] | valid_114; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_660 = 9'h73 == array_addr[13:5] | valid_115; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_661 = 9'h74 == array_addr[13:5] | valid_116; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_662 = 9'h75 == array_addr[13:5] | valid_117; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_663 = 9'h76 == array_addr[13:5] | valid_118; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_664 = 9'h77 == array_addr[13:5] | valid_119; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_665 = 9'h78 == array_addr[13:5] | valid_120; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_666 = 9'h79 == array_addr[13:5] | valid_121; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_667 = 9'h7a == array_addr[13:5] | valid_122; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_668 = 9'h7b == array_addr[13:5] | valid_123; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_669 = 9'h7c == array_addr[13:5] | valid_124; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_670 = 9'h7d == array_addr[13:5] | valid_125; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_671 = 9'h7e == array_addr[13:5] | valid_126; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_672 = 9'h7f == array_addr[13:5] | valid_127; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_673 = 9'h80 == array_addr[13:5] | valid_128; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_674 = 9'h81 == array_addr[13:5] | valid_129; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_675 = 9'h82 == array_addr[13:5] | valid_130; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_676 = 9'h83 == array_addr[13:5] | valid_131; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_677 = 9'h84 == array_addr[13:5] | valid_132; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_678 = 9'h85 == array_addr[13:5] | valid_133; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_679 = 9'h86 == array_addr[13:5] | valid_134; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_680 = 9'h87 == array_addr[13:5] | valid_135; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_681 = 9'h88 == array_addr[13:5] | valid_136; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_682 = 9'h89 == array_addr[13:5] | valid_137; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_683 = 9'h8a == array_addr[13:5] | valid_138; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_684 = 9'h8b == array_addr[13:5] | valid_139; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_685 = 9'h8c == array_addr[13:5] | valid_140; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_686 = 9'h8d == array_addr[13:5] | valid_141; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_687 = 9'h8e == array_addr[13:5] | valid_142; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_688 = 9'h8f == array_addr[13:5] | valid_143; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_689 = 9'h90 == array_addr[13:5] | valid_144; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_690 = 9'h91 == array_addr[13:5] | valid_145; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_691 = 9'h92 == array_addr[13:5] | valid_146; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_692 = 9'h93 == array_addr[13:5] | valid_147; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_693 = 9'h94 == array_addr[13:5] | valid_148; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_694 = 9'h95 == array_addr[13:5] | valid_149; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_695 = 9'h96 == array_addr[13:5] | valid_150; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_696 = 9'h97 == array_addr[13:5] | valid_151; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_697 = 9'h98 == array_addr[13:5] | valid_152; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_698 = 9'h99 == array_addr[13:5] | valid_153; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_699 = 9'h9a == array_addr[13:5] | valid_154; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_700 = 9'h9b == array_addr[13:5] | valid_155; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_701 = 9'h9c == array_addr[13:5] | valid_156; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_702 = 9'h9d == array_addr[13:5] | valid_157; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_703 = 9'h9e == array_addr[13:5] | valid_158; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_704 = 9'h9f == array_addr[13:5] | valid_159; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_705 = 9'ha0 == array_addr[13:5] | valid_160; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_706 = 9'ha1 == array_addr[13:5] | valid_161; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_707 = 9'ha2 == array_addr[13:5] | valid_162; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_708 = 9'ha3 == array_addr[13:5] | valid_163; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_709 = 9'ha4 == array_addr[13:5] | valid_164; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_710 = 9'ha5 == array_addr[13:5] | valid_165; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_711 = 9'ha6 == array_addr[13:5] | valid_166; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_712 = 9'ha7 == array_addr[13:5] | valid_167; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_713 = 9'ha8 == array_addr[13:5] | valid_168; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_714 = 9'ha9 == array_addr[13:5] | valid_169; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_715 = 9'haa == array_addr[13:5] | valid_170; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_716 = 9'hab == array_addr[13:5] | valid_171; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_717 = 9'hac == array_addr[13:5] | valid_172; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_718 = 9'had == array_addr[13:5] | valid_173; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_719 = 9'hae == array_addr[13:5] | valid_174; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_720 = 9'haf == array_addr[13:5] | valid_175; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_721 = 9'hb0 == array_addr[13:5] | valid_176; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_722 = 9'hb1 == array_addr[13:5] | valid_177; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_723 = 9'hb2 == array_addr[13:5] | valid_178; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_724 = 9'hb3 == array_addr[13:5] | valid_179; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_725 = 9'hb4 == array_addr[13:5] | valid_180; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_726 = 9'hb5 == array_addr[13:5] | valid_181; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_727 = 9'hb6 == array_addr[13:5] | valid_182; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_728 = 9'hb7 == array_addr[13:5] | valid_183; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_729 = 9'hb8 == array_addr[13:5] | valid_184; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_730 = 9'hb9 == array_addr[13:5] | valid_185; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_731 = 9'hba == array_addr[13:5] | valid_186; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_732 = 9'hbb == array_addr[13:5] | valid_187; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_733 = 9'hbc == array_addr[13:5] | valid_188; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_734 = 9'hbd == array_addr[13:5] | valid_189; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_735 = 9'hbe == array_addr[13:5] | valid_190; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_736 = 9'hbf == array_addr[13:5] | valid_191; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_737 = 9'hc0 == array_addr[13:5] | valid_192; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_738 = 9'hc1 == array_addr[13:5] | valid_193; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_739 = 9'hc2 == array_addr[13:5] | valid_194; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_740 = 9'hc3 == array_addr[13:5] | valid_195; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_741 = 9'hc4 == array_addr[13:5] | valid_196; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_742 = 9'hc5 == array_addr[13:5] | valid_197; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_743 = 9'hc6 == array_addr[13:5] | valid_198; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_744 = 9'hc7 == array_addr[13:5] | valid_199; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_745 = 9'hc8 == array_addr[13:5] | valid_200; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_746 = 9'hc9 == array_addr[13:5] | valid_201; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_747 = 9'hca == array_addr[13:5] | valid_202; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_748 = 9'hcb == array_addr[13:5] | valid_203; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_749 = 9'hcc == array_addr[13:5] | valid_204; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_750 = 9'hcd == array_addr[13:5] | valid_205; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_751 = 9'hce == array_addr[13:5] | valid_206; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_752 = 9'hcf == array_addr[13:5] | valid_207; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_753 = 9'hd0 == array_addr[13:5] | valid_208; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_754 = 9'hd1 == array_addr[13:5] | valid_209; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_755 = 9'hd2 == array_addr[13:5] | valid_210; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_756 = 9'hd3 == array_addr[13:5] | valid_211; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_757 = 9'hd4 == array_addr[13:5] | valid_212; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_758 = 9'hd5 == array_addr[13:5] | valid_213; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_759 = 9'hd6 == array_addr[13:5] | valid_214; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_760 = 9'hd7 == array_addr[13:5] | valid_215; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_761 = 9'hd8 == array_addr[13:5] | valid_216; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_762 = 9'hd9 == array_addr[13:5] | valid_217; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_763 = 9'hda == array_addr[13:5] | valid_218; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_764 = 9'hdb == array_addr[13:5] | valid_219; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_765 = 9'hdc == array_addr[13:5] | valid_220; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_766 = 9'hdd == array_addr[13:5] | valid_221; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_767 = 9'hde == array_addr[13:5] | valid_222; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_768 = 9'hdf == array_addr[13:5] | valid_223; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_769 = 9'he0 == array_addr[13:5] | valid_224; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_770 = 9'he1 == array_addr[13:5] | valid_225; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_771 = 9'he2 == array_addr[13:5] | valid_226; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_772 = 9'he3 == array_addr[13:5] | valid_227; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_773 = 9'he4 == array_addr[13:5] | valid_228; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_774 = 9'he5 == array_addr[13:5] | valid_229; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_775 = 9'he6 == array_addr[13:5] | valid_230; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_776 = 9'he7 == array_addr[13:5] | valid_231; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_777 = 9'he8 == array_addr[13:5] | valid_232; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_778 = 9'he9 == array_addr[13:5] | valid_233; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_779 = 9'hea == array_addr[13:5] | valid_234; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_780 = 9'heb == array_addr[13:5] | valid_235; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_781 = 9'hec == array_addr[13:5] | valid_236; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_782 = 9'hed == array_addr[13:5] | valid_237; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_783 = 9'hee == array_addr[13:5] | valid_238; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_784 = 9'hef == array_addr[13:5] | valid_239; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_785 = 9'hf0 == array_addr[13:5] | valid_240; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_786 = 9'hf1 == array_addr[13:5] | valid_241; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_787 = 9'hf2 == array_addr[13:5] | valid_242; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_788 = 9'hf3 == array_addr[13:5] | valid_243; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_789 = 9'hf4 == array_addr[13:5] | valid_244; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_790 = 9'hf5 == array_addr[13:5] | valid_245; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_791 = 9'hf6 == array_addr[13:5] | valid_246; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_792 = 9'hf7 == array_addr[13:5] | valid_247; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_793 = 9'hf8 == array_addr[13:5] | valid_248; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_794 = 9'hf9 == array_addr[13:5] | valid_249; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_795 = 9'hfa == array_addr[13:5] | valid_250; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_796 = 9'hfb == array_addr[13:5] | valid_251; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_797 = 9'hfc == array_addr[13:5] | valid_252; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_798 = 9'hfd == array_addr[13:5] | valid_253; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_799 = 9'hfe == array_addr[13:5] | valid_254; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_800 = 9'hff == array_addr[13:5] | valid_255; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_801 = 9'h100 == array_addr[13:5] | valid_256; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_802 = 9'h101 == array_addr[13:5] | valid_257; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_803 = 9'h102 == array_addr[13:5] | valid_258; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_804 = 9'h103 == array_addr[13:5] | valid_259; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_805 = 9'h104 == array_addr[13:5] | valid_260; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_806 = 9'h105 == array_addr[13:5] | valid_261; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_807 = 9'h106 == array_addr[13:5] | valid_262; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_808 = 9'h107 == array_addr[13:5] | valid_263; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_809 = 9'h108 == array_addr[13:5] | valid_264; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_810 = 9'h109 == array_addr[13:5] | valid_265; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_811 = 9'h10a == array_addr[13:5] | valid_266; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_812 = 9'h10b == array_addr[13:5] | valid_267; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_813 = 9'h10c == array_addr[13:5] | valid_268; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_814 = 9'h10d == array_addr[13:5] | valid_269; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_815 = 9'h10e == array_addr[13:5] | valid_270; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_816 = 9'h10f == array_addr[13:5] | valid_271; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_817 = 9'h110 == array_addr[13:5] | valid_272; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_818 = 9'h111 == array_addr[13:5] | valid_273; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_819 = 9'h112 == array_addr[13:5] | valid_274; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_820 = 9'h113 == array_addr[13:5] | valid_275; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_821 = 9'h114 == array_addr[13:5] | valid_276; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_822 = 9'h115 == array_addr[13:5] | valid_277; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_823 = 9'h116 == array_addr[13:5] | valid_278; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_824 = 9'h117 == array_addr[13:5] | valid_279; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_825 = 9'h118 == array_addr[13:5] | valid_280; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_826 = 9'h119 == array_addr[13:5] | valid_281; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_827 = 9'h11a == array_addr[13:5] | valid_282; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_828 = 9'h11b == array_addr[13:5] | valid_283; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_829 = 9'h11c == array_addr[13:5] | valid_284; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_830 = 9'h11d == array_addr[13:5] | valid_285; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_831 = 9'h11e == array_addr[13:5] | valid_286; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_832 = 9'h11f == array_addr[13:5] | valid_287; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_833 = 9'h120 == array_addr[13:5] | valid_288; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_834 = 9'h121 == array_addr[13:5] | valid_289; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_835 = 9'h122 == array_addr[13:5] | valid_290; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_836 = 9'h123 == array_addr[13:5] | valid_291; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_837 = 9'h124 == array_addr[13:5] | valid_292; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_838 = 9'h125 == array_addr[13:5] | valid_293; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_839 = 9'h126 == array_addr[13:5] | valid_294; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_840 = 9'h127 == array_addr[13:5] | valid_295; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_841 = 9'h128 == array_addr[13:5] | valid_296; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_842 = 9'h129 == array_addr[13:5] | valid_297; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_843 = 9'h12a == array_addr[13:5] | valid_298; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_844 = 9'h12b == array_addr[13:5] | valid_299; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_845 = 9'h12c == array_addr[13:5] | valid_300; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_846 = 9'h12d == array_addr[13:5] | valid_301; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_847 = 9'h12e == array_addr[13:5] | valid_302; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_848 = 9'h12f == array_addr[13:5] | valid_303; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_849 = 9'h130 == array_addr[13:5] | valid_304; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_850 = 9'h131 == array_addr[13:5] | valid_305; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_851 = 9'h132 == array_addr[13:5] | valid_306; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_852 = 9'h133 == array_addr[13:5] | valid_307; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_853 = 9'h134 == array_addr[13:5] | valid_308; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_854 = 9'h135 == array_addr[13:5] | valid_309; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_855 = 9'h136 == array_addr[13:5] | valid_310; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_856 = 9'h137 == array_addr[13:5] | valid_311; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_857 = 9'h138 == array_addr[13:5] | valid_312; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_858 = 9'h139 == array_addr[13:5] | valid_313; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_859 = 9'h13a == array_addr[13:5] | valid_314; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_860 = 9'h13b == array_addr[13:5] | valid_315; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_861 = 9'h13c == array_addr[13:5] | valid_316; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_862 = 9'h13d == array_addr[13:5] | valid_317; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_863 = 9'h13e == array_addr[13:5] | valid_318; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_864 = 9'h13f == array_addr[13:5] | valid_319; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_865 = 9'h140 == array_addr[13:5] | valid_320; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_866 = 9'h141 == array_addr[13:5] | valid_321; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_867 = 9'h142 == array_addr[13:5] | valid_322; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_868 = 9'h143 == array_addr[13:5] | valid_323; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_869 = 9'h144 == array_addr[13:5] | valid_324; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_870 = 9'h145 == array_addr[13:5] | valid_325; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_871 = 9'h146 == array_addr[13:5] | valid_326; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_872 = 9'h147 == array_addr[13:5] | valid_327; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_873 = 9'h148 == array_addr[13:5] | valid_328; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_874 = 9'h149 == array_addr[13:5] | valid_329; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_875 = 9'h14a == array_addr[13:5] | valid_330; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_876 = 9'h14b == array_addr[13:5] | valid_331; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_877 = 9'h14c == array_addr[13:5] | valid_332; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_878 = 9'h14d == array_addr[13:5] | valid_333; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_879 = 9'h14e == array_addr[13:5] | valid_334; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_880 = 9'h14f == array_addr[13:5] | valid_335; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_881 = 9'h150 == array_addr[13:5] | valid_336; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_882 = 9'h151 == array_addr[13:5] | valid_337; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_883 = 9'h152 == array_addr[13:5] | valid_338; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_884 = 9'h153 == array_addr[13:5] | valid_339; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_885 = 9'h154 == array_addr[13:5] | valid_340; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_886 = 9'h155 == array_addr[13:5] | valid_341; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_887 = 9'h156 == array_addr[13:5] | valid_342; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_888 = 9'h157 == array_addr[13:5] | valid_343; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_889 = 9'h158 == array_addr[13:5] | valid_344; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_890 = 9'h159 == array_addr[13:5] | valid_345; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_891 = 9'h15a == array_addr[13:5] | valid_346; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_892 = 9'h15b == array_addr[13:5] | valid_347; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_893 = 9'h15c == array_addr[13:5] | valid_348; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_894 = 9'h15d == array_addr[13:5] | valid_349; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_895 = 9'h15e == array_addr[13:5] | valid_350; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_896 = 9'h15f == array_addr[13:5] | valid_351; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_897 = 9'h160 == array_addr[13:5] | valid_352; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_898 = 9'h161 == array_addr[13:5] | valid_353; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_899 = 9'h162 == array_addr[13:5] | valid_354; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_900 = 9'h163 == array_addr[13:5] | valid_355; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_901 = 9'h164 == array_addr[13:5] | valid_356; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_902 = 9'h165 == array_addr[13:5] | valid_357; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_903 = 9'h166 == array_addr[13:5] | valid_358; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_904 = 9'h167 == array_addr[13:5] | valid_359; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_905 = 9'h168 == array_addr[13:5] | valid_360; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_906 = 9'h169 == array_addr[13:5] | valid_361; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_907 = 9'h16a == array_addr[13:5] | valid_362; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_908 = 9'h16b == array_addr[13:5] | valid_363; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_909 = 9'h16c == array_addr[13:5] | valid_364; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_910 = 9'h16d == array_addr[13:5] | valid_365; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_911 = 9'h16e == array_addr[13:5] | valid_366; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_912 = 9'h16f == array_addr[13:5] | valid_367; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_913 = 9'h170 == array_addr[13:5] | valid_368; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_914 = 9'h171 == array_addr[13:5] | valid_369; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_915 = 9'h172 == array_addr[13:5] | valid_370; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_916 = 9'h173 == array_addr[13:5] | valid_371; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_917 = 9'h174 == array_addr[13:5] | valid_372; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_918 = 9'h175 == array_addr[13:5] | valid_373; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_919 = 9'h176 == array_addr[13:5] | valid_374; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_920 = 9'h177 == array_addr[13:5] | valid_375; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_921 = 9'h178 == array_addr[13:5] | valid_376; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_922 = 9'h179 == array_addr[13:5] | valid_377; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_923 = 9'h17a == array_addr[13:5] | valid_378; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_924 = 9'h17b == array_addr[13:5] | valid_379; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_925 = 9'h17c == array_addr[13:5] | valid_380; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_926 = 9'h17d == array_addr[13:5] | valid_381; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_927 = 9'h17e == array_addr[13:5] | valid_382; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_928 = 9'h17f == array_addr[13:5] | valid_383; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_929 = 9'h180 == array_addr[13:5] | valid_384; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_930 = 9'h181 == array_addr[13:5] | valid_385; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_931 = 9'h182 == array_addr[13:5] | valid_386; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_932 = 9'h183 == array_addr[13:5] | valid_387; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_933 = 9'h184 == array_addr[13:5] | valid_388; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_934 = 9'h185 == array_addr[13:5] | valid_389; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_935 = 9'h186 == array_addr[13:5] | valid_390; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_936 = 9'h187 == array_addr[13:5] | valid_391; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_937 = 9'h188 == array_addr[13:5] | valid_392; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_938 = 9'h189 == array_addr[13:5] | valid_393; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_939 = 9'h18a == array_addr[13:5] | valid_394; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_940 = 9'h18b == array_addr[13:5] | valid_395; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_941 = 9'h18c == array_addr[13:5] | valid_396; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_942 = 9'h18d == array_addr[13:5] | valid_397; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_943 = 9'h18e == array_addr[13:5] | valid_398; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_944 = 9'h18f == array_addr[13:5] | valid_399; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_945 = 9'h190 == array_addr[13:5] | valid_400; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_946 = 9'h191 == array_addr[13:5] | valid_401; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_947 = 9'h192 == array_addr[13:5] | valid_402; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_948 = 9'h193 == array_addr[13:5] | valid_403; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_949 = 9'h194 == array_addr[13:5] | valid_404; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_950 = 9'h195 == array_addr[13:5] | valid_405; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_951 = 9'h196 == array_addr[13:5] | valid_406; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_952 = 9'h197 == array_addr[13:5] | valid_407; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_953 = 9'h198 == array_addr[13:5] | valid_408; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_954 = 9'h199 == array_addr[13:5] | valid_409; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_955 = 9'h19a == array_addr[13:5] | valid_410; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_956 = 9'h19b == array_addr[13:5] | valid_411; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_957 = 9'h19c == array_addr[13:5] | valid_412; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_958 = 9'h19d == array_addr[13:5] | valid_413; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_959 = 9'h19e == array_addr[13:5] | valid_414; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_960 = 9'h19f == array_addr[13:5] | valid_415; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_961 = 9'h1a0 == array_addr[13:5] | valid_416; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_962 = 9'h1a1 == array_addr[13:5] | valid_417; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_963 = 9'h1a2 == array_addr[13:5] | valid_418; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_964 = 9'h1a3 == array_addr[13:5] | valid_419; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_965 = 9'h1a4 == array_addr[13:5] | valid_420; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_966 = 9'h1a5 == array_addr[13:5] | valid_421; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_967 = 9'h1a6 == array_addr[13:5] | valid_422; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_968 = 9'h1a7 == array_addr[13:5] | valid_423; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_969 = 9'h1a8 == array_addr[13:5] | valid_424; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_970 = 9'h1a9 == array_addr[13:5] | valid_425; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_971 = 9'h1aa == array_addr[13:5] | valid_426; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_972 = 9'h1ab == array_addr[13:5] | valid_427; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_973 = 9'h1ac == array_addr[13:5] | valid_428; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_974 = 9'h1ad == array_addr[13:5] | valid_429; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_975 = 9'h1ae == array_addr[13:5] | valid_430; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_976 = 9'h1af == array_addr[13:5] | valid_431; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_977 = 9'h1b0 == array_addr[13:5] | valid_432; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_978 = 9'h1b1 == array_addr[13:5] | valid_433; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_979 = 9'h1b2 == array_addr[13:5] | valid_434; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_980 = 9'h1b3 == array_addr[13:5] | valid_435; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_981 = 9'h1b4 == array_addr[13:5] | valid_436; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_982 = 9'h1b5 == array_addr[13:5] | valid_437; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_983 = 9'h1b6 == array_addr[13:5] | valid_438; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_984 = 9'h1b7 == array_addr[13:5] | valid_439; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_985 = 9'h1b8 == array_addr[13:5] | valid_440; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_986 = 9'h1b9 == array_addr[13:5] | valid_441; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_987 = 9'h1ba == array_addr[13:5] | valid_442; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_988 = 9'h1bb == array_addr[13:5] | valid_443; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_989 = 9'h1bc == array_addr[13:5] | valid_444; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_990 = 9'h1bd == array_addr[13:5] | valid_445; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_991 = 9'h1be == array_addr[13:5] | valid_446; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_992 = 9'h1bf == array_addr[13:5] | valid_447; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_993 = 9'h1c0 == array_addr[13:5] | valid_448; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_994 = 9'h1c1 == array_addr[13:5] | valid_449; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_995 = 9'h1c2 == array_addr[13:5] | valid_450; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_996 = 9'h1c3 == array_addr[13:5] | valid_451; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_997 = 9'h1c4 == array_addr[13:5] | valid_452; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_998 = 9'h1c5 == array_addr[13:5] | valid_453; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_999 = 9'h1c6 == array_addr[13:5] | valid_454; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1000 = 9'h1c7 == array_addr[13:5] | valid_455; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1001 = 9'h1c8 == array_addr[13:5] | valid_456; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1002 = 9'h1c9 == array_addr[13:5] | valid_457; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1003 = 9'h1ca == array_addr[13:5] | valid_458; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1004 = 9'h1cb == array_addr[13:5] | valid_459; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1005 = 9'h1cc == array_addr[13:5] | valid_460; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1006 = 9'h1cd == array_addr[13:5] | valid_461; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1007 = 9'h1ce == array_addr[13:5] | valid_462; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1008 = 9'h1cf == array_addr[13:5] | valid_463; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1009 = 9'h1d0 == array_addr[13:5] | valid_464; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1010 = 9'h1d1 == array_addr[13:5] | valid_465; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1011 = 9'h1d2 == array_addr[13:5] | valid_466; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1012 = 9'h1d3 == array_addr[13:5] | valid_467; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1013 = 9'h1d4 == array_addr[13:5] | valid_468; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1014 = 9'h1d5 == array_addr[13:5] | valid_469; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1015 = 9'h1d6 == array_addr[13:5] | valid_470; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1016 = 9'h1d7 == array_addr[13:5] | valid_471; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1017 = 9'h1d8 == array_addr[13:5] | valid_472; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1018 = 9'h1d9 == array_addr[13:5] | valid_473; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1019 = 9'h1da == array_addr[13:5] | valid_474; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1020 = 9'h1db == array_addr[13:5] | valid_475; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1021 = 9'h1dc == array_addr[13:5] | valid_476; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1022 = 9'h1dd == array_addr[13:5] | valid_477; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1023 = 9'h1de == array_addr[13:5] | valid_478; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1024 = 9'h1df == array_addr[13:5] | valid_479; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1025 = 9'h1e0 == array_addr[13:5] | valid_480; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1026 = 9'h1e1 == array_addr[13:5] | valid_481; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1027 = 9'h1e2 == array_addr[13:5] | valid_482; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1028 = 9'h1e3 == array_addr[13:5] | valid_483; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1029 = 9'h1e4 == array_addr[13:5] | valid_484; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1030 = 9'h1e5 == array_addr[13:5] | valid_485; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1031 = 9'h1e6 == array_addr[13:5] | valid_486; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1032 = 9'h1e7 == array_addr[13:5] | valid_487; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1033 = 9'h1e8 == array_addr[13:5] | valid_488; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1034 = 9'h1e9 == array_addr[13:5] | valid_489; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1035 = 9'h1ea == array_addr[13:5] | valid_490; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1036 = 9'h1eb == array_addr[13:5] | valid_491; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1037 = 9'h1ec == array_addr[13:5] | valid_492; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1038 = 9'h1ed == array_addr[13:5] | valid_493; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1039 = 9'h1ee == array_addr[13:5] | valid_494; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1040 = 9'h1ef == array_addr[13:5] | valid_495; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1041 = 9'h1f0 == array_addr[13:5] | valid_496; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1042 = 9'h1f1 == array_addr[13:5] | valid_497; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1043 = 9'h1f2 == array_addr[13:5] | valid_498; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1044 = 9'h1f3 == array_addr[13:5] | valid_499; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1045 = 9'h1f4 == array_addr[13:5] | valid_500; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1046 = 9'h1f5 == array_addr[13:5] | valid_501; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1047 = 9'h1f6 == array_addr[13:5] | valid_502; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1048 = 9'h1f7 == array_addr[13:5] | valid_503; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1049 = 9'h1f8 == array_addr[13:5] | valid_504; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1050 = 9'h1f9 == array_addr[13:5] | valid_505; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1051 = 9'h1fa == array_addr[13:5] | valid_506; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1052 = 9'h1fb == array_addr[13:5] | valid_507; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1053 = 9'h1fc == array_addr[13:5] | valid_508; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1054 = 9'h1fd == array_addr[13:5] | valid_509; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1055 = 9'h1fe == array_addr[13:5] | valid_510; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1056 = 9'h1ff == array_addr[13:5] | valid_511; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1058 = ~sc_fail_r ? _GEN_545 : valid_0; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1059 = ~sc_fail_r ? _GEN_546 : valid_1; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1060 = ~sc_fail_r ? _GEN_547 : valid_2; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1061 = ~sc_fail_r ? _GEN_548 : valid_3; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1062 = ~sc_fail_r ? _GEN_549 : valid_4; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1063 = ~sc_fail_r ? _GEN_550 : valid_5; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1064 = ~sc_fail_r ? _GEN_551 : valid_6; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1065 = ~sc_fail_r ? _GEN_552 : valid_7; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1066 = ~sc_fail_r ? _GEN_553 : valid_8; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1067 = ~sc_fail_r ? _GEN_554 : valid_9; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1068 = ~sc_fail_r ? _GEN_555 : valid_10; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1069 = ~sc_fail_r ? _GEN_556 : valid_11; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1070 = ~sc_fail_r ? _GEN_557 : valid_12; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1071 = ~sc_fail_r ? _GEN_558 : valid_13; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1072 = ~sc_fail_r ? _GEN_559 : valid_14; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1073 = ~sc_fail_r ? _GEN_560 : valid_15; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1074 = ~sc_fail_r ? _GEN_561 : valid_16; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1075 = ~sc_fail_r ? _GEN_562 : valid_17; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1076 = ~sc_fail_r ? _GEN_563 : valid_18; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1077 = ~sc_fail_r ? _GEN_564 : valid_19; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1078 = ~sc_fail_r ? _GEN_565 : valid_20; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1079 = ~sc_fail_r ? _GEN_566 : valid_21; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1080 = ~sc_fail_r ? _GEN_567 : valid_22; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1081 = ~sc_fail_r ? _GEN_568 : valid_23; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1082 = ~sc_fail_r ? _GEN_569 : valid_24; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1083 = ~sc_fail_r ? _GEN_570 : valid_25; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1084 = ~sc_fail_r ? _GEN_571 : valid_26; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1085 = ~sc_fail_r ? _GEN_572 : valid_27; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1086 = ~sc_fail_r ? _GEN_573 : valid_28; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1087 = ~sc_fail_r ? _GEN_574 : valid_29; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1088 = ~sc_fail_r ? _GEN_575 : valid_30; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1089 = ~sc_fail_r ? _GEN_576 : valid_31; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1090 = ~sc_fail_r ? _GEN_577 : valid_32; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1091 = ~sc_fail_r ? _GEN_578 : valid_33; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1092 = ~sc_fail_r ? _GEN_579 : valid_34; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1093 = ~sc_fail_r ? _GEN_580 : valid_35; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1094 = ~sc_fail_r ? _GEN_581 : valid_36; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1095 = ~sc_fail_r ? _GEN_582 : valid_37; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1096 = ~sc_fail_r ? _GEN_583 : valid_38; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1097 = ~sc_fail_r ? _GEN_584 : valid_39; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1098 = ~sc_fail_r ? _GEN_585 : valid_40; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1099 = ~sc_fail_r ? _GEN_586 : valid_41; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1100 = ~sc_fail_r ? _GEN_587 : valid_42; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1101 = ~sc_fail_r ? _GEN_588 : valid_43; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1102 = ~sc_fail_r ? _GEN_589 : valid_44; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1103 = ~sc_fail_r ? _GEN_590 : valid_45; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1104 = ~sc_fail_r ? _GEN_591 : valid_46; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1105 = ~sc_fail_r ? _GEN_592 : valid_47; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1106 = ~sc_fail_r ? _GEN_593 : valid_48; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1107 = ~sc_fail_r ? _GEN_594 : valid_49; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1108 = ~sc_fail_r ? _GEN_595 : valid_50; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1109 = ~sc_fail_r ? _GEN_596 : valid_51; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1110 = ~sc_fail_r ? _GEN_597 : valid_52; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1111 = ~sc_fail_r ? _GEN_598 : valid_53; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1112 = ~sc_fail_r ? _GEN_599 : valid_54; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1113 = ~sc_fail_r ? _GEN_600 : valid_55; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1114 = ~sc_fail_r ? _GEN_601 : valid_56; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1115 = ~sc_fail_r ? _GEN_602 : valid_57; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1116 = ~sc_fail_r ? _GEN_603 : valid_58; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1117 = ~sc_fail_r ? _GEN_604 : valid_59; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1118 = ~sc_fail_r ? _GEN_605 : valid_60; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1119 = ~sc_fail_r ? _GEN_606 : valid_61; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1120 = ~sc_fail_r ? _GEN_607 : valid_62; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1121 = ~sc_fail_r ? _GEN_608 : valid_63; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1122 = ~sc_fail_r ? _GEN_609 : valid_64; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1123 = ~sc_fail_r ? _GEN_610 : valid_65; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1124 = ~sc_fail_r ? _GEN_611 : valid_66; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1125 = ~sc_fail_r ? _GEN_612 : valid_67; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1126 = ~sc_fail_r ? _GEN_613 : valid_68; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1127 = ~sc_fail_r ? _GEN_614 : valid_69; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1128 = ~sc_fail_r ? _GEN_615 : valid_70; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1129 = ~sc_fail_r ? _GEN_616 : valid_71; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1130 = ~sc_fail_r ? _GEN_617 : valid_72; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1131 = ~sc_fail_r ? _GEN_618 : valid_73; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1132 = ~sc_fail_r ? _GEN_619 : valid_74; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1133 = ~sc_fail_r ? _GEN_620 : valid_75; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1134 = ~sc_fail_r ? _GEN_621 : valid_76; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1135 = ~sc_fail_r ? _GEN_622 : valid_77; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1136 = ~sc_fail_r ? _GEN_623 : valid_78; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1137 = ~sc_fail_r ? _GEN_624 : valid_79; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1138 = ~sc_fail_r ? _GEN_625 : valid_80; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1139 = ~sc_fail_r ? _GEN_626 : valid_81; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1140 = ~sc_fail_r ? _GEN_627 : valid_82; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1141 = ~sc_fail_r ? _GEN_628 : valid_83; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1142 = ~sc_fail_r ? _GEN_629 : valid_84; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1143 = ~sc_fail_r ? _GEN_630 : valid_85; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1144 = ~sc_fail_r ? _GEN_631 : valid_86; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1145 = ~sc_fail_r ? _GEN_632 : valid_87; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1146 = ~sc_fail_r ? _GEN_633 : valid_88; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1147 = ~sc_fail_r ? _GEN_634 : valid_89; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1148 = ~sc_fail_r ? _GEN_635 : valid_90; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1149 = ~sc_fail_r ? _GEN_636 : valid_91; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1150 = ~sc_fail_r ? _GEN_637 : valid_92; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1151 = ~sc_fail_r ? _GEN_638 : valid_93; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1152 = ~sc_fail_r ? _GEN_639 : valid_94; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1153 = ~sc_fail_r ? _GEN_640 : valid_95; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1154 = ~sc_fail_r ? _GEN_641 : valid_96; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1155 = ~sc_fail_r ? _GEN_642 : valid_97; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1156 = ~sc_fail_r ? _GEN_643 : valid_98; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1157 = ~sc_fail_r ? _GEN_644 : valid_99; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1158 = ~sc_fail_r ? _GEN_645 : valid_100; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1159 = ~sc_fail_r ? _GEN_646 : valid_101; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1160 = ~sc_fail_r ? _GEN_647 : valid_102; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1161 = ~sc_fail_r ? _GEN_648 : valid_103; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1162 = ~sc_fail_r ? _GEN_649 : valid_104; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1163 = ~sc_fail_r ? _GEN_650 : valid_105; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1164 = ~sc_fail_r ? _GEN_651 : valid_106; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1165 = ~sc_fail_r ? _GEN_652 : valid_107; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1166 = ~sc_fail_r ? _GEN_653 : valid_108; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1167 = ~sc_fail_r ? _GEN_654 : valid_109; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1168 = ~sc_fail_r ? _GEN_655 : valid_110; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1169 = ~sc_fail_r ? _GEN_656 : valid_111; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1170 = ~sc_fail_r ? _GEN_657 : valid_112; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1171 = ~sc_fail_r ? _GEN_658 : valid_113; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1172 = ~sc_fail_r ? _GEN_659 : valid_114; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1173 = ~sc_fail_r ? _GEN_660 : valid_115; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1174 = ~sc_fail_r ? _GEN_661 : valid_116; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1175 = ~sc_fail_r ? _GEN_662 : valid_117; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1176 = ~sc_fail_r ? _GEN_663 : valid_118; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1177 = ~sc_fail_r ? _GEN_664 : valid_119; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1178 = ~sc_fail_r ? _GEN_665 : valid_120; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1179 = ~sc_fail_r ? _GEN_666 : valid_121; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1180 = ~sc_fail_r ? _GEN_667 : valid_122; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1181 = ~sc_fail_r ? _GEN_668 : valid_123; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1182 = ~sc_fail_r ? _GEN_669 : valid_124; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1183 = ~sc_fail_r ? _GEN_670 : valid_125; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1184 = ~sc_fail_r ? _GEN_671 : valid_126; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1185 = ~sc_fail_r ? _GEN_672 : valid_127; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1186 = ~sc_fail_r ? _GEN_673 : valid_128; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1187 = ~sc_fail_r ? _GEN_674 : valid_129; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1188 = ~sc_fail_r ? _GEN_675 : valid_130; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1189 = ~sc_fail_r ? _GEN_676 : valid_131; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1190 = ~sc_fail_r ? _GEN_677 : valid_132; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1191 = ~sc_fail_r ? _GEN_678 : valid_133; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1192 = ~sc_fail_r ? _GEN_679 : valid_134; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1193 = ~sc_fail_r ? _GEN_680 : valid_135; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1194 = ~sc_fail_r ? _GEN_681 : valid_136; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1195 = ~sc_fail_r ? _GEN_682 : valid_137; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1196 = ~sc_fail_r ? _GEN_683 : valid_138; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1197 = ~sc_fail_r ? _GEN_684 : valid_139; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1198 = ~sc_fail_r ? _GEN_685 : valid_140; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1199 = ~sc_fail_r ? _GEN_686 : valid_141; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1200 = ~sc_fail_r ? _GEN_687 : valid_142; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1201 = ~sc_fail_r ? _GEN_688 : valid_143; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1202 = ~sc_fail_r ? _GEN_689 : valid_144; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1203 = ~sc_fail_r ? _GEN_690 : valid_145; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1204 = ~sc_fail_r ? _GEN_691 : valid_146; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1205 = ~sc_fail_r ? _GEN_692 : valid_147; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1206 = ~sc_fail_r ? _GEN_693 : valid_148; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1207 = ~sc_fail_r ? _GEN_694 : valid_149; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1208 = ~sc_fail_r ? _GEN_695 : valid_150; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1209 = ~sc_fail_r ? _GEN_696 : valid_151; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1210 = ~sc_fail_r ? _GEN_697 : valid_152; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1211 = ~sc_fail_r ? _GEN_698 : valid_153; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1212 = ~sc_fail_r ? _GEN_699 : valid_154; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1213 = ~sc_fail_r ? _GEN_700 : valid_155; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1214 = ~sc_fail_r ? _GEN_701 : valid_156; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1215 = ~sc_fail_r ? _GEN_702 : valid_157; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1216 = ~sc_fail_r ? _GEN_703 : valid_158; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1217 = ~sc_fail_r ? _GEN_704 : valid_159; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1218 = ~sc_fail_r ? _GEN_705 : valid_160; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1219 = ~sc_fail_r ? _GEN_706 : valid_161; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1220 = ~sc_fail_r ? _GEN_707 : valid_162; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1221 = ~sc_fail_r ? _GEN_708 : valid_163; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1222 = ~sc_fail_r ? _GEN_709 : valid_164; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1223 = ~sc_fail_r ? _GEN_710 : valid_165; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1224 = ~sc_fail_r ? _GEN_711 : valid_166; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1225 = ~sc_fail_r ? _GEN_712 : valid_167; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1226 = ~sc_fail_r ? _GEN_713 : valid_168; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1227 = ~sc_fail_r ? _GEN_714 : valid_169; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1228 = ~sc_fail_r ? _GEN_715 : valid_170; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1229 = ~sc_fail_r ? _GEN_716 : valid_171; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1230 = ~sc_fail_r ? _GEN_717 : valid_172; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1231 = ~sc_fail_r ? _GEN_718 : valid_173; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1232 = ~sc_fail_r ? _GEN_719 : valid_174; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1233 = ~sc_fail_r ? _GEN_720 : valid_175; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1234 = ~sc_fail_r ? _GEN_721 : valid_176; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1235 = ~sc_fail_r ? _GEN_722 : valid_177; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1236 = ~sc_fail_r ? _GEN_723 : valid_178; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1237 = ~sc_fail_r ? _GEN_724 : valid_179; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1238 = ~sc_fail_r ? _GEN_725 : valid_180; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1239 = ~sc_fail_r ? _GEN_726 : valid_181; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1240 = ~sc_fail_r ? _GEN_727 : valid_182; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1241 = ~sc_fail_r ? _GEN_728 : valid_183; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1242 = ~sc_fail_r ? _GEN_729 : valid_184; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1243 = ~sc_fail_r ? _GEN_730 : valid_185; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1244 = ~sc_fail_r ? _GEN_731 : valid_186; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1245 = ~sc_fail_r ? _GEN_732 : valid_187; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1246 = ~sc_fail_r ? _GEN_733 : valid_188; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1247 = ~sc_fail_r ? _GEN_734 : valid_189; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1248 = ~sc_fail_r ? _GEN_735 : valid_190; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1249 = ~sc_fail_r ? _GEN_736 : valid_191; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1250 = ~sc_fail_r ? _GEN_737 : valid_192; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1251 = ~sc_fail_r ? _GEN_738 : valid_193; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1252 = ~sc_fail_r ? _GEN_739 : valid_194; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1253 = ~sc_fail_r ? _GEN_740 : valid_195; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1254 = ~sc_fail_r ? _GEN_741 : valid_196; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1255 = ~sc_fail_r ? _GEN_742 : valid_197; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1256 = ~sc_fail_r ? _GEN_743 : valid_198; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1257 = ~sc_fail_r ? _GEN_744 : valid_199; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1258 = ~sc_fail_r ? _GEN_745 : valid_200; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1259 = ~sc_fail_r ? _GEN_746 : valid_201; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1260 = ~sc_fail_r ? _GEN_747 : valid_202; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1261 = ~sc_fail_r ? _GEN_748 : valid_203; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1262 = ~sc_fail_r ? _GEN_749 : valid_204; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1263 = ~sc_fail_r ? _GEN_750 : valid_205; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1264 = ~sc_fail_r ? _GEN_751 : valid_206; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1265 = ~sc_fail_r ? _GEN_752 : valid_207; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1266 = ~sc_fail_r ? _GEN_753 : valid_208; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1267 = ~sc_fail_r ? _GEN_754 : valid_209; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1268 = ~sc_fail_r ? _GEN_755 : valid_210; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1269 = ~sc_fail_r ? _GEN_756 : valid_211; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1270 = ~sc_fail_r ? _GEN_757 : valid_212; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1271 = ~sc_fail_r ? _GEN_758 : valid_213; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1272 = ~sc_fail_r ? _GEN_759 : valid_214; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1273 = ~sc_fail_r ? _GEN_760 : valid_215; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1274 = ~sc_fail_r ? _GEN_761 : valid_216; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1275 = ~sc_fail_r ? _GEN_762 : valid_217; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1276 = ~sc_fail_r ? _GEN_763 : valid_218; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1277 = ~sc_fail_r ? _GEN_764 : valid_219; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1278 = ~sc_fail_r ? _GEN_765 : valid_220; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1279 = ~sc_fail_r ? _GEN_766 : valid_221; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1280 = ~sc_fail_r ? _GEN_767 : valid_222; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1281 = ~sc_fail_r ? _GEN_768 : valid_223; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1282 = ~sc_fail_r ? _GEN_769 : valid_224; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1283 = ~sc_fail_r ? _GEN_770 : valid_225; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1284 = ~sc_fail_r ? _GEN_771 : valid_226; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1285 = ~sc_fail_r ? _GEN_772 : valid_227; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1286 = ~sc_fail_r ? _GEN_773 : valid_228; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1287 = ~sc_fail_r ? _GEN_774 : valid_229; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1288 = ~sc_fail_r ? _GEN_775 : valid_230; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1289 = ~sc_fail_r ? _GEN_776 : valid_231; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1290 = ~sc_fail_r ? _GEN_777 : valid_232; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1291 = ~sc_fail_r ? _GEN_778 : valid_233; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1292 = ~sc_fail_r ? _GEN_779 : valid_234; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1293 = ~sc_fail_r ? _GEN_780 : valid_235; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1294 = ~sc_fail_r ? _GEN_781 : valid_236; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1295 = ~sc_fail_r ? _GEN_782 : valid_237; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1296 = ~sc_fail_r ? _GEN_783 : valid_238; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1297 = ~sc_fail_r ? _GEN_784 : valid_239; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1298 = ~sc_fail_r ? _GEN_785 : valid_240; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1299 = ~sc_fail_r ? _GEN_786 : valid_241; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1300 = ~sc_fail_r ? _GEN_787 : valid_242; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1301 = ~sc_fail_r ? _GEN_788 : valid_243; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1302 = ~sc_fail_r ? _GEN_789 : valid_244; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1303 = ~sc_fail_r ? _GEN_790 : valid_245; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1304 = ~sc_fail_r ? _GEN_791 : valid_246; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1305 = ~sc_fail_r ? _GEN_792 : valid_247; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1306 = ~sc_fail_r ? _GEN_793 : valid_248; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1307 = ~sc_fail_r ? _GEN_794 : valid_249; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1308 = ~sc_fail_r ? _GEN_795 : valid_250; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1309 = ~sc_fail_r ? _GEN_796 : valid_251; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1310 = ~sc_fail_r ? _GEN_797 : valid_252; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1311 = ~sc_fail_r ? _GEN_798 : valid_253; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1312 = ~sc_fail_r ? _GEN_799 : valid_254; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1313 = ~sc_fail_r ? _GEN_800 : valid_255; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1314 = ~sc_fail_r ? _GEN_801 : valid_256; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1315 = ~sc_fail_r ? _GEN_802 : valid_257; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1316 = ~sc_fail_r ? _GEN_803 : valid_258; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1317 = ~sc_fail_r ? _GEN_804 : valid_259; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1318 = ~sc_fail_r ? _GEN_805 : valid_260; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1319 = ~sc_fail_r ? _GEN_806 : valid_261; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1320 = ~sc_fail_r ? _GEN_807 : valid_262; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1321 = ~sc_fail_r ? _GEN_808 : valid_263; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1322 = ~sc_fail_r ? _GEN_809 : valid_264; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1323 = ~sc_fail_r ? _GEN_810 : valid_265; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1324 = ~sc_fail_r ? _GEN_811 : valid_266; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1325 = ~sc_fail_r ? _GEN_812 : valid_267; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1326 = ~sc_fail_r ? _GEN_813 : valid_268; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1327 = ~sc_fail_r ? _GEN_814 : valid_269; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1328 = ~sc_fail_r ? _GEN_815 : valid_270; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1329 = ~sc_fail_r ? _GEN_816 : valid_271; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1330 = ~sc_fail_r ? _GEN_817 : valid_272; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1331 = ~sc_fail_r ? _GEN_818 : valid_273; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1332 = ~sc_fail_r ? _GEN_819 : valid_274; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1333 = ~sc_fail_r ? _GEN_820 : valid_275; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1334 = ~sc_fail_r ? _GEN_821 : valid_276; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1335 = ~sc_fail_r ? _GEN_822 : valid_277; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1336 = ~sc_fail_r ? _GEN_823 : valid_278; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1337 = ~sc_fail_r ? _GEN_824 : valid_279; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1338 = ~sc_fail_r ? _GEN_825 : valid_280; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1339 = ~sc_fail_r ? _GEN_826 : valid_281; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1340 = ~sc_fail_r ? _GEN_827 : valid_282; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1341 = ~sc_fail_r ? _GEN_828 : valid_283; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1342 = ~sc_fail_r ? _GEN_829 : valid_284; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1343 = ~sc_fail_r ? _GEN_830 : valid_285; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1344 = ~sc_fail_r ? _GEN_831 : valid_286; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1345 = ~sc_fail_r ? _GEN_832 : valid_287; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1346 = ~sc_fail_r ? _GEN_833 : valid_288; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1347 = ~sc_fail_r ? _GEN_834 : valid_289; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1348 = ~sc_fail_r ? _GEN_835 : valid_290; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1349 = ~sc_fail_r ? _GEN_836 : valid_291; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1350 = ~sc_fail_r ? _GEN_837 : valid_292; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1351 = ~sc_fail_r ? _GEN_838 : valid_293; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1352 = ~sc_fail_r ? _GEN_839 : valid_294; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1353 = ~sc_fail_r ? _GEN_840 : valid_295; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1354 = ~sc_fail_r ? _GEN_841 : valid_296; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1355 = ~sc_fail_r ? _GEN_842 : valid_297; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1356 = ~sc_fail_r ? _GEN_843 : valid_298; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1357 = ~sc_fail_r ? _GEN_844 : valid_299; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1358 = ~sc_fail_r ? _GEN_845 : valid_300; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1359 = ~sc_fail_r ? _GEN_846 : valid_301; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1360 = ~sc_fail_r ? _GEN_847 : valid_302; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1361 = ~sc_fail_r ? _GEN_848 : valid_303; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1362 = ~sc_fail_r ? _GEN_849 : valid_304; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1363 = ~sc_fail_r ? _GEN_850 : valid_305; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1364 = ~sc_fail_r ? _GEN_851 : valid_306; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1365 = ~sc_fail_r ? _GEN_852 : valid_307; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1366 = ~sc_fail_r ? _GEN_853 : valid_308; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1367 = ~sc_fail_r ? _GEN_854 : valid_309; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1368 = ~sc_fail_r ? _GEN_855 : valid_310; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1369 = ~sc_fail_r ? _GEN_856 : valid_311; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1370 = ~sc_fail_r ? _GEN_857 : valid_312; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1371 = ~sc_fail_r ? _GEN_858 : valid_313; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1372 = ~sc_fail_r ? _GEN_859 : valid_314; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1373 = ~sc_fail_r ? _GEN_860 : valid_315; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1374 = ~sc_fail_r ? _GEN_861 : valid_316; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1375 = ~sc_fail_r ? _GEN_862 : valid_317; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1376 = ~sc_fail_r ? _GEN_863 : valid_318; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1377 = ~sc_fail_r ? _GEN_864 : valid_319; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1378 = ~sc_fail_r ? _GEN_865 : valid_320; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1379 = ~sc_fail_r ? _GEN_866 : valid_321; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1380 = ~sc_fail_r ? _GEN_867 : valid_322; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1381 = ~sc_fail_r ? _GEN_868 : valid_323; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1382 = ~sc_fail_r ? _GEN_869 : valid_324; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1383 = ~sc_fail_r ? _GEN_870 : valid_325; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1384 = ~sc_fail_r ? _GEN_871 : valid_326; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1385 = ~sc_fail_r ? _GEN_872 : valid_327; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1386 = ~sc_fail_r ? _GEN_873 : valid_328; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1387 = ~sc_fail_r ? _GEN_874 : valid_329; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1388 = ~sc_fail_r ? _GEN_875 : valid_330; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1389 = ~sc_fail_r ? _GEN_876 : valid_331; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1390 = ~sc_fail_r ? _GEN_877 : valid_332; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1391 = ~sc_fail_r ? _GEN_878 : valid_333; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1392 = ~sc_fail_r ? _GEN_879 : valid_334; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1393 = ~sc_fail_r ? _GEN_880 : valid_335; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1394 = ~sc_fail_r ? _GEN_881 : valid_336; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1395 = ~sc_fail_r ? _GEN_882 : valid_337; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1396 = ~sc_fail_r ? _GEN_883 : valid_338; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1397 = ~sc_fail_r ? _GEN_884 : valid_339; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1398 = ~sc_fail_r ? _GEN_885 : valid_340; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1399 = ~sc_fail_r ? _GEN_886 : valid_341; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1400 = ~sc_fail_r ? _GEN_887 : valid_342; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1401 = ~sc_fail_r ? _GEN_888 : valid_343; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1402 = ~sc_fail_r ? _GEN_889 : valid_344; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1403 = ~sc_fail_r ? _GEN_890 : valid_345; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1404 = ~sc_fail_r ? _GEN_891 : valid_346; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1405 = ~sc_fail_r ? _GEN_892 : valid_347; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1406 = ~sc_fail_r ? _GEN_893 : valid_348; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1407 = ~sc_fail_r ? _GEN_894 : valid_349; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1408 = ~sc_fail_r ? _GEN_895 : valid_350; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1409 = ~sc_fail_r ? _GEN_896 : valid_351; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1410 = ~sc_fail_r ? _GEN_897 : valid_352; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1411 = ~sc_fail_r ? _GEN_898 : valid_353; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1412 = ~sc_fail_r ? _GEN_899 : valid_354; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1413 = ~sc_fail_r ? _GEN_900 : valid_355; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1414 = ~sc_fail_r ? _GEN_901 : valid_356; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1415 = ~sc_fail_r ? _GEN_902 : valid_357; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1416 = ~sc_fail_r ? _GEN_903 : valid_358; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1417 = ~sc_fail_r ? _GEN_904 : valid_359; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1418 = ~sc_fail_r ? _GEN_905 : valid_360; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1419 = ~sc_fail_r ? _GEN_906 : valid_361; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1420 = ~sc_fail_r ? _GEN_907 : valid_362; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1421 = ~sc_fail_r ? _GEN_908 : valid_363; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1422 = ~sc_fail_r ? _GEN_909 : valid_364; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1423 = ~sc_fail_r ? _GEN_910 : valid_365; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1424 = ~sc_fail_r ? _GEN_911 : valid_366; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1425 = ~sc_fail_r ? _GEN_912 : valid_367; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1426 = ~sc_fail_r ? _GEN_913 : valid_368; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1427 = ~sc_fail_r ? _GEN_914 : valid_369; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1428 = ~sc_fail_r ? _GEN_915 : valid_370; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1429 = ~sc_fail_r ? _GEN_916 : valid_371; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1430 = ~sc_fail_r ? _GEN_917 : valid_372; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1431 = ~sc_fail_r ? _GEN_918 : valid_373; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1432 = ~sc_fail_r ? _GEN_919 : valid_374; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1433 = ~sc_fail_r ? _GEN_920 : valid_375; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1434 = ~sc_fail_r ? _GEN_921 : valid_376; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1435 = ~sc_fail_r ? _GEN_922 : valid_377; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1436 = ~sc_fail_r ? _GEN_923 : valid_378; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1437 = ~sc_fail_r ? _GEN_924 : valid_379; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1438 = ~sc_fail_r ? _GEN_925 : valid_380; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1439 = ~sc_fail_r ? _GEN_926 : valid_381; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1440 = ~sc_fail_r ? _GEN_927 : valid_382; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1441 = ~sc_fail_r ? _GEN_928 : valid_383; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1442 = ~sc_fail_r ? _GEN_929 : valid_384; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1443 = ~sc_fail_r ? _GEN_930 : valid_385; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1444 = ~sc_fail_r ? _GEN_931 : valid_386; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1445 = ~sc_fail_r ? _GEN_932 : valid_387; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1446 = ~sc_fail_r ? _GEN_933 : valid_388; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1447 = ~sc_fail_r ? _GEN_934 : valid_389; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1448 = ~sc_fail_r ? _GEN_935 : valid_390; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1449 = ~sc_fail_r ? _GEN_936 : valid_391; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1450 = ~sc_fail_r ? _GEN_937 : valid_392; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1451 = ~sc_fail_r ? _GEN_938 : valid_393; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1452 = ~sc_fail_r ? _GEN_939 : valid_394; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1453 = ~sc_fail_r ? _GEN_940 : valid_395; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1454 = ~sc_fail_r ? _GEN_941 : valid_396; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1455 = ~sc_fail_r ? _GEN_942 : valid_397; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1456 = ~sc_fail_r ? _GEN_943 : valid_398; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1457 = ~sc_fail_r ? _GEN_944 : valid_399; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1458 = ~sc_fail_r ? _GEN_945 : valid_400; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1459 = ~sc_fail_r ? _GEN_946 : valid_401; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1460 = ~sc_fail_r ? _GEN_947 : valid_402; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1461 = ~sc_fail_r ? _GEN_948 : valid_403; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1462 = ~sc_fail_r ? _GEN_949 : valid_404; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1463 = ~sc_fail_r ? _GEN_950 : valid_405; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1464 = ~sc_fail_r ? _GEN_951 : valid_406; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1465 = ~sc_fail_r ? _GEN_952 : valid_407; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1466 = ~sc_fail_r ? _GEN_953 : valid_408; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1467 = ~sc_fail_r ? _GEN_954 : valid_409; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1468 = ~sc_fail_r ? _GEN_955 : valid_410; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1469 = ~sc_fail_r ? _GEN_956 : valid_411; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1470 = ~sc_fail_r ? _GEN_957 : valid_412; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1471 = ~sc_fail_r ? _GEN_958 : valid_413; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1472 = ~sc_fail_r ? _GEN_959 : valid_414; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1473 = ~sc_fail_r ? _GEN_960 : valid_415; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1474 = ~sc_fail_r ? _GEN_961 : valid_416; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1475 = ~sc_fail_r ? _GEN_962 : valid_417; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1476 = ~sc_fail_r ? _GEN_963 : valid_418; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1477 = ~sc_fail_r ? _GEN_964 : valid_419; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1478 = ~sc_fail_r ? _GEN_965 : valid_420; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1479 = ~sc_fail_r ? _GEN_966 : valid_421; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1480 = ~sc_fail_r ? _GEN_967 : valid_422; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1481 = ~sc_fail_r ? _GEN_968 : valid_423; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1482 = ~sc_fail_r ? _GEN_969 : valid_424; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1483 = ~sc_fail_r ? _GEN_970 : valid_425; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1484 = ~sc_fail_r ? _GEN_971 : valid_426; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1485 = ~sc_fail_r ? _GEN_972 : valid_427; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1486 = ~sc_fail_r ? _GEN_973 : valid_428; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1487 = ~sc_fail_r ? _GEN_974 : valid_429; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1488 = ~sc_fail_r ? _GEN_975 : valid_430; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1489 = ~sc_fail_r ? _GEN_976 : valid_431; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1490 = ~sc_fail_r ? _GEN_977 : valid_432; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1491 = ~sc_fail_r ? _GEN_978 : valid_433; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1492 = ~sc_fail_r ? _GEN_979 : valid_434; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1493 = ~sc_fail_r ? _GEN_980 : valid_435; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1494 = ~sc_fail_r ? _GEN_981 : valid_436; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1495 = ~sc_fail_r ? _GEN_982 : valid_437; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1496 = ~sc_fail_r ? _GEN_983 : valid_438; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1497 = ~sc_fail_r ? _GEN_984 : valid_439; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1498 = ~sc_fail_r ? _GEN_985 : valid_440; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1499 = ~sc_fail_r ? _GEN_986 : valid_441; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1500 = ~sc_fail_r ? _GEN_987 : valid_442; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1501 = ~sc_fail_r ? _GEN_988 : valid_443; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1502 = ~sc_fail_r ? _GEN_989 : valid_444; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1503 = ~sc_fail_r ? _GEN_990 : valid_445; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1504 = ~sc_fail_r ? _GEN_991 : valid_446; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1505 = ~sc_fail_r ? _GEN_992 : valid_447; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1506 = ~sc_fail_r ? _GEN_993 : valid_448; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1507 = ~sc_fail_r ? _GEN_994 : valid_449; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1508 = ~sc_fail_r ? _GEN_995 : valid_450; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1509 = ~sc_fail_r ? _GEN_996 : valid_451; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1510 = ~sc_fail_r ? _GEN_997 : valid_452; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1511 = ~sc_fail_r ? _GEN_998 : valid_453; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1512 = ~sc_fail_r ? _GEN_999 : valid_454; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1513 = ~sc_fail_r ? _GEN_1000 : valid_455; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1514 = ~sc_fail_r ? _GEN_1001 : valid_456; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1515 = ~sc_fail_r ? _GEN_1002 : valid_457; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1516 = ~sc_fail_r ? _GEN_1003 : valid_458; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1517 = ~sc_fail_r ? _GEN_1004 : valid_459; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1518 = ~sc_fail_r ? _GEN_1005 : valid_460; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1519 = ~sc_fail_r ? _GEN_1006 : valid_461; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1520 = ~sc_fail_r ? _GEN_1007 : valid_462; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1521 = ~sc_fail_r ? _GEN_1008 : valid_463; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1522 = ~sc_fail_r ? _GEN_1009 : valid_464; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1523 = ~sc_fail_r ? _GEN_1010 : valid_465; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1524 = ~sc_fail_r ? _GEN_1011 : valid_466; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1525 = ~sc_fail_r ? _GEN_1012 : valid_467; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1526 = ~sc_fail_r ? _GEN_1013 : valid_468; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1527 = ~sc_fail_r ? _GEN_1014 : valid_469; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1528 = ~sc_fail_r ? _GEN_1015 : valid_470; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1529 = ~sc_fail_r ? _GEN_1016 : valid_471; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1530 = ~sc_fail_r ? _GEN_1017 : valid_472; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1531 = ~sc_fail_r ? _GEN_1018 : valid_473; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1532 = ~sc_fail_r ? _GEN_1019 : valid_474; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1533 = ~sc_fail_r ? _GEN_1020 : valid_475; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1534 = ~sc_fail_r ? _GEN_1021 : valid_476; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1535 = ~sc_fail_r ? _GEN_1022 : valid_477; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1536 = ~sc_fail_r ? _GEN_1023 : valid_478; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1537 = ~sc_fail_r ? _GEN_1024 : valid_479; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1538 = ~sc_fail_r ? _GEN_1025 : valid_480; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1539 = ~sc_fail_r ? _GEN_1026 : valid_481; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1540 = ~sc_fail_r ? _GEN_1027 : valid_482; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1541 = ~sc_fail_r ? _GEN_1028 : valid_483; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1542 = ~sc_fail_r ? _GEN_1029 : valid_484; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1543 = ~sc_fail_r ? _GEN_1030 : valid_485; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1544 = ~sc_fail_r ? _GEN_1031 : valid_486; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1545 = ~sc_fail_r ? _GEN_1032 : valid_487; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1546 = ~sc_fail_r ? _GEN_1033 : valid_488; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1547 = ~sc_fail_r ? _GEN_1034 : valid_489; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1548 = ~sc_fail_r ? _GEN_1035 : valid_490; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1549 = ~sc_fail_r ? _GEN_1036 : valid_491; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1550 = ~sc_fail_r ? _GEN_1037 : valid_492; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1551 = ~sc_fail_r ? _GEN_1038 : valid_493; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1552 = ~sc_fail_r ? _GEN_1039 : valid_494; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1553 = ~sc_fail_r ? _GEN_1040 : valid_495; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1554 = ~sc_fail_r ? _GEN_1041 : valid_496; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1555 = ~sc_fail_r ? _GEN_1042 : valid_497; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1556 = ~sc_fail_r ? _GEN_1043 : valid_498; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1557 = ~sc_fail_r ? _GEN_1044 : valid_499; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1558 = ~sc_fail_r ? _GEN_1045 : valid_500; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1559 = ~sc_fail_r ? _GEN_1046 : valid_501; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1560 = ~sc_fail_r ? _GEN_1047 : valid_502; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1561 = ~sc_fail_r ? _GEN_1048 : valid_503; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1562 = ~sc_fail_r ? _GEN_1049 : valid_504; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1563 = ~sc_fail_r ? _GEN_1050 : valid_505; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1564 = ~sc_fail_r ? _GEN_1051 : valid_506; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1565 = ~sc_fail_r ? _GEN_1052 : valid_507; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1566 = ~sc_fail_r ? _GEN_1053 : valid_508; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1567 = ~sc_fail_r ? _GEN_1054 : valid_509; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1568 = ~sc_fail_r ? _GEN_1055 : valid_510; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1569 = ~sc_fail_r ? _GEN_1056 : valid_511; // @[DCache.scala 171:24 56:22]
  wire  _GEN_1571 = state == 3'h7 ? _T_12 : req_r_wen & array_hit; // @[DCache.scala 165:26 177:24]
  wire  _GEN_1572 = state == 3'h7 ? _GEN_1058 : valid_0; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1573 = state == 3'h7 ? _GEN_1059 : valid_1; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1574 = state == 3'h7 ? _GEN_1060 : valid_2; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1575 = state == 3'h7 ? _GEN_1061 : valid_3; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1576 = state == 3'h7 ? _GEN_1062 : valid_4; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1577 = state == 3'h7 ? _GEN_1063 : valid_5; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1578 = state == 3'h7 ? _GEN_1064 : valid_6; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1579 = state == 3'h7 ? _GEN_1065 : valid_7; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1580 = state == 3'h7 ? _GEN_1066 : valid_8; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1581 = state == 3'h7 ? _GEN_1067 : valid_9; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1582 = state == 3'h7 ? _GEN_1068 : valid_10; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1583 = state == 3'h7 ? _GEN_1069 : valid_11; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1584 = state == 3'h7 ? _GEN_1070 : valid_12; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1585 = state == 3'h7 ? _GEN_1071 : valid_13; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1586 = state == 3'h7 ? _GEN_1072 : valid_14; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1587 = state == 3'h7 ? _GEN_1073 : valid_15; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1588 = state == 3'h7 ? _GEN_1074 : valid_16; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1589 = state == 3'h7 ? _GEN_1075 : valid_17; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1590 = state == 3'h7 ? _GEN_1076 : valid_18; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1591 = state == 3'h7 ? _GEN_1077 : valid_19; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1592 = state == 3'h7 ? _GEN_1078 : valid_20; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1593 = state == 3'h7 ? _GEN_1079 : valid_21; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1594 = state == 3'h7 ? _GEN_1080 : valid_22; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1595 = state == 3'h7 ? _GEN_1081 : valid_23; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1596 = state == 3'h7 ? _GEN_1082 : valid_24; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1597 = state == 3'h7 ? _GEN_1083 : valid_25; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1598 = state == 3'h7 ? _GEN_1084 : valid_26; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1599 = state == 3'h7 ? _GEN_1085 : valid_27; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1600 = state == 3'h7 ? _GEN_1086 : valid_28; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1601 = state == 3'h7 ? _GEN_1087 : valid_29; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1602 = state == 3'h7 ? _GEN_1088 : valid_30; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1603 = state == 3'h7 ? _GEN_1089 : valid_31; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1604 = state == 3'h7 ? _GEN_1090 : valid_32; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1605 = state == 3'h7 ? _GEN_1091 : valid_33; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1606 = state == 3'h7 ? _GEN_1092 : valid_34; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1607 = state == 3'h7 ? _GEN_1093 : valid_35; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1608 = state == 3'h7 ? _GEN_1094 : valid_36; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1609 = state == 3'h7 ? _GEN_1095 : valid_37; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1610 = state == 3'h7 ? _GEN_1096 : valid_38; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1611 = state == 3'h7 ? _GEN_1097 : valid_39; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1612 = state == 3'h7 ? _GEN_1098 : valid_40; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1613 = state == 3'h7 ? _GEN_1099 : valid_41; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1614 = state == 3'h7 ? _GEN_1100 : valid_42; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1615 = state == 3'h7 ? _GEN_1101 : valid_43; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1616 = state == 3'h7 ? _GEN_1102 : valid_44; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1617 = state == 3'h7 ? _GEN_1103 : valid_45; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1618 = state == 3'h7 ? _GEN_1104 : valid_46; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1619 = state == 3'h7 ? _GEN_1105 : valid_47; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1620 = state == 3'h7 ? _GEN_1106 : valid_48; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1621 = state == 3'h7 ? _GEN_1107 : valid_49; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1622 = state == 3'h7 ? _GEN_1108 : valid_50; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1623 = state == 3'h7 ? _GEN_1109 : valid_51; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1624 = state == 3'h7 ? _GEN_1110 : valid_52; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1625 = state == 3'h7 ? _GEN_1111 : valid_53; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1626 = state == 3'h7 ? _GEN_1112 : valid_54; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1627 = state == 3'h7 ? _GEN_1113 : valid_55; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1628 = state == 3'h7 ? _GEN_1114 : valid_56; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1629 = state == 3'h7 ? _GEN_1115 : valid_57; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1630 = state == 3'h7 ? _GEN_1116 : valid_58; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1631 = state == 3'h7 ? _GEN_1117 : valid_59; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1632 = state == 3'h7 ? _GEN_1118 : valid_60; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1633 = state == 3'h7 ? _GEN_1119 : valid_61; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1634 = state == 3'h7 ? _GEN_1120 : valid_62; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1635 = state == 3'h7 ? _GEN_1121 : valid_63; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1636 = state == 3'h7 ? _GEN_1122 : valid_64; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1637 = state == 3'h7 ? _GEN_1123 : valid_65; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1638 = state == 3'h7 ? _GEN_1124 : valid_66; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1639 = state == 3'h7 ? _GEN_1125 : valid_67; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1640 = state == 3'h7 ? _GEN_1126 : valid_68; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1641 = state == 3'h7 ? _GEN_1127 : valid_69; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1642 = state == 3'h7 ? _GEN_1128 : valid_70; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1643 = state == 3'h7 ? _GEN_1129 : valid_71; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1644 = state == 3'h7 ? _GEN_1130 : valid_72; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1645 = state == 3'h7 ? _GEN_1131 : valid_73; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1646 = state == 3'h7 ? _GEN_1132 : valid_74; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1647 = state == 3'h7 ? _GEN_1133 : valid_75; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1648 = state == 3'h7 ? _GEN_1134 : valid_76; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1649 = state == 3'h7 ? _GEN_1135 : valid_77; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1650 = state == 3'h7 ? _GEN_1136 : valid_78; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1651 = state == 3'h7 ? _GEN_1137 : valid_79; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1652 = state == 3'h7 ? _GEN_1138 : valid_80; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1653 = state == 3'h7 ? _GEN_1139 : valid_81; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1654 = state == 3'h7 ? _GEN_1140 : valid_82; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1655 = state == 3'h7 ? _GEN_1141 : valid_83; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1656 = state == 3'h7 ? _GEN_1142 : valid_84; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1657 = state == 3'h7 ? _GEN_1143 : valid_85; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1658 = state == 3'h7 ? _GEN_1144 : valid_86; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1659 = state == 3'h7 ? _GEN_1145 : valid_87; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1660 = state == 3'h7 ? _GEN_1146 : valid_88; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1661 = state == 3'h7 ? _GEN_1147 : valid_89; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1662 = state == 3'h7 ? _GEN_1148 : valid_90; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1663 = state == 3'h7 ? _GEN_1149 : valid_91; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1664 = state == 3'h7 ? _GEN_1150 : valid_92; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1665 = state == 3'h7 ? _GEN_1151 : valid_93; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1666 = state == 3'h7 ? _GEN_1152 : valid_94; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1667 = state == 3'h7 ? _GEN_1153 : valid_95; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1668 = state == 3'h7 ? _GEN_1154 : valid_96; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1669 = state == 3'h7 ? _GEN_1155 : valid_97; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1670 = state == 3'h7 ? _GEN_1156 : valid_98; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1671 = state == 3'h7 ? _GEN_1157 : valid_99; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1672 = state == 3'h7 ? _GEN_1158 : valid_100; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1673 = state == 3'h7 ? _GEN_1159 : valid_101; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1674 = state == 3'h7 ? _GEN_1160 : valid_102; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1675 = state == 3'h7 ? _GEN_1161 : valid_103; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1676 = state == 3'h7 ? _GEN_1162 : valid_104; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1677 = state == 3'h7 ? _GEN_1163 : valid_105; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1678 = state == 3'h7 ? _GEN_1164 : valid_106; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1679 = state == 3'h7 ? _GEN_1165 : valid_107; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1680 = state == 3'h7 ? _GEN_1166 : valid_108; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1681 = state == 3'h7 ? _GEN_1167 : valid_109; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1682 = state == 3'h7 ? _GEN_1168 : valid_110; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1683 = state == 3'h7 ? _GEN_1169 : valid_111; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1684 = state == 3'h7 ? _GEN_1170 : valid_112; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1685 = state == 3'h7 ? _GEN_1171 : valid_113; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1686 = state == 3'h7 ? _GEN_1172 : valid_114; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1687 = state == 3'h7 ? _GEN_1173 : valid_115; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1688 = state == 3'h7 ? _GEN_1174 : valid_116; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1689 = state == 3'h7 ? _GEN_1175 : valid_117; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1690 = state == 3'h7 ? _GEN_1176 : valid_118; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1691 = state == 3'h7 ? _GEN_1177 : valid_119; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1692 = state == 3'h7 ? _GEN_1178 : valid_120; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1693 = state == 3'h7 ? _GEN_1179 : valid_121; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1694 = state == 3'h7 ? _GEN_1180 : valid_122; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1695 = state == 3'h7 ? _GEN_1181 : valid_123; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1696 = state == 3'h7 ? _GEN_1182 : valid_124; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1697 = state == 3'h7 ? _GEN_1183 : valid_125; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1698 = state == 3'h7 ? _GEN_1184 : valid_126; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1699 = state == 3'h7 ? _GEN_1185 : valid_127; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1700 = state == 3'h7 ? _GEN_1186 : valid_128; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1701 = state == 3'h7 ? _GEN_1187 : valid_129; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1702 = state == 3'h7 ? _GEN_1188 : valid_130; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1703 = state == 3'h7 ? _GEN_1189 : valid_131; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1704 = state == 3'h7 ? _GEN_1190 : valid_132; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1705 = state == 3'h7 ? _GEN_1191 : valid_133; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1706 = state == 3'h7 ? _GEN_1192 : valid_134; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1707 = state == 3'h7 ? _GEN_1193 : valid_135; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1708 = state == 3'h7 ? _GEN_1194 : valid_136; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1709 = state == 3'h7 ? _GEN_1195 : valid_137; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1710 = state == 3'h7 ? _GEN_1196 : valid_138; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1711 = state == 3'h7 ? _GEN_1197 : valid_139; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1712 = state == 3'h7 ? _GEN_1198 : valid_140; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1713 = state == 3'h7 ? _GEN_1199 : valid_141; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1714 = state == 3'h7 ? _GEN_1200 : valid_142; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1715 = state == 3'h7 ? _GEN_1201 : valid_143; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1716 = state == 3'h7 ? _GEN_1202 : valid_144; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1717 = state == 3'h7 ? _GEN_1203 : valid_145; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1718 = state == 3'h7 ? _GEN_1204 : valid_146; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1719 = state == 3'h7 ? _GEN_1205 : valid_147; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1720 = state == 3'h7 ? _GEN_1206 : valid_148; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1721 = state == 3'h7 ? _GEN_1207 : valid_149; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1722 = state == 3'h7 ? _GEN_1208 : valid_150; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1723 = state == 3'h7 ? _GEN_1209 : valid_151; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1724 = state == 3'h7 ? _GEN_1210 : valid_152; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1725 = state == 3'h7 ? _GEN_1211 : valid_153; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1726 = state == 3'h7 ? _GEN_1212 : valid_154; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1727 = state == 3'h7 ? _GEN_1213 : valid_155; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1728 = state == 3'h7 ? _GEN_1214 : valid_156; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1729 = state == 3'h7 ? _GEN_1215 : valid_157; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1730 = state == 3'h7 ? _GEN_1216 : valid_158; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1731 = state == 3'h7 ? _GEN_1217 : valid_159; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1732 = state == 3'h7 ? _GEN_1218 : valid_160; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1733 = state == 3'h7 ? _GEN_1219 : valid_161; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1734 = state == 3'h7 ? _GEN_1220 : valid_162; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1735 = state == 3'h7 ? _GEN_1221 : valid_163; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1736 = state == 3'h7 ? _GEN_1222 : valid_164; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1737 = state == 3'h7 ? _GEN_1223 : valid_165; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1738 = state == 3'h7 ? _GEN_1224 : valid_166; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1739 = state == 3'h7 ? _GEN_1225 : valid_167; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1740 = state == 3'h7 ? _GEN_1226 : valid_168; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1741 = state == 3'h7 ? _GEN_1227 : valid_169; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1742 = state == 3'h7 ? _GEN_1228 : valid_170; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1743 = state == 3'h7 ? _GEN_1229 : valid_171; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1744 = state == 3'h7 ? _GEN_1230 : valid_172; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1745 = state == 3'h7 ? _GEN_1231 : valid_173; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1746 = state == 3'h7 ? _GEN_1232 : valid_174; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1747 = state == 3'h7 ? _GEN_1233 : valid_175; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1748 = state == 3'h7 ? _GEN_1234 : valid_176; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1749 = state == 3'h7 ? _GEN_1235 : valid_177; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1750 = state == 3'h7 ? _GEN_1236 : valid_178; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1751 = state == 3'h7 ? _GEN_1237 : valid_179; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1752 = state == 3'h7 ? _GEN_1238 : valid_180; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1753 = state == 3'h7 ? _GEN_1239 : valid_181; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1754 = state == 3'h7 ? _GEN_1240 : valid_182; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1755 = state == 3'h7 ? _GEN_1241 : valid_183; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1756 = state == 3'h7 ? _GEN_1242 : valid_184; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1757 = state == 3'h7 ? _GEN_1243 : valid_185; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1758 = state == 3'h7 ? _GEN_1244 : valid_186; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1759 = state == 3'h7 ? _GEN_1245 : valid_187; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1760 = state == 3'h7 ? _GEN_1246 : valid_188; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1761 = state == 3'h7 ? _GEN_1247 : valid_189; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1762 = state == 3'h7 ? _GEN_1248 : valid_190; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1763 = state == 3'h7 ? _GEN_1249 : valid_191; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1764 = state == 3'h7 ? _GEN_1250 : valid_192; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1765 = state == 3'h7 ? _GEN_1251 : valid_193; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1766 = state == 3'h7 ? _GEN_1252 : valid_194; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1767 = state == 3'h7 ? _GEN_1253 : valid_195; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1768 = state == 3'h7 ? _GEN_1254 : valid_196; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1769 = state == 3'h7 ? _GEN_1255 : valid_197; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1770 = state == 3'h7 ? _GEN_1256 : valid_198; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1771 = state == 3'h7 ? _GEN_1257 : valid_199; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1772 = state == 3'h7 ? _GEN_1258 : valid_200; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1773 = state == 3'h7 ? _GEN_1259 : valid_201; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1774 = state == 3'h7 ? _GEN_1260 : valid_202; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1775 = state == 3'h7 ? _GEN_1261 : valid_203; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1776 = state == 3'h7 ? _GEN_1262 : valid_204; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1777 = state == 3'h7 ? _GEN_1263 : valid_205; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1778 = state == 3'h7 ? _GEN_1264 : valid_206; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1779 = state == 3'h7 ? _GEN_1265 : valid_207; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1780 = state == 3'h7 ? _GEN_1266 : valid_208; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1781 = state == 3'h7 ? _GEN_1267 : valid_209; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1782 = state == 3'h7 ? _GEN_1268 : valid_210; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1783 = state == 3'h7 ? _GEN_1269 : valid_211; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1784 = state == 3'h7 ? _GEN_1270 : valid_212; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1785 = state == 3'h7 ? _GEN_1271 : valid_213; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1786 = state == 3'h7 ? _GEN_1272 : valid_214; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1787 = state == 3'h7 ? _GEN_1273 : valid_215; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1788 = state == 3'h7 ? _GEN_1274 : valid_216; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1789 = state == 3'h7 ? _GEN_1275 : valid_217; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1790 = state == 3'h7 ? _GEN_1276 : valid_218; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1791 = state == 3'h7 ? _GEN_1277 : valid_219; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1792 = state == 3'h7 ? _GEN_1278 : valid_220; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1793 = state == 3'h7 ? _GEN_1279 : valid_221; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1794 = state == 3'h7 ? _GEN_1280 : valid_222; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1795 = state == 3'h7 ? _GEN_1281 : valid_223; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1796 = state == 3'h7 ? _GEN_1282 : valid_224; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1797 = state == 3'h7 ? _GEN_1283 : valid_225; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1798 = state == 3'h7 ? _GEN_1284 : valid_226; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1799 = state == 3'h7 ? _GEN_1285 : valid_227; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1800 = state == 3'h7 ? _GEN_1286 : valid_228; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1801 = state == 3'h7 ? _GEN_1287 : valid_229; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1802 = state == 3'h7 ? _GEN_1288 : valid_230; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1803 = state == 3'h7 ? _GEN_1289 : valid_231; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1804 = state == 3'h7 ? _GEN_1290 : valid_232; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1805 = state == 3'h7 ? _GEN_1291 : valid_233; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1806 = state == 3'h7 ? _GEN_1292 : valid_234; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1807 = state == 3'h7 ? _GEN_1293 : valid_235; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1808 = state == 3'h7 ? _GEN_1294 : valid_236; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1809 = state == 3'h7 ? _GEN_1295 : valid_237; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1810 = state == 3'h7 ? _GEN_1296 : valid_238; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1811 = state == 3'h7 ? _GEN_1297 : valid_239; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1812 = state == 3'h7 ? _GEN_1298 : valid_240; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1813 = state == 3'h7 ? _GEN_1299 : valid_241; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1814 = state == 3'h7 ? _GEN_1300 : valid_242; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1815 = state == 3'h7 ? _GEN_1301 : valid_243; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1816 = state == 3'h7 ? _GEN_1302 : valid_244; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1817 = state == 3'h7 ? _GEN_1303 : valid_245; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1818 = state == 3'h7 ? _GEN_1304 : valid_246; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1819 = state == 3'h7 ? _GEN_1305 : valid_247; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1820 = state == 3'h7 ? _GEN_1306 : valid_248; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1821 = state == 3'h7 ? _GEN_1307 : valid_249; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1822 = state == 3'h7 ? _GEN_1308 : valid_250; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1823 = state == 3'h7 ? _GEN_1309 : valid_251; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1824 = state == 3'h7 ? _GEN_1310 : valid_252; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1825 = state == 3'h7 ? _GEN_1311 : valid_253; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1826 = state == 3'h7 ? _GEN_1312 : valid_254; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1827 = state == 3'h7 ? _GEN_1313 : valid_255; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1828 = state == 3'h7 ? _GEN_1314 : valid_256; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1829 = state == 3'h7 ? _GEN_1315 : valid_257; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1830 = state == 3'h7 ? _GEN_1316 : valid_258; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1831 = state == 3'h7 ? _GEN_1317 : valid_259; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1832 = state == 3'h7 ? _GEN_1318 : valid_260; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1833 = state == 3'h7 ? _GEN_1319 : valid_261; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1834 = state == 3'h7 ? _GEN_1320 : valid_262; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1835 = state == 3'h7 ? _GEN_1321 : valid_263; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1836 = state == 3'h7 ? _GEN_1322 : valid_264; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1837 = state == 3'h7 ? _GEN_1323 : valid_265; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1838 = state == 3'h7 ? _GEN_1324 : valid_266; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1839 = state == 3'h7 ? _GEN_1325 : valid_267; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1840 = state == 3'h7 ? _GEN_1326 : valid_268; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1841 = state == 3'h7 ? _GEN_1327 : valid_269; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1842 = state == 3'h7 ? _GEN_1328 : valid_270; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1843 = state == 3'h7 ? _GEN_1329 : valid_271; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1844 = state == 3'h7 ? _GEN_1330 : valid_272; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1845 = state == 3'h7 ? _GEN_1331 : valid_273; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1846 = state == 3'h7 ? _GEN_1332 : valid_274; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1847 = state == 3'h7 ? _GEN_1333 : valid_275; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1848 = state == 3'h7 ? _GEN_1334 : valid_276; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1849 = state == 3'h7 ? _GEN_1335 : valid_277; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1850 = state == 3'h7 ? _GEN_1336 : valid_278; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1851 = state == 3'h7 ? _GEN_1337 : valid_279; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1852 = state == 3'h7 ? _GEN_1338 : valid_280; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1853 = state == 3'h7 ? _GEN_1339 : valid_281; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1854 = state == 3'h7 ? _GEN_1340 : valid_282; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1855 = state == 3'h7 ? _GEN_1341 : valid_283; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1856 = state == 3'h7 ? _GEN_1342 : valid_284; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1857 = state == 3'h7 ? _GEN_1343 : valid_285; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1858 = state == 3'h7 ? _GEN_1344 : valid_286; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1859 = state == 3'h7 ? _GEN_1345 : valid_287; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1860 = state == 3'h7 ? _GEN_1346 : valid_288; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1861 = state == 3'h7 ? _GEN_1347 : valid_289; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1862 = state == 3'h7 ? _GEN_1348 : valid_290; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1863 = state == 3'h7 ? _GEN_1349 : valid_291; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1864 = state == 3'h7 ? _GEN_1350 : valid_292; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1865 = state == 3'h7 ? _GEN_1351 : valid_293; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1866 = state == 3'h7 ? _GEN_1352 : valid_294; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1867 = state == 3'h7 ? _GEN_1353 : valid_295; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1868 = state == 3'h7 ? _GEN_1354 : valid_296; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1869 = state == 3'h7 ? _GEN_1355 : valid_297; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1870 = state == 3'h7 ? _GEN_1356 : valid_298; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1871 = state == 3'h7 ? _GEN_1357 : valid_299; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1872 = state == 3'h7 ? _GEN_1358 : valid_300; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1873 = state == 3'h7 ? _GEN_1359 : valid_301; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1874 = state == 3'h7 ? _GEN_1360 : valid_302; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1875 = state == 3'h7 ? _GEN_1361 : valid_303; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1876 = state == 3'h7 ? _GEN_1362 : valid_304; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1877 = state == 3'h7 ? _GEN_1363 : valid_305; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1878 = state == 3'h7 ? _GEN_1364 : valid_306; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1879 = state == 3'h7 ? _GEN_1365 : valid_307; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1880 = state == 3'h7 ? _GEN_1366 : valid_308; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1881 = state == 3'h7 ? _GEN_1367 : valid_309; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1882 = state == 3'h7 ? _GEN_1368 : valid_310; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1883 = state == 3'h7 ? _GEN_1369 : valid_311; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1884 = state == 3'h7 ? _GEN_1370 : valid_312; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1885 = state == 3'h7 ? _GEN_1371 : valid_313; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1886 = state == 3'h7 ? _GEN_1372 : valid_314; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1887 = state == 3'h7 ? _GEN_1373 : valid_315; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1888 = state == 3'h7 ? _GEN_1374 : valid_316; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1889 = state == 3'h7 ? _GEN_1375 : valid_317; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1890 = state == 3'h7 ? _GEN_1376 : valid_318; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1891 = state == 3'h7 ? _GEN_1377 : valid_319; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1892 = state == 3'h7 ? _GEN_1378 : valid_320; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1893 = state == 3'h7 ? _GEN_1379 : valid_321; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1894 = state == 3'h7 ? _GEN_1380 : valid_322; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1895 = state == 3'h7 ? _GEN_1381 : valid_323; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1896 = state == 3'h7 ? _GEN_1382 : valid_324; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1897 = state == 3'h7 ? _GEN_1383 : valid_325; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1898 = state == 3'h7 ? _GEN_1384 : valid_326; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1899 = state == 3'h7 ? _GEN_1385 : valid_327; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1900 = state == 3'h7 ? _GEN_1386 : valid_328; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1901 = state == 3'h7 ? _GEN_1387 : valid_329; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1902 = state == 3'h7 ? _GEN_1388 : valid_330; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1903 = state == 3'h7 ? _GEN_1389 : valid_331; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1904 = state == 3'h7 ? _GEN_1390 : valid_332; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1905 = state == 3'h7 ? _GEN_1391 : valid_333; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1906 = state == 3'h7 ? _GEN_1392 : valid_334; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1907 = state == 3'h7 ? _GEN_1393 : valid_335; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1908 = state == 3'h7 ? _GEN_1394 : valid_336; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1909 = state == 3'h7 ? _GEN_1395 : valid_337; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1910 = state == 3'h7 ? _GEN_1396 : valid_338; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1911 = state == 3'h7 ? _GEN_1397 : valid_339; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1912 = state == 3'h7 ? _GEN_1398 : valid_340; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1913 = state == 3'h7 ? _GEN_1399 : valid_341; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1914 = state == 3'h7 ? _GEN_1400 : valid_342; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1915 = state == 3'h7 ? _GEN_1401 : valid_343; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1916 = state == 3'h7 ? _GEN_1402 : valid_344; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1917 = state == 3'h7 ? _GEN_1403 : valid_345; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1918 = state == 3'h7 ? _GEN_1404 : valid_346; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1919 = state == 3'h7 ? _GEN_1405 : valid_347; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1920 = state == 3'h7 ? _GEN_1406 : valid_348; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1921 = state == 3'h7 ? _GEN_1407 : valid_349; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1922 = state == 3'h7 ? _GEN_1408 : valid_350; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1923 = state == 3'h7 ? _GEN_1409 : valid_351; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1924 = state == 3'h7 ? _GEN_1410 : valid_352; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1925 = state == 3'h7 ? _GEN_1411 : valid_353; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1926 = state == 3'h7 ? _GEN_1412 : valid_354; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1927 = state == 3'h7 ? _GEN_1413 : valid_355; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1928 = state == 3'h7 ? _GEN_1414 : valid_356; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1929 = state == 3'h7 ? _GEN_1415 : valid_357; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1930 = state == 3'h7 ? _GEN_1416 : valid_358; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1931 = state == 3'h7 ? _GEN_1417 : valid_359; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1932 = state == 3'h7 ? _GEN_1418 : valid_360; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1933 = state == 3'h7 ? _GEN_1419 : valid_361; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1934 = state == 3'h7 ? _GEN_1420 : valid_362; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1935 = state == 3'h7 ? _GEN_1421 : valid_363; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1936 = state == 3'h7 ? _GEN_1422 : valid_364; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1937 = state == 3'h7 ? _GEN_1423 : valid_365; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1938 = state == 3'h7 ? _GEN_1424 : valid_366; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1939 = state == 3'h7 ? _GEN_1425 : valid_367; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1940 = state == 3'h7 ? _GEN_1426 : valid_368; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1941 = state == 3'h7 ? _GEN_1427 : valid_369; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1942 = state == 3'h7 ? _GEN_1428 : valid_370; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1943 = state == 3'h7 ? _GEN_1429 : valid_371; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1944 = state == 3'h7 ? _GEN_1430 : valid_372; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1945 = state == 3'h7 ? _GEN_1431 : valid_373; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1946 = state == 3'h7 ? _GEN_1432 : valid_374; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1947 = state == 3'h7 ? _GEN_1433 : valid_375; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1948 = state == 3'h7 ? _GEN_1434 : valid_376; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1949 = state == 3'h7 ? _GEN_1435 : valid_377; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1950 = state == 3'h7 ? _GEN_1436 : valid_378; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1951 = state == 3'h7 ? _GEN_1437 : valid_379; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1952 = state == 3'h7 ? _GEN_1438 : valid_380; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1953 = state == 3'h7 ? _GEN_1439 : valid_381; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1954 = state == 3'h7 ? _GEN_1440 : valid_382; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1955 = state == 3'h7 ? _GEN_1441 : valid_383; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1956 = state == 3'h7 ? _GEN_1442 : valid_384; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1957 = state == 3'h7 ? _GEN_1443 : valid_385; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1958 = state == 3'h7 ? _GEN_1444 : valid_386; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1959 = state == 3'h7 ? _GEN_1445 : valid_387; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1960 = state == 3'h7 ? _GEN_1446 : valid_388; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1961 = state == 3'h7 ? _GEN_1447 : valid_389; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1962 = state == 3'h7 ? _GEN_1448 : valid_390; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1963 = state == 3'h7 ? _GEN_1449 : valid_391; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1964 = state == 3'h7 ? _GEN_1450 : valid_392; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1965 = state == 3'h7 ? _GEN_1451 : valid_393; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1966 = state == 3'h7 ? _GEN_1452 : valid_394; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1967 = state == 3'h7 ? _GEN_1453 : valid_395; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1968 = state == 3'h7 ? _GEN_1454 : valid_396; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1969 = state == 3'h7 ? _GEN_1455 : valid_397; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1970 = state == 3'h7 ? _GEN_1456 : valid_398; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1971 = state == 3'h7 ? _GEN_1457 : valid_399; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1972 = state == 3'h7 ? _GEN_1458 : valid_400; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1973 = state == 3'h7 ? _GEN_1459 : valid_401; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1974 = state == 3'h7 ? _GEN_1460 : valid_402; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1975 = state == 3'h7 ? _GEN_1461 : valid_403; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1976 = state == 3'h7 ? _GEN_1462 : valid_404; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1977 = state == 3'h7 ? _GEN_1463 : valid_405; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1978 = state == 3'h7 ? _GEN_1464 : valid_406; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1979 = state == 3'h7 ? _GEN_1465 : valid_407; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1980 = state == 3'h7 ? _GEN_1466 : valid_408; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1981 = state == 3'h7 ? _GEN_1467 : valid_409; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1982 = state == 3'h7 ? _GEN_1468 : valid_410; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1983 = state == 3'h7 ? _GEN_1469 : valid_411; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1984 = state == 3'h7 ? _GEN_1470 : valid_412; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1985 = state == 3'h7 ? _GEN_1471 : valid_413; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1986 = state == 3'h7 ? _GEN_1472 : valid_414; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1987 = state == 3'h7 ? _GEN_1473 : valid_415; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1988 = state == 3'h7 ? _GEN_1474 : valid_416; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1989 = state == 3'h7 ? _GEN_1475 : valid_417; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1990 = state == 3'h7 ? _GEN_1476 : valid_418; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1991 = state == 3'h7 ? _GEN_1477 : valid_419; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1992 = state == 3'h7 ? _GEN_1478 : valid_420; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1993 = state == 3'h7 ? _GEN_1479 : valid_421; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1994 = state == 3'h7 ? _GEN_1480 : valid_422; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1995 = state == 3'h7 ? _GEN_1481 : valid_423; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1996 = state == 3'h7 ? _GEN_1482 : valid_424; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1997 = state == 3'h7 ? _GEN_1483 : valid_425; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1998 = state == 3'h7 ? _GEN_1484 : valid_426; // @[DCache.scala 165:26 56:22]
  wire  _GEN_1999 = state == 3'h7 ? _GEN_1485 : valid_427; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2000 = state == 3'h7 ? _GEN_1486 : valid_428; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2001 = state == 3'h7 ? _GEN_1487 : valid_429; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2002 = state == 3'h7 ? _GEN_1488 : valid_430; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2003 = state == 3'h7 ? _GEN_1489 : valid_431; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2004 = state == 3'h7 ? _GEN_1490 : valid_432; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2005 = state == 3'h7 ? _GEN_1491 : valid_433; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2006 = state == 3'h7 ? _GEN_1492 : valid_434; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2007 = state == 3'h7 ? _GEN_1493 : valid_435; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2008 = state == 3'h7 ? _GEN_1494 : valid_436; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2009 = state == 3'h7 ? _GEN_1495 : valid_437; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2010 = state == 3'h7 ? _GEN_1496 : valid_438; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2011 = state == 3'h7 ? _GEN_1497 : valid_439; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2012 = state == 3'h7 ? _GEN_1498 : valid_440; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2013 = state == 3'h7 ? _GEN_1499 : valid_441; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2014 = state == 3'h7 ? _GEN_1500 : valid_442; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2015 = state == 3'h7 ? _GEN_1501 : valid_443; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2016 = state == 3'h7 ? _GEN_1502 : valid_444; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2017 = state == 3'h7 ? _GEN_1503 : valid_445; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2018 = state == 3'h7 ? _GEN_1504 : valid_446; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2019 = state == 3'h7 ? _GEN_1505 : valid_447; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2020 = state == 3'h7 ? _GEN_1506 : valid_448; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2021 = state == 3'h7 ? _GEN_1507 : valid_449; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2022 = state == 3'h7 ? _GEN_1508 : valid_450; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2023 = state == 3'h7 ? _GEN_1509 : valid_451; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2024 = state == 3'h7 ? _GEN_1510 : valid_452; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2025 = state == 3'h7 ? _GEN_1511 : valid_453; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2026 = state == 3'h7 ? _GEN_1512 : valid_454; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2027 = state == 3'h7 ? _GEN_1513 : valid_455; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2028 = state == 3'h7 ? _GEN_1514 : valid_456; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2029 = state == 3'h7 ? _GEN_1515 : valid_457; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2030 = state == 3'h7 ? _GEN_1516 : valid_458; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2031 = state == 3'h7 ? _GEN_1517 : valid_459; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2032 = state == 3'h7 ? _GEN_1518 : valid_460; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2033 = state == 3'h7 ? _GEN_1519 : valid_461; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2034 = state == 3'h7 ? _GEN_1520 : valid_462; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2035 = state == 3'h7 ? _GEN_1521 : valid_463; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2036 = state == 3'h7 ? _GEN_1522 : valid_464; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2037 = state == 3'h7 ? _GEN_1523 : valid_465; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2038 = state == 3'h7 ? _GEN_1524 : valid_466; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2039 = state == 3'h7 ? _GEN_1525 : valid_467; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2040 = state == 3'h7 ? _GEN_1526 : valid_468; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2041 = state == 3'h7 ? _GEN_1527 : valid_469; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2042 = state == 3'h7 ? _GEN_1528 : valid_470; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2043 = state == 3'h7 ? _GEN_1529 : valid_471; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2044 = state == 3'h7 ? _GEN_1530 : valid_472; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2045 = state == 3'h7 ? _GEN_1531 : valid_473; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2046 = state == 3'h7 ? _GEN_1532 : valid_474; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2047 = state == 3'h7 ? _GEN_1533 : valid_475; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2048 = state == 3'h7 ? _GEN_1534 : valid_476; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2049 = state == 3'h7 ? _GEN_1535 : valid_477; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2050 = state == 3'h7 ? _GEN_1536 : valid_478; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2051 = state == 3'h7 ? _GEN_1537 : valid_479; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2052 = state == 3'h7 ? _GEN_1538 : valid_480; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2053 = state == 3'h7 ? _GEN_1539 : valid_481; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2054 = state == 3'h7 ? _GEN_1540 : valid_482; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2055 = state == 3'h7 ? _GEN_1541 : valid_483; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2056 = state == 3'h7 ? _GEN_1542 : valid_484; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2057 = state == 3'h7 ? _GEN_1543 : valid_485; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2058 = state == 3'h7 ? _GEN_1544 : valid_486; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2059 = state == 3'h7 ? _GEN_1545 : valid_487; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2060 = state == 3'h7 ? _GEN_1546 : valid_488; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2061 = state == 3'h7 ? _GEN_1547 : valid_489; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2062 = state == 3'h7 ? _GEN_1548 : valid_490; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2063 = state == 3'h7 ? _GEN_1549 : valid_491; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2064 = state == 3'h7 ? _GEN_1550 : valid_492; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2065 = state == 3'h7 ? _GEN_1551 : valid_493; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2066 = state == 3'h7 ? _GEN_1552 : valid_494; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2067 = state == 3'h7 ? _GEN_1553 : valid_495; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2068 = state == 3'h7 ? _GEN_1554 : valid_496; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2069 = state == 3'h7 ? _GEN_1555 : valid_497; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2070 = state == 3'h7 ? _GEN_1556 : valid_498; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2071 = state == 3'h7 ? _GEN_1557 : valid_499; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2072 = state == 3'h7 ? _GEN_1558 : valid_500; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2073 = state == 3'h7 ? _GEN_1559 : valid_501; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2074 = state == 3'h7 ? _GEN_1560 : valid_502; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2075 = state == 3'h7 ? _GEN_1561 : valid_503; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2076 = state == 3'h7 ? _GEN_1562 : valid_504; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2077 = state == 3'h7 ? _GEN_1563 : valid_505; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2078 = state == 3'h7 ? _GEN_1564 : valid_506; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2079 = state == 3'h7 ? _GEN_1565 : valid_507; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2080 = state == 3'h7 ? _GEN_1566 : valid_508; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2081 = state == 3'h7 ? _GEN_1567 : valid_509; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2082 = state == 3'h7 ? _GEN_1568 : valid_510; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2083 = state == 3'h7 ? _GEN_1569 : valid_511; // @[DCache.scala 165:26 56:22]
  wire  _GEN_2086 = _array_io_en_T_1 ? _GEN_1572 : valid_0; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2087 = _array_io_en_T_1 ? _GEN_1573 : valid_1; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2088 = _array_io_en_T_1 ? _GEN_1574 : valid_2; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2089 = _array_io_en_T_1 ? _GEN_1575 : valid_3; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2090 = _array_io_en_T_1 ? _GEN_1576 : valid_4; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2091 = _array_io_en_T_1 ? _GEN_1577 : valid_5; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2092 = _array_io_en_T_1 ? _GEN_1578 : valid_6; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2093 = _array_io_en_T_1 ? _GEN_1579 : valid_7; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2094 = _array_io_en_T_1 ? _GEN_1580 : valid_8; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2095 = _array_io_en_T_1 ? _GEN_1581 : valid_9; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2096 = _array_io_en_T_1 ? _GEN_1582 : valid_10; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2097 = _array_io_en_T_1 ? _GEN_1583 : valid_11; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2098 = _array_io_en_T_1 ? _GEN_1584 : valid_12; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2099 = _array_io_en_T_1 ? _GEN_1585 : valid_13; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2100 = _array_io_en_T_1 ? _GEN_1586 : valid_14; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2101 = _array_io_en_T_1 ? _GEN_1587 : valid_15; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2102 = _array_io_en_T_1 ? _GEN_1588 : valid_16; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2103 = _array_io_en_T_1 ? _GEN_1589 : valid_17; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2104 = _array_io_en_T_1 ? _GEN_1590 : valid_18; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2105 = _array_io_en_T_1 ? _GEN_1591 : valid_19; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2106 = _array_io_en_T_1 ? _GEN_1592 : valid_20; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2107 = _array_io_en_T_1 ? _GEN_1593 : valid_21; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2108 = _array_io_en_T_1 ? _GEN_1594 : valid_22; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2109 = _array_io_en_T_1 ? _GEN_1595 : valid_23; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2110 = _array_io_en_T_1 ? _GEN_1596 : valid_24; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2111 = _array_io_en_T_1 ? _GEN_1597 : valid_25; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2112 = _array_io_en_T_1 ? _GEN_1598 : valid_26; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2113 = _array_io_en_T_1 ? _GEN_1599 : valid_27; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2114 = _array_io_en_T_1 ? _GEN_1600 : valid_28; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2115 = _array_io_en_T_1 ? _GEN_1601 : valid_29; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2116 = _array_io_en_T_1 ? _GEN_1602 : valid_30; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2117 = _array_io_en_T_1 ? _GEN_1603 : valid_31; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2118 = _array_io_en_T_1 ? _GEN_1604 : valid_32; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2119 = _array_io_en_T_1 ? _GEN_1605 : valid_33; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2120 = _array_io_en_T_1 ? _GEN_1606 : valid_34; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2121 = _array_io_en_T_1 ? _GEN_1607 : valid_35; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2122 = _array_io_en_T_1 ? _GEN_1608 : valid_36; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2123 = _array_io_en_T_1 ? _GEN_1609 : valid_37; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2124 = _array_io_en_T_1 ? _GEN_1610 : valid_38; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2125 = _array_io_en_T_1 ? _GEN_1611 : valid_39; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2126 = _array_io_en_T_1 ? _GEN_1612 : valid_40; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2127 = _array_io_en_T_1 ? _GEN_1613 : valid_41; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2128 = _array_io_en_T_1 ? _GEN_1614 : valid_42; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2129 = _array_io_en_T_1 ? _GEN_1615 : valid_43; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2130 = _array_io_en_T_1 ? _GEN_1616 : valid_44; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2131 = _array_io_en_T_1 ? _GEN_1617 : valid_45; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2132 = _array_io_en_T_1 ? _GEN_1618 : valid_46; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2133 = _array_io_en_T_1 ? _GEN_1619 : valid_47; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2134 = _array_io_en_T_1 ? _GEN_1620 : valid_48; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2135 = _array_io_en_T_1 ? _GEN_1621 : valid_49; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2136 = _array_io_en_T_1 ? _GEN_1622 : valid_50; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2137 = _array_io_en_T_1 ? _GEN_1623 : valid_51; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2138 = _array_io_en_T_1 ? _GEN_1624 : valid_52; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2139 = _array_io_en_T_1 ? _GEN_1625 : valid_53; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2140 = _array_io_en_T_1 ? _GEN_1626 : valid_54; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2141 = _array_io_en_T_1 ? _GEN_1627 : valid_55; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2142 = _array_io_en_T_1 ? _GEN_1628 : valid_56; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2143 = _array_io_en_T_1 ? _GEN_1629 : valid_57; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2144 = _array_io_en_T_1 ? _GEN_1630 : valid_58; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2145 = _array_io_en_T_1 ? _GEN_1631 : valid_59; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2146 = _array_io_en_T_1 ? _GEN_1632 : valid_60; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2147 = _array_io_en_T_1 ? _GEN_1633 : valid_61; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2148 = _array_io_en_T_1 ? _GEN_1634 : valid_62; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2149 = _array_io_en_T_1 ? _GEN_1635 : valid_63; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2150 = _array_io_en_T_1 ? _GEN_1636 : valid_64; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2151 = _array_io_en_T_1 ? _GEN_1637 : valid_65; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2152 = _array_io_en_T_1 ? _GEN_1638 : valid_66; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2153 = _array_io_en_T_1 ? _GEN_1639 : valid_67; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2154 = _array_io_en_T_1 ? _GEN_1640 : valid_68; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2155 = _array_io_en_T_1 ? _GEN_1641 : valid_69; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2156 = _array_io_en_T_1 ? _GEN_1642 : valid_70; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2157 = _array_io_en_T_1 ? _GEN_1643 : valid_71; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2158 = _array_io_en_T_1 ? _GEN_1644 : valid_72; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2159 = _array_io_en_T_1 ? _GEN_1645 : valid_73; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2160 = _array_io_en_T_1 ? _GEN_1646 : valid_74; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2161 = _array_io_en_T_1 ? _GEN_1647 : valid_75; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2162 = _array_io_en_T_1 ? _GEN_1648 : valid_76; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2163 = _array_io_en_T_1 ? _GEN_1649 : valid_77; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2164 = _array_io_en_T_1 ? _GEN_1650 : valid_78; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2165 = _array_io_en_T_1 ? _GEN_1651 : valid_79; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2166 = _array_io_en_T_1 ? _GEN_1652 : valid_80; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2167 = _array_io_en_T_1 ? _GEN_1653 : valid_81; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2168 = _array_io_en_T_1 ? _GEN_1654 : valid_82; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2169 = _array_io_en_T_1 ? _GEN_1655 : valid_83; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2170 = _array_io_en_T_1 ? _GEN_1656 : valid_84; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2171 = _array_io_en_T_1 ? _GEN_1657 : valid_85; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2172 = _array_io_en_T_1 ? _GEN_1658 : valid_86; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2173 = _array_io_en_T_1 ? _GEN_1659 : valid_87; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2174 = _array_io_en_T_1 ? _GEN_1660 : valid_88; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2175 = _array_io_en_T_1 ? _GEN_1661 : valid_89; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2176 = _array_io_en_T_1 ? _GEN_1662 : valid_90; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2177 = _array_io_en_T_1 ? _GEN_1663 : valid_91; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2178 = _array_io_en_T_1 ? _GEN_1664 : valid_92; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2179 = _array_io_en_T_1 ? _GEN_1665 : valid_93; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2180 = _array_io_en_T_1 ? _GEN_1666 : valid_94; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2181 = _array_io_en_T_1 ? _GEN_1667 : valid_95; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2182 = _array_io_en_T_1 ? _GEN_1668 : valid_96; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2183 = _array_io_en_T_1 ? _GEN_1669 : valid_97; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2184 = _array_io_en_T_1 ? _GEN_1670 : valid_98; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2185 = _array_io_en_T_1 ? _GEN_1671 : valid_99; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2186 = _array_io_en_T_1 ? _GEN_1672 : valid_100; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2187 = _array_io_en_T_1 ? _GEN_1673 : valid_101; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2188 = _array_io_en_T_1 ? _GEN_1674 : valid_102; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2189 = _array_io_en_T_1 ? _GEN_1675 : valid_103; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2190 = _array_io_en_T_1 ? _GEN_1676 : valid_104; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2191 = _array_io_en_T_1 ? _GEN_1677 : valid_105; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2192 = _array_io_en_T_1 ? _GEN_1678 : valid_106; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2193 = _array_io_en_T_1 ? _GEN_1679 : valid_107; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2194 = _array_io_en_T_1 ? _GEN_1680 : valid_108; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2195 = _array_io_en_T_1 ? _GEN_1681 : valid_109; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2196 = _array_io_en_T_1 ? _GEN_1682 : valid_110; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2197 = _array_io_en_T_1 ? _GEN_1683 : valid_111; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2198 = _array_io_en_T_1 ? _GEN_1684 : valid_112; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2199 = _array_io_en_T_1 ? _GEN_1685 : valid_113; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2200 = _array_io_en_T_1 ? _GEN_1686 : valid_114; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2201 = _array_io_en_T_1 ? _GEN_1687 : valid_115; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2202 = _array_io_en_T_1 ? _GEN_1688 : valid_116; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2203 = _array_io_en_T_1 ? _GEN_1689 : valid_117; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2204 = _array_io_en_T_1 ? _GEN_1690 : valid_118; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2205 = _array_io_en_T_1 ? _GEN_1691 : valid_119; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2206 = _array_io_en_T_1 ? _GEN_1692 : valid_120; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2207 = _array_io_en_T_1 ? _GEN_1693 : valid_121; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2208 = _array_io_en_T_1 ? _GEN_1694 : valid_122; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2209 = _array_io_en_T_1 ? _GEN_1695 : valid_123; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2210 = _array_io_en_T_1 ? _GEN_1696 : valid_124; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2211 = _array_io_en_T_1 ? _GEN_1697 : valid_125; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2212 = _array_io_en_T_1 ? _GEN_1698 : valid_126; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2213 = _array_io_en_T_1 ? _GEN_1699 : valid_127; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2214 = _array_io_en_T_1 ? _GEN_1700 : valid_128; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2215 = _array_io_en_T_1 ? _GEN_1701 : valid_129; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2216 = _array_io_en_T_1 ? _GEN_1702 : valid_130; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2217 = _array_io_en_T_1 ? _GEN_1703 : valid_131; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2218 = _array_io_en_T_1 ? _GEN_1704 : valid_132; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2219 = _array_io_en_T_1 ? _GEN_1705 : valid_133; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2220 = _array_io_en_T_1 ? _GEN_1706 : valid_134; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2221 = _array_io_en_T_1 ? _GEN_1707 : valid_135; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2222 = _array_io_en_T_1 ? _GEN_1708 : valid_136; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2223 = _array_io_en_T_1 ? _GEN_1709 : valid_137; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2224 = _array_io_en_T_1 ? _GEN_1710 : valid_138; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2225 = _array_io_en_T_1 ? _GEN_1711 : valid_139; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2226 = _array_io_en_T_1 ? _GEN_1712 : valid_140; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2227 = _array_io_en_T_1 ? _GEN_1713 : valid_141; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2228 = _array_io_en_T_1 ? _GEN_1714 : valid_142; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2229 = _array_io_en_T_1 ? _GEN_1715 : valid_143; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2230 = _array_io_en_T_1 ? _GEN_1716 : valid_144; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2231 = _array_io_en_T_1 ? _GEN_1717 : valid_145; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2232 = _array_io_en_T_1 ? _GEN_1718 : valid_146; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2233 = _array_io_en_T_1 ? _GEN_1719 : valid_147; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2234 = _array_io_en_T_1 ? _GEN_1720 : valid_148; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2235 = _array_io_en_T_1 ? _GEN_1721 : valid_149; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2236 = _array_io_en_T_1 ? _GEN_1722 : valid_150; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2237 = _array_io_en_T_1 ? _GEN_1723 : valid_151; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2238 = _array_io_en_T_1 ? _GEN_1724 : valid_152; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2239 = _array_io_en_T_1 ? _GEN_1725 : valid_153; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2240 = _array_io_en_T_1 ? _GEN_1726 : valid_154; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2241 = _array_io_en_T_1 ? _GEN_1727 : valid_155; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2242 = _array_io_en_T_1 ? _GEN_1728 : valid_156; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2243 = _array_io_en_T_1 ? _GEN_1729 : valid_157; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2244 = _array_io_en_T_1 ? _GEN_1730 : valid_158; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2245 = _array_io_en_T_1 ? _GEN_1731 : valid_159; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2246 = _array_io_en_T_1 ? _GEN_1732 : valid_160; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2247 = _array_io_en_T_1 ? _GEN_1733 : valid_161; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2248 = _array_io_en_T_1 ? _GEN_1734 : valid_162; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2249 = _array_io_en_T_1 ? _GEN_1735 : valid_163; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2250 = _array_io_en_T_1 ? _GEN_1736 : valid_164; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2251 = _array_io_en_T_1 ? _GEN_1737 : valid_165; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2252 = _array_io_en_T_1 ? _GEN_1738 : valid_166; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2253 = _array_io_en_T_1 ? _GEN_1739 : valid_167; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2254 = _array_io_en_T_1 ? _GEN_1740 : valid_168; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2255 = _array_io_en_T_1 ? _GEN_1741 : valid_169; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2256 = _array_io_en_T_1 ? _GEN_1742 : valid_170; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2257 = _array_io_en_T_1 ? _GEN_1743 : valid_171; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2258 = _array_io_en_T_1 ? _GEN_1744 : valid_172; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2259 = _array_io_en_T_1 ? _GEN_1745 : valid_173; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2260 = _array_io_en_T_1 ? _GEN_1746 : valid_174; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2261 = _array_io_en_T_1 ? _GEN_1747 : valid_175; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2262 = _array_io_en_T_1 ? _GEN_1748 : valid_176; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2263 = _array_io_en_T_1 ? _GEN_1749 : valid_177; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2264 = _array_io_en_T_1 ? _GEN_1750 : valid_178; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2265 = _array_io_en_T_1 ? _GEN_1751 : valid_179; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2266 = _array_io_en_T_1 ? _GEN_1752 : valid_180; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2267 = _array_io_en_T_1 ? _GEN_1753 : valid_181; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2268 = _array_io_en_T_1 ? _GEN_1754 : valid_182; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2269 = _array_io_en_T_1 ? _GEN_1755 : valid_183; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2270 = _array_io_en_T_1 ? _GEN_1756 : valid_184; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2271 = _array_io_en_T_1 ? _GEN_1757 : valid_185; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2272 = _array_io_en_T_1 ? _GEN_1758 : valid_186; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2273 = _array_io_en_T_1 ? _GEN_1759 : valid_187; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2274 = _array_io_en_T_1 ? _GEN_1760 : valid_188; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2275 = _array_io_en_T_1 ? _GEN_1761 : valid_189; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2276 = _array_io_en_T_1 ? _GEN_1762 : valid_190; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2277 = _array_io_en_T_1 ? _GEN_1763 : valid_191; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2278 = _array_io_en_T_1 ? _GEN_1764 : valid_192; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2279 = _array_io_en_T_1 ? _GEN_1765 : valid_193; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2280 = _array_io_en_T_1 ? _GEN_1766 : valid_194; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2281 = _array_io_en_T_1 ? _GEN_1767 : valid_195; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2282 = _array_io_en_T_1 ? _GEN_1768 : valid_196; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2283 = _array_io_en_T_1 ? _GEN_1769 : valid_197; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2284 = _array_io_en_T_1 ? _GEN_1770 : valid_198; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2285 = _array_io_en_T_1 ? _GEN_1771 : valid_199; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2286 = _array_io_en_T_1 ? _GEN_1772 : valid_200; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2287 = _array_io_en_T_1 ? _GEN_1773 : valid_201; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2288 = _array_io_en_T_1 ? _GEN_1774 : valid_202; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2289 = _array_io_en_T_1 ? _GEN_1775 : valid_203; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2290 = _array_io_en_T_1 ? _GEN_1776 : valid_204; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2291 = _array_io_en_T_1 ? _GEN_1777 : valid_205; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2292 = _array_io_en_T_1 ? _GEN_1778 : valid_206; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2293 = _array_io_en_T_1 ? _GEN_1779 : valid_207; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2294 = _array_io_en_T_1 ? _GEN_1780 : valid_208; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2295 = _array_io_en_T_1 ? _GEN_1781 : valid_209; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2296 = _array_io_en_T_1 ? _GEN_1782 : valid_210; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2297 = _array_io_en_T_1 ? _GEN_1783 : valid_211; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2298 = _array_io_en_T_1 ? _GEN_1784 : valid_212; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2299 = _array_io_en_T_1 ? _GEN_1785 : valid_213; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2300 = _array_io_en_T_1 ? _GEN_1786 : valid_214; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2301 = _array_io_en_T_1 ? _GEN_1787 : valid_215; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2302 = _array_io_en_T_1 ? _GEN_1788 : valid_216; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2303 = _array_io_en_T_1 ? _GEN_1789 : valid_217; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2304 = _array_io_en_T_1 ? _GEN_1790 : valid_218; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2305 = _array_io_en_T_1 ? _GEN_1791 : valid_219; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2306 = _array_io_en_T_1 ? _GEN_1792 : valid_220; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2307 = _array_io_en_T_1 ? _GEN_1793 : valid_221; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2308 = _array_io_en_T_1 ? _GEN_1794 : valid_222; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2309 = _array_io_en_T_1 ? _GEN_1795 : valid_223; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2310 = _array_io_en_T_1 ? _GEN_1796 : valid_224; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2311 = _array_io_en_T_1 ? _GEN_1797 : valid_225; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2312 = _array_io_en_T_1 ? _GEN_1798 : valid_226; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2313 = _array_io_en_T_1 ? _GEN_1799 : valid_227; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2314 = _array_io_en_T_1 ? _GEN_1800 : valid_228; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2315 = _array_io_en_T_1 ? _GEN_1801 : valid_229; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2316 = _array_io_en_T_1 ? _GEN_1802 : valid_230; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2317 = _array_io_en_T_1 ? _GEN_1803 : valid_231; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2318 = _array_io_en_T_1 ? _GEN_1804 : valid_232; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2319 = _array_io_en_T_1 ? _GEN_1805 : valid_233; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2320 = _array_io_en_T_1 ? _GEN_1806 : valid_234; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2321 = _array_io_en_T_1 ? _GEN_1807 : valid_235; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2322 = _array_io_en_T_1 ? _GEN_1808 : valid_236; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2323 = _array_io_en_T_1 ? _GEN_1809 : valid_237; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2324 = _array_io_en_T_1 ? _GEN_1810 : valid_238; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2325 = _array_io_en_T_1 ? _GEN_1811 : valid_239; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2326 = _array_io_en_T_1 ? _GEN_1812 : valid_240; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2327 = _array_io_en_T_1 ? _GEN_1813 : valid_241; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2328 = _array_io_en_T_1 ? _GEN_1814 : valid_242; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2329 = _array_io_en_T_1 ? _GEN_1815 : valid_243; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2330 = _array_io_en_T_1 ? _GEN_1816 : valid_244; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2331 = _array_io_en_T_1 ? _GEN_1817 : valid_245; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2332 = _array_io_en_T_1 ? _GEN_1818 : valid_246; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2333 = _array_io_en_T_1 ? _GEN_1819 : valid_247; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2334 = _array_io_en_T_1 ? _GEN_1820 : valid_248; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2335 = _array_io_en_T_1 ? _GEN_1821 : valid_249; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2336 = _array_io_en_T_1 ? _GEN_1822 : valid_250; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2337 = _array_io_en_T_1 ? _GEN_1823 : valid_251; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2338 = _array_io_en_T_1 ? _GEN_1824 : valid_252; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2339 = _array_io_en_T_1 ? _GEN_1825 : valid_253; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2340 = _array_io_en_T_1 ? _GEN_1826 : valid_254; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2341 = _array_io_en_T_1 ? _GEN_1827 : valid_255; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2342 = _array_io_en_T_1 ? _GEN_1828 : valid_256; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2343 = _array_io_en_T_1 ? _GEN_1829 : valid_257; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2344 = _array_io_en_T_1 ? _GEN_1830 : valid_258; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2345 = _array_io_en_T_1 ? _GEN_1831 : valid_259; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2346 = _array_io_en_T_1 ? _GEN_1832 : valid_260; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2347 = _array_io_en_T_1 ? _GEN_1833 : valid_261; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2348 = _array_io_en_T_1 ? _GEN_1834 : valid_262; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2349 = _array_io_en_T_1 ? _GEN_1835 : valid_263; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2350 = _array_io_en_T_1 ? _GEN_1836 : valid_264; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2351 = _array_io_en_T_1 ? _GEN_1837 : valid_265; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2352 = _array_io_en_T_1 ? _GEN_1838 : valid_266; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2353 = _array_io_en_T_1 ? _GEN_1839 : valid_267; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2354 = _array_io_en_T_1 ? _GEN_1840 : valid_268; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2355 = _array_io_en_T_1 ? _GEN_1841 : valid_269; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2356 = _array_io_en_T_1 ? _GEN_1842 : valid_270; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2357 = _array_io_en_T_1 ? _GEN_1843 : valid_271; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2358 = _array_io_en_T_1 ? _GEN_1844 : valid_272; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2359 = _array_io_en_T_1 ? _GEN_1845 : valid_273; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2360 = _array_io_en_T_1 ? _GEN_1846 : valid_274; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2361 = _array_io_en_T_1 ? _GEN_1847 : valid_275; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2362 = _array_io_en_T_1 ? _GEN_1848 : valid_276; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2363 = _array_io_en_T_1 ? _GEN_1849 : valid_277; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2364 = _array_io_en_T_1 ? _GEN_1850 : valid_278; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2365 = _array_io_en_T_1 ? _GEN_1851 : valid_279; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2366 = _array_io_en_T_1 ? _GEN_1852 : valid_280; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2367 = _array_io_en_T_1 ? _GEN_1853 : valid_281; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2368 = _array_io_en_T_1 ? _GEN_1854 : valid_282; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2369 = _array_io_en_T_1 ? _GEN_1855 : valid_283; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2370 = _array_io_en_T_1 ? _GEN_1856 : valid_284; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2371 = _array_io_en_T_1 ? _GEN_1857 : valid_285; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2372 = _array_io_en_T_1 ? _GEN_1858 : valid_286; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2373 = _array_io_en_T_1 ? _GEN_1859 : valid_287; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2374 = _array_io_en_T_1 ? _GEN_1860 : valid_288; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2375 = _array_io_en_T_1 ? _GEN_1861 : valid_289; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2376 = _array_io_en_T_1 ? _GEN_1862 : valid_290; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2377 = _array_io_en_T_1 ? _GEN_1863 : valid_291; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2378 = _array_io_en_T_1 ? _GEN_1864 : valid_292; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2379 = _array_io_en_T_1 ? _GEN_1865 : valid_293; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2380 = _array_io_en_T_1 ? _GEN_1866 : valid_294; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2381 = _array_io_en_T_1 ? _GEN_1867 : valid_295; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2382 = _array_io_en_T_1 ? _GEN_1868 : valid_296; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2383 = _array_io_en_T_1 ? _GEN_1869 : valid_297; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2384 = _array_io_en_T_1 ? _GEN_1870 : valid_298; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2385 = _array_io_en_T_1 ? _GEN_1871 : valid_299; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2386 = _array_io_en_T_1 ? _GEN_1872 : valid_300; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2387 = _array_io_en_T_1 ? _GEN_1873 : valid_301; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2388 = _array_io_en_T_1 ? _GEN_1874 : valid_302; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2389 = _array_io_en_T_1 ? _GEN_1875 : valid_303; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2390 = _array_io_en_T_1 ? _GEN_1876 : valid_304; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2391 = _array_io_en_T_1 ? _GEN_1877 : valid_305; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2392 = _array_io_en_T_1 ? _GEN_1878 : valid_306; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2393 = _array_io_en_T_1 ? _GEN_1879 : valid_307; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2394 = _array_io_en_T_1 ? _GEN_1880 : valid_308; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2395 = _array_io_en_T_1 ? _GEN_1881 : valid_309; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2396 = _array_io_en_T_1 ? _GEN_1882 : valid_310; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2397 = _array_io_en_T_1 ? _GEN_1883 : valid_311; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2398 = _array_io_en_T_1 ? _GEN_1884 : valid_312; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2399 = _array_io_en_T_1 ? _GEN_1885 : valid_313; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2400 = _array_io_en_T_1 ? _GEN_1886 : valid_314; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2401 = _array_io_en_T_1 ? _GEN_1887 : valid_315; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2402 = _array_io_en_T_1 ? _GEN_1888 : valid_316; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2403 = _array_io_en_T_1 ? _GEN_1889 : valid_317; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2404 = _array_io_en_T_1 ? _GEN_1890 : valid_318; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2405 = _array_io_en_T_1 ? _GEN_1891 : valid_319; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2406 = _array_io_en_T_1 ? _GEN_1892 : valid_320; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2407 = _array_io_en_T_1 ? _GEN_1893 : valid_321; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2408 = _array_io_en_T_1 ? _GEN_1894 : valid_322; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2409 = _array_io_en_T_1 ? _GEN_1895 : valid_323; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2410 = _array_io_en_T_1 ? _GEN_1896 : valid_324; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2411 = _array_io_en_T_1 ? _GEN_1897 : valid_325; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2412 = _array_io_en_T_1 ? _GEN_1898 : valid_326; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2413 = _array_io_en_T_1 ? _GEN_1899 : valid_327; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2414 = _array_io_en_T_1 ? _GEN_1900 : valid_328; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2415 = _array_io_en_T_1 ? _GEN_1901 : valid_329; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2416 = _array_io_en_T_1 ? _GEN_1902 : valid_330; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2417 = _array_io_en_T_1 ? _GEN_1903 : valid_331; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2418 = _array_io_en_T_1 ? _GEN_1904 : valid_332; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2419 = _array_io_en_T_1 ? _GEN_1905 : valid_333; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2420 = _array_io_en_T_1 ? _GEN_1906 : valid_334; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2421 = _array_io_en_T_1 ? _GEN_1907 : valid_335; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2422 = _array_io_en_T_1 ? _GEN_1908 : valid_336; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2423 = _array_io_en_T_1 ? _GEN_1909 : valid_337; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2424 = _array_io_en_T_1 ? _GEN_1910 : valid_338; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2425 = _array_io_en_T_1 ? _GEN_1911 : valid_339; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2426 = _array_io_en_T_1 ? _GEN_1912 : valid_340; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2427 = _array_io_en_T_1 ? _GEN_1913 : valid_341; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2428 = _array_io_en_T_1 ? _GEN_1914 : valid_342; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2429 = _array_io_en_T_1 ? _GEN_1915 : valid_343; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2430 = _array_io_en_T_1 ? _GEN_1916 : valid_344; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2431 = _array_io_en_T_1 ? _GEN_1917 : valid_345; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2432 = _array_io_en_T_1 ? _GEN_1918 : valid_346; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2433 = _array_io_en_T_1 ? _GEN_1919 : valid_347; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2434 = _array_io_en_T_1 ? _GEN_1920 : valid_348; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2435 = _array_io_en_T_1 ? _GEN_1921 : valid_349; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2436 = _array_io_en_T_1 ? _GEN_1922 : valid_350; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2437 = _array_io_en_T_1 ? _GEN_1923 : valid_351; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2438 = _array_io_en_T_1 ? _GEN_1924 : valid_352; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2439 = _array_io_en_T_1 ? _GEN_1925 : valid_353; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2440 = _array_io_en_T_1 ? _GEN_1926 : valid_354; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2441 = _array_io_en_T_1 ? _GEN_1927 : valid_355; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2442 = _array_io_en_T_1 ? _GEN_1928 : valid_356; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2443 = _array_io_en_T_1 ? _GEN_1929 : valid_357; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2444 = _array_io_en_T_1 ? _GEN_1930 : valid_358; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2445 = _array_io_en_T_1 ? _GEN_1931 : valid_359; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2446 = _array_io_en_T_1 ? _GEN_1932 : valid_360; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2447 = _array_io_en_T_1 ? _GEN_1933 : valid_361; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2448 = _array_io_en_T_1 ? _GEN_1934 : valid_362; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2449 = _array_io_en_T_1 ? _GEN_1935 : valid_363; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2450 = _array_io_en_T_1 ? _GEN_1936 : valid_364; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2451 = _array_io_en_T_1 ? _GEN_1937 : valid_365; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2452 = _array_io_en_T_1 ? _GEN_1938 : valid_366; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2453 = _array_io_en_T_1 ? _GEN_1939 : valid_367; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2454 = _array_io_en_T_1 ? _GEN_1940 : valid_368; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2455 = _array_io_en_T_1 ? _GEN_1941 : valid_369; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2456 = _array_io_en_T_1 ? _GEN_1942 : valid_370; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2457 = _array_io_en_T_1 ? _GEN_1943 : valid_371; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2458 = _array_io_en_T_1 ? _GEN_1944 : valid_372; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2459 = _array_io_en_T_1 ? _GEN_1945 : valid_373; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2460 = _array_io_en_T_1 ? _GEN_1946 : valid_374; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2461 = _array_io_en_T_1 ? _GEN_1947 : valid_375; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2462 = _array_io_en_T_1 ? _GEN_1948 : valid_376; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2463 = _array_io_en_T_1 ? _GEN_1949 : valid_377; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2464 = _array_io_en_T_1 ? _GEN_1950 : valid_378; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2465 = _array_io_en_T_1 ? _GEN_1951 : valid_379; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2466 = _array_io_en_T_1 ? _GEN_1952 : valid_380; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2467 = _array_io_en_T_1 ? _GEN_1953 : valid_381; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2468 = _array_io_en_T_1 ? _GEN_1954 : valid_382; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2469 = _array_io_en_T_1 ? _GEN_1955 : valid_383; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2470 = _array_io_en_T_1 ? _GEN_1956 : valid_384; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2471 = _array_io_en_T_1 ? _GEN_1957 : valid_385; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2472 = _array_io_en_T_1 ? _GEN_1958 : valid_386; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2473 = _array_io_en_T_1 ? _GEN_1959 : valid_387; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2474 = _array_io_en_T_1 ? _GEN_1960 : valid_388; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2475 = _array_io_en_T_1 ? _GEN_1961 : valid_389; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2476 = _array_io_en_T_1 ? _GEN_1962 : valid_390; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2477 = _array_io_en_T_1 ? _GEN_1963 : valid_391; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2478 = _array_io_en_T_1 ? _GEN_1964 : valid_392; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2479 = _array_io_en_T_1 ? _GEN_1965 : valid_393; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2480 = _array_io_en_T_1 ? _GEN_1966 : valid_394; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2481 = _array_io_en_T_1 ? _GEN_1967 : valid_395; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2482 = _array_io_en_T_1 ? _GEN_1968 : valid_396; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2483 = _array_io_en_T_1 ? _GEN_1969 : valid_397; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2484 = _array_io_en_T_1 ? _GEN_1970 : valid_398; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2485 = _array_io_en_T_1 ? _GEN_1971 : valid_399; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2486 = _array_io_en_T_1 ? _GEN_1972 : valid_400; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2487 = _array_io_en_T_1 ? _GEN_1973 : valid_401; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2488 = _array_io_en_T_1 ? _GEN_1974 : valid_402; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2489 = _array_io_en_T_1 ? _GEN_1975 : valid_403; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2490 = _array_io_en_T_1 ? _GEN_1976 : valid_404; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2491 = _array_io_en_T_1 ? _GEN_1977 : valid_405; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2492 = _array_io_en_T_1 ? _GEN_1978 : valid_406; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2493 = _array_io_en_T_1 ? _GEN_1979 : valid_407; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2494 = _array_io_en_T_1 ? _GEN_1980 : valid_408; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2495 = _array_io_en_T_1 ? _GEN_1981 : valid_409; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2496 = _array_io_en_T_1 ? _GEN_1982 : valid_410; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2497 = _array_io_en_T_1 ? _GEN_1983 : valid_411; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2498 = _array_io_en_T_1 ? _GEN_1984 : valid_412; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2499 = _array_io_en_T_1 ? _GEN_1985 : valid_413; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2500 = _array_io_en_T_1 ? _GEN_1986 : valid_414; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2501 = _array_io_en_T_1 ? _GEN_1987 : valid_415; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2502 = _array_io_en_T_1 ? _GEN_1988 : valid_416; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2503 = _array_io_en_T_1 ? _GEN_1989 : valid_417; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2504 = _array_io_en_T_1 ? _GEN_1990 : valid_418; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2505 = _array_io_en_T_1 ? _GEN_1991 : valid_419; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2506 = _array_io_en_T_1 ? _GEN_1992 : valid_420; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2507 = _array_io_en_T_1 ? _GEN_1993 : valid_421; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2508 = _array_io_en_T_1 ? _GEN_1994 : valid_422; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2509 = _array_io_en_T_1 ? _GEN_1995 : valid_423; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2510 = _array_io_en_T_1 ? _GEN_1996 : valid_424; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2511 = _array_io_en_T_1 ? _GEN_1997 : valid_425; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2512 = _array_io_en_T_1 ? _GEN_1998 : valid_426; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2513 = _array_io_en_T_1 ? _GEN_1999 : valid_427; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2514 = _array_io_en_T_1 ? _GEN_2000 : valid_428; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2515 = _array_io_en_T_1 ? _GEN_2001 : valid_429; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2516 = _array_io_en_T_1 ? _GEN_2002 : valid_430; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2517 = _array_io_en_T_1 ? _GEN_2003 : valid_431; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2518 = _array_io_en_T_1 ? _GEN_2004 : valid_432; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2519 = _array_io_en_T_1 ? _GEN_2005 : valid_433; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2520 = _array_io_en_T_1 ? _GEN_2006 : valid_434; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2521 = _array_io_en_T_1 ? _GEN_2007 : valid_435; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2522 = _array_io_en_T_1 ? _GEN_2008 : valid_436; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2523 = _array_io_en_T_1 ? _GEN_2009 : valid_437; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2524 = _array_io_en_T_1 ? _GEN_2010 : valid_438; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2525 = _array_io_en_T_1 ? _GEN_2011 : valid_439; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2526 = _array_io_en_T_1 ? _GEN_2012 : valid_440; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2527 = _array_io_en_T_1 ? _GEN_2013 : valid_441; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2528 = _array_io_en_T_1 ? _GEN_2014 : valid_442; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2529 = _array_io_en_T_1 ? _GEN_2015 : valid_443; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2530 = _array_io_en_T_1 ? _GEN_2016 : valid_444; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2531 = _array_io_en_T_1 ? _GEN_2017 : valid_445; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2532 = _array_io_en_T_1 ? _GEN_2018 : valid_446; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2533 = _array_io_en_T_1 ? _GEN_2019 : valid_447; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2534 = _array_io_en_T_1 ? _GEN_2020 : valid_448; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2535 = _array_io_en_T_1 ? _GEN_2021 : valid_449; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2536 = _array_io_en_T_1 ? _GEN_2022 : valid_450; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2537 = _array_io_en_T_1 ? _GEN_2023 : valid_451; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2538 = _array_io_en_T_1 ? _GEN_2024 : valid_452; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2539 = _array_io_en_T_1 ? _GEN_2025 : valid_453; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2540 = _array_io_en_T_1 ? _GEN_2026 : valid_454; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2541 = _array_io_en_T_1 ? _GEN_2027 : valid_455; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2542 = _array_io_en_T_1 ? _GEN_2028 : valid_456; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2543 = _array_io_en_T_1 ? _GEN_2029 : valid_457; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2544 = _array_io_en_T_1 ? _GEN_2030 : valid_458; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2545 = _array_io_en_T_1 ? _GEN_2031 : valid_459; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2546 = _array_io_en_T_1 ? _GEN_2032 : valid_460; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2547 = _array_io_en_T_1 ? _GEN_2033 : valid_461; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2548 = _array_io_en_T_1 ? _GEN_2034 : valid_462; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2549 = _array_io_en_T_1 ? _GEN_2035 : valid_463; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2550 = _array_io_en_T_1 ? _GEN_2036 : valid_464; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2551 = _array_io_en_T_1 ? _GEN_2037 : valid_465; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2552 = _array_io_en_T_1 ? _GEN_2038 : valid_466; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2553 = _array_io_en_T_1 ? _GEN_2039 : valid_467; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2554 = _array_io_en_T_1 ? _GEN_2040 : valid_468; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2555 = _array_io_en_T_1 ? _GEN_2041 : valid_469; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2556 = _array_io_en_T_1 ? _GEN_2042 : valid_470; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2557 = _array_io_en_T_1 ? _GEN_2043 : valid_471; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2558 = _array_io_en_T_1 ? _GEN_2044 : valid_472; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2559 = _array_io_en_T_1 ? _GEN_2045 : valid_473; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2560 = _array_io_en_T_1 ? _GEN_2046 : valid_474; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2561 = _array_io_en_T_1 ? _GEN_2047 : valid_475; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2562 = _array_io_en_T_1 ? _GEN_2048 : valid_476; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2563 = _array_io_en_T_1 ? _GEN_2049 : valid_477; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2564 = _array_io_en_T_1 ? _GEN_2050 : valid_478; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2565 = _array_io_en_T_1 ? _GEN_2051 : valid_479; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2566 = _array_io_en_T_1 ? _GEN_2052 : valid_480; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2567 = _array_io_en_T_1 ? _GEN_2053 : valid_481; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2568 = _array_io_en_T_1 ? _GEN_2054 : valid_482; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2569 = _array_io_en_T_1 ? _GEN_2055 : valid_483; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2570 = _array_io_en_T_1 ? _GEN_2056 : valid_484; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2571 = _array_io_en_T_1 ? _GEN_2057 : valid_485; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2572 = _array_io_en_T_1 ? _GEN_2058 : valid_486; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2573 = _array_io_en_T_1 ? _GEN_2059 : valid_487; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2574 = _array_io_en_T_1 ? _GEN_2060 : valid_488; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2575 = _array_io_en_T_1 ? _GEN_2061 : valid_489; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2576 = _array_io_en_T_1 ? _GEN_2062 : valid_490; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2577 = _array_io_en_T_1 ? _GEN_2063 : valid_491; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2578 = _array_io_en_T_1 ? _GEN_2064 : valid_492; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2579 = _array_io_en_T_1 ? _GEN_2065 : valid_493; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2580 = _array_io_en_T_1 ? _GEN_2066 : valid_494; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2581 = _array_io_en_T_1 ? _GEN_2067 : valid_495; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2582 = _array_io_en_T_1 ? _GEN_2068 : valid_496; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2583 = _array_io_en_T_1 ? _GEN_2069 : valid_497; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2584 = _array_io_en_T_1 ? _GEN_2070 : valid_498; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2585 = _array_io_en_T_1 ? _GEN_2071 : valid_499; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2586 = _array_io_en_T_1 ? _GEN_2072 : valid_500; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2587 = _array_io_en_T_1 ? _GEN_2073 : valid_501; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2588 = _array_io_en_T_1 ? _GEN_2074 : valid_502; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2589 = _array_io_en_T_1 ? _GEN_2075 : valid_503; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2590 = _array_io_en_T_1 ? _GEN_2076 : valid_504; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2591 = _array_io_en_T_1 ? _GEN_2077 : valid_505; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2592 = _array_io_en_T_1 ? _GEN_2078 : valid_506; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2593 = _array_io_en_T_1 ? _GEN_2079 : valid_507; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2594 = _array_io_en_T_1 ? _GEN_2080 : valid_508; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2595 = _array_io_en_T_1 ? _GEN_2081 : valid_509; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2596 = _array_io_en_T_1 ? _GEN_2082 : valid_510; // @[DCache.scala 164:19 56:22]
  wire  _GEN_2597 = _array_io_en_T_1 ? _GEN_2083 : valid_511; // @[DCache.scala 164:19 56:22]
  wire  tl_c_valid = probing | state == 3'h2 & _GEN_535; // @[DCache.scala 260:25]
  wire  _probing_T_1 = auto_out_c_ready & tl_c_valid; // @[Decoupled.scala 51:35]
  wire  _GEN_2598 = _probing_T_1 ? 1'h0 : probing; // @[Utils.scala 38:18 36:20 38:22]
  wire  _GEN_2599 = _tl_b_bits_r_T | _GEN_2598; // @[Utils.scala 39:{19,23}]
  wire [2:0] _state_T_1 = _GEN_535 ? 3'h2 : 3'h4; // @[DCache.scala 194:21]
  wire [2:0] _GEN_2601 = ~array_hit ? _state_T_1 : state; // @[DCache.scala 193:30 194:15 60:118]
  wire [2:0] _GEN_2603 = _probing_T_1 & _x1_b_ready_T ? 3'h3 : state; // @[DCache.scala 200:41 201:15 60:118]
  wire [2:0] _GEN_2604 = ~_GEN_535 ? 3'h4 : _GEN_2603; // @[DCache.scala 198:26 199:15]
  wire [2:0] _GEN_2605 = _tl_d_bits_r_T ? 3'h4 : state; // @[DCache.scala 205:23 206:15 60:118]
  wire  tl_a_valid = state == 3'h4; // @[DCache.scala 257:24]
  wire  _T_27 = auto_out_a_ready & tl_a_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_2606 = _T_27 ? 3'h5 : state; // @[DCache.scala 210:23 211:15 60:118]
  wire [2:0] _GEN_2607 = _tl_d_bits_r_T ? 3'h6 : state; // @[DCache.scala 215:23 216:15 60:118]
  wire  tl_e_valid = state == 3'h6; // @[DCache.scala 263:24]
  wire  _T_31 = auto_out_e_ready & tl_e_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_2608 = _T_31 ? 3'h7 : state; // @[DCache.scala 220:23 221:15 60:118]
  wire [2:0] _GEN_2609 = _array_io_en_T_1 ? 3'h0 : state; // @[DCache.scala 225:23 226:15 60:118]
  wire [2:0] _GEN_2610 = 3'h7 == state ? _GEN_2609 : state; // @[DCache.scala 184:17 60:118]
  wire [2:0] _GEN_2611 = 3'h6 == state ? _GEN_2608 : _GEN_2610; // @[DCache.scala 184:17]
  wire [2:0] _GEN_2612 = 3'h5 == state ? _GEN_2607 : _GEN_2611; // @[DCache.scala 184:17]
  wire [2:0] _GEN_2613 = 3'h4 == state ? _GEN_2606 : _GEN_2612; // @[DCache.scala 184:17]
  wire [2:0] _GEN_2614 = 3'h3 == state ? _GEN_2605 : _GEN_2613; // @[DCache.scala 184:17]
  reg  probe_out_REG; // @[DCache.scala 233:54]
  reg [273:0] probe_out_r; // @[Reg.scala 35:20]
  wire [273:0] _GEN_2618 = probe_out_REG ? array_io_rdata : probe_out_r; // @[Reg.scala 36:18 35:20 36:22]
  wire [255:0] probe_out_data = _GEN_2618[255:0]; // @[DCache.scala 233:75]
  wire [17:0] probe_out_tag = _GEN_2618[273:256]; // @[DCache.scala 233:75]
  wire  _GEN_2620 = 9'h1 == _GEN_4[13:5] ? valid_1 : valid_0; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2621 = 9'h2 == _GEN_4[13:5] ? valid_2 : _GEN_2620; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2622 = 9'h3 == _GEN_4[13:5] ? valid_3 : _GEN_2621; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2623 = 9'h4 == _GEN_4[13:5] ? valid_4 : _GEN_2622; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2624 = 9'h5 == _GEN_4[13:5] ? valid_5 : _GEN_2623; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2625 = 9'h6 == _GEN_4[13:5] ? valid_6 : _GEN_2624; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2626 = 9'h7 == _GEN_4[13:5] ? valid_7 : _GEN_2625; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2627 = 9'h8 == _GEN_4[13:5] ? valid_8 : _GEN_2626; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2628 = 9'h9 == _GEN_4[13:5] ? valid_9 : _GEN_2627; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2629 = 9'ha == _GEN_4[13:5] ? valid_10 : _GEN_2628; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2630 = 9'hb == _GEN_4[13:5] ? valid_11 : _GEN_2629; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2631 = 9'hc == _GEN_4[13:5] ? valid_12 : _GEN_2630; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2632 = 9'hd == _GEN_4[13:5] ? valid_13 : _GEN_2631; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2633 = 9'he == _GEN_4[13:5] ? valid_14 : _GEN_2632; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2634 = 9'hf == _GEN_4[13:5] ? valid_15 : _GEN_2633; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2635 = 9'h10 == _GEN_4[13:5] ? valid_16 : _GEN_2634; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2636 = 9'h11 == _GEN_4[13:5] ? valid_17 : _GEN_2635; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2637 = 9'h12 == _GEN_4[13:5] ? valid_18 : _GEN_2636; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2638 = 9'h13 == _GEN_4[13:5] ? valid_19 : _GEN_2637; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2639 = 9'h14 == _GEN_4[13:5] ? valid_20 : _GEN_2638; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2640 = 9'h15 == _GEN_4[13:5] ? valid_21 : _GEN_2639; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2641 = 9'h16 == _GEN_4[13:5] ? valid_22 : _GEN_2640; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2642 = 9'h17 == _GEN_4[13:5] ? valid_23 : _GEN_2641; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2643 = 9'h18 == _GEN_4[13:5] ? valid_24 : _GEN_2642; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2644 = 9'h19 == _GEN_4[13:5] ? valid_25 : _GEN_2643; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2645 = 9'h1a == _GEN_4[13:5] ? valid_26 : _GEN_2644; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2646 = 9'h1b == _GEN_4[13:5] ? valid_27 : _GEN_2645; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2647 = 9'h1c == _GEN_4[13:5] ? valid_28 : _GEN_2646; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2648 = 9'h1d == _GEN_4[13:5] ? valid_29 : _GEN_2647; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2649 = 9'h1e == _GEN_4[13:5] ? valid_30 : _GEN_2648; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2650 = 9'h1f == _GEN_4[13:5] ? valid_31 : _GEN_2649; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2651 = 9'h20 == _GEN_4[13:5] ? valid_32 : _GEN_2650; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2652 = 9'h21 == _GEN_4[13:5] ? valid_33 : _GEN_2651; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2653 = 9'h22 == _GEN_4[13:5] ? valid_34 : _GEN_2652; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2654 = 9'h23 == _GEN_4[13:5] ? valid_35 : _GEN_2653; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2655 = 9'h24 == _GEN_4[13:5] ? valid_36 : _GEN_2654; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2656 = 9'h25 == _GEN_4[13:5] ? valid_37 : _GEN_2655; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2657 = 9'h26 == _GEN_4[13:5] ? valid_38 : _GEN_2656; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2658 = 9'h27 == _GEN_4[13:5] ? valid_39 : _GEN_2657; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2659 = 9'h28 == _GEN_4[13:5] ? valid_40 : _GEN_2658; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2660 = 9'h29 == _GEN_4[13:5] ? valid_41 : _GEN_2659; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2661 = 9'h2a == _GEN_4[13:5] ? valid_42 : _GEN_2660; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2662 = 9'h2b == _GEN_4[13:5] ? valid_43 : _GEN_2661; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2663 = 9'h2c == _GEN_4[13:5] ? valid_44 : _GEN_2662; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2664 = 9'h2d == _GEN_4[13:5] ? valid_45 : _GEN_2663; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2665 = 9'h2e == _GEN_4[13:5] ? valid_46 : _GEN_2664; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2666 = 9'h2f == _GEN_4[13:5] ? valid_47 : _GEN_2665; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2667 = 9'h30 == _GEN_4[13:5] ? valid_48 : _GEN_2666; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2668 = 9'h31 == _GEN_4[13:5] ? valid_49 : _GEN_2667; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2669 = 9'h32 == _GEN_4[13:5] ? valid_50 : _GEN_2668; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2670 = 9'h33 == _GEN_4[13:5] ? valid_51 : _GEN_2669; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2671 = 9'h34 == _GEN_4[13:5] ? valid_52 : _GEN_2670; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2672 = 9'h35 == _GEN_4[13:5] ? valid_53 : _GEN_2671; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2673 = 9'h36 == _GEN_4[13:5] ? valid_54 : _GEN_2672; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2674 = 9'h37 == _GEN_4[13:5] ? valid_55 : _GEN_2673; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2675 = 9'h38 == _GEN_4[13:5] ? valid_56 : _GEN_2674; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2676 = 9'h39 == _GEN_4[13:5] ? valid_57 : _GEN_2675; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2677 = 9'h3a == _GEN_4[13:5] ? valid_58 : _GEN_2676; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2678 = 9'h3b == _GEN_4[13:5] ? valid_59 : _GEN_2677; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2679 = 9'h3c == _GEN_4[13:5] ? valid_60 : _GEN_2678; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2680 = 9'h3d == _GEN_4[13:5] ? valid_61 : _GEN_2679; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2681 = 9'h3e == _GEN_4[13:5] ? valid_62 : _GEN_2680; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2682 = 9'h3f == _GEN_4[13:5] ? valid_63 : _GEN_2681; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2683 = 9'h40 == _GEN_4[13:5] ? valid_64 : _GEN_2682; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2684 = 9'h41 == _GEN_4[13:5] ? valid_65 : _GEN_2683; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2685 = 9'h42 == _GEN_4[13:5] ? valid_66 : _GEN_2684; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2686 = 9'h43 == _GEN_4[13:5] ? valid_67 : _GEN_2685; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2687 = 9'h44 == _GEN_4[13:5] ? valid_68 : _GEN_2686; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2688 = 9'h45 == _GEN_4[13:5] ? valid_69 : _GEN_2687; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2689 = 9'h46 == _GEN_4[13:5] ? valid_70 : _GEN_2688; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2690 = 9'h47 == _GEN_4[13:5] ? valid_71 : _GEN_2689; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2691 = 9'h48 == _GEN_4[13:5] ? valid_72 : _GEN_2690; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2692 = 9'h49 == _GEN_4[13:5] ? valid_73 : _GEN_2691; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2693 = 9'h4a == _GEN_4[13:5] ? valid_74 : _GEN_2692; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2694 = 9'h4b == _GEN_4[13:5] ? valid_75 : _GEN_2693; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2695 = 9'h4c == _GEN_4[13:5] ? valid_76 : _GEN_2694; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2696 = 9'h4d == _GEN_4[13:5] ? valid_77 : _GEN_2695; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2697 = 9'h4e == _GEN_4[13:5] ? valid_78 : _GEN_2696; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2698 = 9'h4f == _GEN_4[13:5] ? valid_79 : _GEN_2697; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2699 = 9'h50 == _GEN_4[13:5] ? valid_80 : _GEN_2698; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2700 = 9'h51 == _GEN_4[13:5] ? valid_81 : _GEN_2699; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2701 = 9'h52 == _GEN_4[13:5] ? valid_82 : _GEN_2700; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2702 = 9'h53 == _GEN_4[13:5] ? valid_83 : _GEN_2701; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2703 = 9'h54 == _GEN_4[13:5] ? valid_84 : _GEN_2702; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2704 = 9'h55 == _GEN_4[13:5] ? valid_85 : _GEN_2703; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2705 = 9'h56 == _GEN_4[13:5] ? valid_86 : _GEN_2704; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2706 = 9'h57 == _GEN_4[13:5] ? valid_87 : _GEN_2705; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2707 = 9'h58 == _GEN_4[13:5] ? valid_88 : _GEN_2706; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2708 = 9'h59 == _GEN_4[13:5] ? valid_89 : _GEN_2707; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2709 = 9'h5a == _GEN_4[13:5] ? valid_90 : _GEN_2708; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2710 = 9'h5b == _GEN_4[13:5] ? valid_91 : _GEN_2709; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2711 = 9'h5c == _GEN_4[13:5] ? valid_92 : _GEN_2710; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2712 = 9'h5d == _GEN_4[13:5] ? valid_93 : _GEN_2711; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2713 = 9'h5e == _GEN_4[13:5] ? valid_94 : _GEN_2712; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2714 = 9'h5f == _GEN_4[13:5] ? valid_95 : _GEN_2713; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2715 = 9'h60 == _GEN_4[13:5] ? valid_96 : _GEN_2714; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2716 = 9'h61 == _GEN_4[13:5] ? valid_97 : _GEN_2715; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2717 = 9'h62 == _GEN_4[13:5] ? valid_98 : _GEN_2716; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2718 = 9'h63 == _GEN_4[13:5] ? valid_99 : _GEN_2717; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2719 = 9'h64 == _GEN_4[13:5] ? valid_100 : _GEN_2718; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2720 = 9'h65 == _GEN_4[13:5] ? valid_101 : _GEN_2719; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2721 = 9'h66 == _GEN_4[13:5] ? valid_102 : _GEN_2720; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2722 = 9'h67 == _GEN_4[13:5] ? valid_103 : _GEN_2721; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2723 = 9'h68 == _GEN_4[13:5] ? valid_104 : _GEN_2722; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2724 = 9'h69 == _GEN_4[13:5] ? valid_105 : _GEN_2723; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2725 = 9'h6a == _GEN_4[13:5] ? valid_106 : _GEN_2724; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2726 = 9'h6b == _GEN_4[13:5] ? valid_107 : _GEN_2725; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2727 = 9'h6c == _GEN_4[13:5] ? valid_108 : _GEN_2726; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2728 = 9'h6d == _GEN_4[13:5] ? valid_109 : _GEN_2727; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2729 = 9'h6e == _GEN_4[13:5] ? valid_110 : _GEN_2728; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2730 = 9'h6f == _GEN_4[13:5] ? valid_111 : _GEN_2729; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2731 = 9'h70 == _GEN_4[13:5] ? valid_112 : _GEN_2730; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2732 = 9'h71 == _GEN_4[13:5] ? valid_113 : _GEN_2731; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2733 = 9'h72 == _GEN_4[13:5] ? valid_114 : _GEN_2732; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2734 = 9'h73 == _GEN_4[13:5] ? valid_115 : _GEN_2733; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2735 = 9'h74 == _GEN_4[13:5] ? valid_116 : _GEN_2734; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2736 = 9'h75 == _GEN_4[13:5] ? valid_117 : _GEN_2735; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2737 = 9'h76 == _GEN_4[13:5] ? valid_118 : _GEN_2736; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2738 = 9'h77 == _GEN_4[13:5] ? valid_119 : _GEN_2737; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2739 = 9'h78 == _GEN_4[13:5] ? valid_120 : _GEN_2738; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2740 = 9'h79 == _GEN_4[13:5] ? valid_121 : _GEN_2739; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2741 = 9'h7a == _GEN_4[13:5] ? valid_122 : _GEN_2740; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2742 = 9'h7b == _GEN_4[13:5] ? valid_123 : _GEN_2741; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2743 = 9'h7c == _GEN_4[13:5] ? valid_124 : _GEN_2742; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2744 = 9'h7d == _GEN_4[13:5] ? valid_125 : _GEN_2743; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2745 = 9'h7e == _GEN_4[13:5] ? valid_126 : _GEN_2744; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2746 = 9'h7f == _GEN_4[13:5] ? valid_127 : _GEN_2745; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2747 = 9'h80 == _GEN_4[13:5] ? valid_128 : _GEN_2746; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2748 = 9'h81 == _GEN_4[13:5] ? valid_129 : _GEN_2747; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2749 = 9'h82 == _GEN_4[13:5] ? valid_130 : _GEN_2748; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2750 = 9'h83 == _GEN_4[13:5] ? valid_131 : _GEN_2749; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2751 = 9'h84 == _GEN_4[13:5] ? valid_132 : _GEN_2750; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2752 = 9'h85 == _GEN_4[13:5] ? valid_133 : _GEN_2751; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2753 = 9'h86 == _GEN_4[13:5] ? valid_134 : _GEN_2752; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2754 = 9'h87 == _GEN_4[13:5] ? valid_135 : _GEN_2753; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2755 = 9'h88 == _GEN_4[13:5] ? valid_136 : _GEN_2754; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2756 = 9'h89 == _GEN_4[13:5] ? valid_137 : _GEN_2755; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2757 = 9'h8a == _GEN_4[13:5] ? valid_138 : _GEN_2756; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2758 = 9'h8b == _GEN_4[13:5] ? valid_139 : _GEN_2757; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2759 = 9'h8c == _GEN_4[13:5] ? valid_140 : _GEN_2758; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2760 = 9'h8d == _GEN_4[13:5] ? valid_141 : _GEN_2759; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2761 = 9'h8e == _GEN_4[13:5] ? valid_142 : _GEN_2760; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2762 = 9'h8f == _GEN_4[13:5] ? valid_143 : _GEN_2761; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2763 = 9'h90 == _GEN_4[13:5] ? valid_144 : _GEN_2762; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2764 = 9'h91 == _GEN_4[13:5] ? valid_145 : _GEN_2763; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2765 = 9'h92 == _GEN_4[13:5] ? valid_146 : _GEN_2764; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2766 = 9'h93 == _GEN_4[13:5] ? valid_147 : _GEN_2765; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2767 = 9'h94 == _GEN_4[13:5] ? valid_148 : _GEN_2766; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2768 = 9'h95 == _GEN_4[13:5] ? valid_149 : _GEN_2767; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2769 = 9'h96 == _GEN_4[13:5] ? valid_150 : _GEN_2768; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2770 = 9'h97 == _GEN_4[13:5] ? valid_151 : _GEN_2769; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2771 = 9'h98 == _GEN_4[13:5] ? valid_152 : _GEN_2770; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2772 = 9'h99 == _GEN_4[13:5] ? valid_153 : _GEN_2771; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2773 = 9'h9a == _GEN_4[13:5] ? valid_154 : _GEN_2772; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2774 = 9'h9b == _GEN_4[13:5] ? valid_155 : _GEN_2773; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2775 = 9'h9c == _GEN_4[13:5] ? valid_156 : _GEN_2774; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2776 = 9'h9d == _GEN_4[13:5] ? valid_157 : _GEN_2775; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2777 = 9'h9e == _GEN_4[13:5] ? valid_158 : _GEN_2776; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2778 = 9'h9f == _GEN_4[13:5] ? valid_159 : _GEN_2777; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2779 = 9'ha0 == _GEN_4[13:5] ? valid_160 : _GEN_2778; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2780 = 9'ha1 == _GEN_4[13:5] ? valid_161 : _GEN_2779; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2781 = 9'ha2 == _GEN_4[13:5] ? valid_162 : _GEN_2780; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2782 = 9'ha3 == _GEN_4[13:5] ? valid_163 : _GEN_2781; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2783 = 9'ha4 == _GEN_4[13:5] ? valid_164 : _GEN_2782; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2784 = 9'ha5 == _GEN_4[13:5] ? valid_165 : _GEN_2783; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2785 = 9'ha6 == _GEN_4[13:5] ? valid_166 : _GEN_2784; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2786 = 9'ha7 == _GEN_4[13:5] ? valid_167 : _GEN_2785; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2787 = 9'ha8 == _GEN_4[13:5] ? valid_168 : _GEN_2786; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2788 = 9'ha9 == _GEN_4[13:5] ? valid_169 : _GEN_2787; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2789 = 9'haa == _GEN_4[13:5] ? valid_170 : _GEN_2788; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2790 = 9'hab == _GEN_4[13:5] ? valid_171 : _GEN_2789; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2791 = 9'hac == _GEN_4[13:5] ? valid_172 : _GEN_2790; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2792 = 9'had == _GEN_4[13:5] ? valid_173 : _GEN_2791; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2793 = 9'hae == _GEN_4[13:5] ? valid_174 : _GEN_2792; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2794 = 9'haf == _GEN_4[13:5] ? valid_175 : _GEN_2793; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2795 = 9'hb0 == _GEN_4[13:5] ? valid_176 : _GEN_2794; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2796 = 9'hb1 == _GEN_4[13:5] ? valid_177 : _GEN_2795; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2797 = 9'hb2 == _GEN_4[13:5] ? valid_178 : _GEN_2796; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2798 = 9'hb3 == _GEN_4[13:5] ? valid_179 : _GEN_2797; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2799 = 9'hb4 == _GEN_4[13:5] ? valid_180 : _GEN_2798; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2800 = 9'hb5 == _GEN_4[13:5] ? valid_181 : _GEN_2799; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2801 = 9'hb6 == _GEN_4[13:5] ? valid_182 : _GEN_2800; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2802 = 9'hb7 == _GEN_4[13:5] ? valid_183 : _GEN_2801; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2803 = 9'hb8 == _GEN_4[13:5] ? valid_184 : _GEN_2802; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2804 = 9'hb9 == _GEN_4[13:5] ? valid_185 : _GEN_2803; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2805 = 9'hba == _GEN_4[13:5] ? valid_186 : _GEN_2804; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2806 = 9'hbb == _GEN_4[13:5] ? valid_187 : _GEN_2805; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2807 = 9'hbc == _GEN_4[13:5] ? valid_188 : _GEN_2806; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2808 = 9'hbd == _GEN_4[13:5] ? valid_189 : _GEN_2807; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2809 = 9'hbe == _GEN_4[13:5] ? valid_190 : _GEN_2808; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2810 = 9'hbf == _GEN_4[13:5] ? valid_191 : _GEN_2809; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2811 = 9'hc0 == _GEN_4[13:5] ? valid_192 : _GEN_2810; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2812 = 9'hc1 == _GEN_4[13:5] ? valid_193 : _GEN_2811; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2813 = 9'hc2 == _GEN_4[13:5] ? valid_194 : _GEN_2812; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2814 = 9'hc3 == _GEN_4[13:5] ? valid_195 : _GEN_2813; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2815 = 9'hc4 == _GEN_4[13:5] ? valid_196 : _GEN_2814; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2816 = 9'hc5 == _GEN_4[13:5] ? valid_197 : _GEN_2815; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2817 = 9'hc6 == _GEN_4[13:5] ? valid_198 : _GEN_2816; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2818 = 9'hc7 == _GEN_4[13:5] ? valid_199 : _GEN_2817; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2819 = 9'hc8 == _GEN_4[13:5] ? valid_200 : _GEN_2818; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2820 = 9'hc9 == _GEN_4[13:5] ? valid_201 : _GEN_2819; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2821 = 9'hca == _GEN_4[13:5] ? valid_202 : _GEN_2820; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2822 = 9'hcb == _GEN_4[13:5] ? valid_203 : _GEN_2821; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2823 = 9'hcc == _GEN_4[13:5] ? valid_204 : _GEN_2822; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2824 = 9'hcd == _GEN_4[13:5] ? valid_205 : _GEN_2823; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2825 = 9'hce == _GEN_4[13:5] ? valid_206 : _GEN_2824; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2826 = 9'hcf == _GEN_4[13:5] ? valid_207 : _GEN_2825; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2827 = 9'hd0 == _GEN_4[13:5] ? valid_208 : _GEN_2826; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2828 = 9'hd1 == _GEN_4[13:5] ? valid_209 : _GEN_2827; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2829 = 9'hd2 == _GEN_4[13:5] ? valid_210 : _GEN_2828; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2830 = 9'hd3 == _GEN_4[13:5] ? valid_211 : _GEN_2829; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2831 = 9'hd4 == _GEN_4[13:5] ? valid_212 : _GEN_2830; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2832 = 9'hd5 == _GEN_4[13:5] ? valid_213 : _GEN_2831; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2833 = 9'hd6 == _GEN_4[13:5] ? valid_214 : _GEN_2832; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2834 = 9'hd7 == _GEN_4[13:5] ? valid_215 : _GEN_2833; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2835 = 9'hd8 == _GEN_4[13:5] ? valid_216 : _GEN_2834; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2836 = 9'hd9 == _GEN_4[13:5] ? valid_217 : _GEN_2835; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2837 = 9'hda == _GEN_4[13:5] ? valid_218 : _GEN_2836; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2838 = 9'hdb == _GEN_4[13:5] ? valid_219 : _GEN_2837; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2839 = 9'hdc == _GEN_4[13:5] ? valid_220 : _GEN_2838; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2840 = 9'hdd == _GEN_4[13:5] ? valid_221 : _GEN_2839; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2841 = 9'hde == _GEN_4[13:5] ? valid_222 : _GEN_2840; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2842 = 9'hdf == _GEN_4[13:5] ? valid_223 : _GEN_2841; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2843 = 9'he0 == _GEN_4[13:5] ? valid_224 : _GEN_2842; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2844 = 9'he1 == _GEN_4[13:5] ? valid_225 : _GEN_2843; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2845 = 9'he2 == _GEN_4[13:5] ? valid_226 : _GEN_2844; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2846 = 9'he3 == _GEN_4[13:5] ? valid_227 : _GEN_2845; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2847 = 9'he4 == _GEN_4[13:5] ? valid_228 : _GEN_2846; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2848 = 9'he5 == _GEN_4[13:5] ? valid_229 : _GEN_2847; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2849 = 9'he6 == _GEN_4[13:5] ? valid_230 : _GEN_2848; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2850 = 9'he7 == _GEN_4[13:5] ? valid_231 : _GEN_2849; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2851 = 9'he8 == _GEN_4[13:5] ? valid_232 : _GEN_2850; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2852 = 9'he9 == _GEN_4[13:5] ? valid_233 : _GEN_2851; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2853 = 9'hea == _GEN_4[13:5] ? valid_234 : _GEN_2852; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2854 = 9'heb == _GEN_4[13:5] ? valid_235 : _GEN_2853; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2855 = 9'hec == _GEN_4[13:5] ? valid_236 : _GEN_2854; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2856 = 9'hed == _GEN_4[13:5] ? valid_237 : _GEN_2855; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2857 = 9'hee == _GEN_4[13:5] ? valid_238 : _GEN_2856; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2858 = 9'hef == _GEN_4[13:5] ? valid_239 : _GEN_2857; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2859 = 9'hf0 == _GEN_4[13:5] ? valid_240 : _GEN_2858; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2860 = 9'hf1 == _GEN_4[13:5] ? valid_241 : _GEN_2859; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2861 = 9'hf2 == _GEN_4[13:5] ? valid_242 : _GEN_2860; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2862 = 9'hf3 == _GEN_4[13:5] ? valid_243 : _GEN_2861; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2863 = 9'hf4 == _GEN_4[13:5] ? valid_244 : _GEN_2862; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2864 = 9'hf5 == _GEN_4[13:5] ? valid_245 : _GEN_2863; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2865 = 9'hf6 == _GEN_4[13:5] ? valid_246 : _GEN_2864; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2866 = 9'hf7 == _GEN_4[13:5] ? valid_247 : _GEN_2865; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2867 = 9'hf8 == _GEN_4[13:5] ? valid_248 : _GEN_2866; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2868 = 9'hf9 == _GEN_4[13:5] ? valid_249 : _GEN_2867; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2869 = 9'hfa == _GEN_4[13:5] ? valid_250 : _GEN_2868; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2870 = 9'hfb == _GEN_4[13:5] ? valid_251 : _GEN_2869; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2871 = 9'hfc == _GEN_4[13:5] ? valid_252 : _GEN_2870; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2872 = 9'hfd == _GEN_4[13:5] ? valid_253 : _GEN_2871; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2873 = 9'hfe == _GEN_4[13:5] ? valid_254 : _GEN_2872; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2874 = 9'hff == _GEN_4[13:5] ? valid_255 : _GEN_2873; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2875 = 9'h100 == _GEN_4[13:5] ? valid_256 : _GEN_2874; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2876 = 9'h101 == _GEN_4[13:5] ? valid_257 : _GEN_2875; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2877 = 9'h102 == _GEN_4[13:5] ? valid_258 : _GEN_2876; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2878 = 9'h103 == _GEN_4[13:5] ? valid_259 : _GEN_2877; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2879 = 9'h104 == _GEN_4[13:5] ? valid_260 : _GEN_2878; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2880 = 9'h105 == _GEN_4[13:5] ? valid_261 : _GEN_2879; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2881 = 9'h106 == _GEN_4[13:5] ? valid_262 : _GEN_2880; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2882 = 9'h107 == _GEN_4[13:5] ? valid_263 : _GEN_2881; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2883 = 9'h108 == _GEN_4[13:5] ? valid_264 : _GEN_2882; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2884 = 9'h109 == _GEN_4[13:5] ? valid_265 : _GEN_2883; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2885 = 9'h10a == _GEN_4[13:5] ? valid_266 : _GEN_2884; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2886 = 9'h10b == _GEN_4[13:5] ? valid_267 : _GEN_2885; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2887 = 9'h10c == _GEN_4[13:5] ? valid_268 : _GEN_2886; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2888 = 9'h10d == _GEN_4[13:5] ? valid_269 : _GEN_2887; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2889 = 9'h10e == _GEN_4[13:5] ? valid_270 : _GEN_2888; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2890 = 9'h10f == _GEN_4[13:5] ? valid_271 : _GEN_2889; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2891 = 9'h110 == _GEN_4[13:5] ? valid_272 : _GEN_2890; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2892 = 9'h111 == _GEN_4[13:5] ? valid_273 : _GEN_2891; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2893 = 9'h112 == _GEN_4[13:5] ? valid_274 : _GEN_2892; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2894 = 9'h113 == _GEN_4[13:5] ? valid_275 : _GEN_2893; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2895 = 9'h114 == _GEN_4[13:5] ? valid_276 : _GEN_2894; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2896 = 9'h115 == _GEN_4[13:5] ? valid_277 : _GEN_2895; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2897 = 9'h116 == _GEN_4[13:5] ? valid_278 : _GEN_2896; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2898 = 9'h117 == _GEN_4[13:5] ? valid_279 : _GEN_2897; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2899 = 9'h118 == _GEN_4[13:5] ? valid_280 : _GEN_2898; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2900 = 9'h119 == _GEN_4[13:5] ? valid_281 : _GEN_2899; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2901 = 9'h11a == _GEN_4[13:5] ? valid_282 : _GEN_2900; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2902 = 9'h11b == _GEN_4[13:5] ? valid_283 : _GEN_2901; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2903 = 9'h11c == _GEN_4[13:5] ? valid_284 : _GEN_2902; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2904 = 9'h11d == _GEN_4[13:5] ? valid_285 : _GEN_2903; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2905 = 9'h11e == _GEN_4[13:5] ? valid_286 : _GEN_2904; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2906 = 9'h11f == _GEN_4[13:5] ? valid_287 : _GEN_2905; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2907 = 9'h120 == _GEN_4[13:5] ? valid_288 : _GEN_2906; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2908 = 9'h121 == _GEN_4[13:5] ? valid_289 : _GEN_2907; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2909 = 9'h122 == _GEN_4[13:5] ? valid_290 : _GEN_2908; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2910 = 9'h123 == _GEN_4[13:5] ? valid_291 : _GEN_2909; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2911 = 9'h124 == _GEN_4[13:5] ? valid_292 : _GEN_2910; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2912 = 9'h125 == _GEN_4[13:5] ? valid_293 : _GEN_2911; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2913 = 9'h126 == _GEN_4[13:5] ? valid_294 : _GEN_2912; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2914 = 9'h127 == _GEN_4[13:5] ? valid_295 : _GEN_2913; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2915 = 9'h128 == _GEN_4[13:5] ? valid_296 : _GEN_2914; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2916 = 9'h129 == _GEN_4[13:5] ? valid_297 : _GEN_2915; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2917 = 9'h12a == _GEN_4[13:5] ? valid_298 : _GEN_2916; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2918 = 9'h12b == _GEN_4[13:5] ? valid_299 : _GEN_2917; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2919 = 9'h12c == _GEN_4[13:5] ? valid_300 : _GEN_2918; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2920 = 9'h12d == _GEN_4[13:5] ? valid_301 : _GEN_2919; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2921 = 9'h12e == _GEN_4[13:5] ? valid_302 : _GEN_2920; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2922 = 9'h12f == _GEN_4[13:5] ? valid_303 : _GEN_2921; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2923 = 9'h130 == _GEN_4[13:5] ? valid_304 : _GEN_2922; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2924 = 9'h131 == _GEN_4[13:5] ? valid_305 : _GEN_2923; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2925 = 9'h132 == _GEN_4[13:5] ? valid_306 : _GEN_2924; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2926 = 9'h133 == _GEN_4[13:5] ? valid_307 : _GEN_2925; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2927 = 9'h134 == _GEN_4[13:5] ? valid_308 : _GEN_2926; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2928 = 9'h135 == _GEN_4[13:5] ? valid_309 : _GEN_2927; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2929 = 9'h136 == _GEN_4[13:5] ? valid_310 : _GEN_2928; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2930 = 9'h137 == _GEN_4[13:5] ? valid_311 : _GEN_2929; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2931 = 9'h138 == _GEN_4[13:5] ? valid_312 : _GEN_2930; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2932 = 9'h139 == _GEN_4[13:5] ? valid_313 : _GEN_2931; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2933 = 9'h13a == _GEN_4[13:5] ? valid_314 : _GEN_2932; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2934 = 9'h13b == _GEN_4[13:5] ? valid_315 : _GEN_2933; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2935 = 9'h13c == _GEN_4[13:5] ? valid_316 : _GEN_2934; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2936 = 9'h13d == _GEN_4[13:5] ? valid_317 : _GEN_2935; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2937 = 9'h13e == _GEN_4[13:5] ? valid_318 : _GEN_2936; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2938 = 9'h13f == _GEN_4[13:5] ? valid_319 : _GEN_2937; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2939 = 9'h140 == _GEN_4[13:5] ? valid_320 : _GEN_2938; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2940 = 9'h141 == _GEN_4[13:5] ? valid_321 : _GEN_2939; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2941 = 9'h142 == _GEN_4[13:5] ? valid_322 : _GEN_2940; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2942 = 9'h143 == _GEN_4[13:5] ? valid_323 : _GEN_2941; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2943 = 9'h144 == _GEN_4[13:5] ? valid_324 : _GEN_2942; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2944 = 9'h145 == _GEN_4[13:5] ? valid_325 : _GEN_2943; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2945 = 9'h146 == _GEN_4[13:5] ? valid_326 : _GEN_2944; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2946 = 9'h147 == _GEN_4[13:5] ? valid_327 : _GEN_2945; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2947 = 9'h148 == _GEN_4[13:5] ? valid_328 : _GEN_2946; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2948 = 9'h149 == _GEN_4[13:5] ? valid_329 : _GEN_2947; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2949 = 9'h14a == _GEN_4[13:5] ? valid_330 : _GEN_2948; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2950 = 9'h14b == _GEN_4[13:5] ? valid_331 : _GEN_2949; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2951 = 9'h14c == _GEN_4[13:5] ? valid_332 : _GEN_2950; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2952 = 9'h14d == _GEN_4[13:5] ? valid_333 : _GEN_2951; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2953 = 9'h14e == _GEN_4[13:5] ? valid_334 : _GEN_2952; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2954 = 9'h14f == _GEN_4[13:5] ? valid_335 : _GEN_2953; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2955 = 9'h150 == _GEN_4[13:5] ? valid_336 : _GEN_2954; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2956 = 9'h151 == _GEN_4[13:5] ? valid_337 : _GEN_2955; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2957 = 9'h152 == _GEN_4[13:5] ? valid_338 : _GEN_2956; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2958 = 9'h153 == _GEN_4[13:5] ? valid_339 : _GEN_2957; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2959 = 9'h154 == _GEN_4[13:5] ? valid_340 : _GEN_2958; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2960 = 9'h155 == _GEN_4[13:5] ? valid_341 : _GEN_2959; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2961 = 9'h156 == _GEN_4[13:5] ? valid_342 : _GEN_2960; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2962 = 9'h157 == _GEN_4[13:5] ? valid_343 : _GEN_2961; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2963 = 9'h158 == _GEN_4[13:5] ? valid_344 : _GEN_2962; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2964 = 9'h159 == _GEN_4[13:5] ? valid_345 : _GEN_2963; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2965 = 9'h15a == _GEN_4[13:5] ? valid_346 : _GEN_2964; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2966 = 9'h15b == _GEN_4[13:5] ? valid_347 : _GEN_2965; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2967 = 9'h15c == _GEN_4[13:5] ? valid_348 : _GEN_2966; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2968 = 9'h15d == _GEN_4[13:5] ? valid_349 : _GEN_2967; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2969 = 9'h15e == _GEN_4[13:5] ? valid_350 : _GEN_2968; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2970 = 9'h15f == _GEN_4[13:5] ? valid_351 : _GEN_2969; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2971 = 9'h160 == _GEN_4[13:5] ? valid_352 : _GEN_2970; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2972 = 9'h161 == _GEN_4[13:5] ? valid_353 : _GEN_2971; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2973 = 9'h162 == _GEN_4[13:5] ? valid_354 : _GEN_2972; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2974 = 9'h163 == _GEN_4[13:5] ? valid_355 : _GEN_2973; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2975 = 9'h164 == _GEN_4[13:5] ? valid_356 : _GEN_2974; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2976 = 9'h165 == _GEN_4[13:5] ? valid_357 : _GEN_2975; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2977 = 9'h166 == _GEN_4[13:5] ? valid_358 : _GEN_2976; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2978 = 9'h167 == _GEN_4[13:5] ? valid_359 : _GEN_2977; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2979 = 9'h168 == _GEN_4[13:5] ? valid_360 : _GEN_2978; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2980 = 9'h169 == _GEN_4[13:5] ? valid_361 : _GEN_2979; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2981 = 9'h16a == _GEN_4[13:5] ? valid_362 : _GEN_2980; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2982 = 9'h16b == _GEN_4[13:5] ? valid_363 : _GEN_2981; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2983 = 9'h16c == _GEN_4[13:5] ? valid_364 : _GEN_2982; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2984 = 9'h16d == _GEN_4[13:5] ? valid_365 : _GEN_2983; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2985 = 9'h16e == _GEN_4[13:5] ? valid_366 : _GEN_2984; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2986 = 9'h16f == _GEN_4[13:5] ? valid_367 : _GEN_2985; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2987 = 9'h170 == _GEN_4[13:5] ? valid_368 : _GEN_2986; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2988 = 9'h171 == _GEN_4[13:5] ? valid_369 : _GEN_2987; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2989 = 9'h172 == _GEN_4[13:5] ? valid_370 : _GEN_2988; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2990 = 9'h173 == _GEN_4[13:5] ? valid_371 : _GEN_2989; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2991 = 9'h174 == _GEN_4[13:5] ? valid_372 : _GEN_2990; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2992 = 9'h175 == _GEN_4[13:5] ? valid_373 : _GEN_2991; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2993 = 9'h176 == _GEN_4[13:5] ? valid_374 : _GEN_2992; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2994 = 9'h177 == _GEN_4[13:5] ? valid_375 : _GEN_2993; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2995 = 9'h178 == _GEN_4[13:5] ? valid_376 : _GEN_2994; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2996 = 9'h179 == _GEN_4[13:5] ? valid_377 : _GEN_2995; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2997 = 9'h17a == _GEN_4[13:5] ? valid_378 : _GEN_2996; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2998 = 9'h17b == _GEN_4[13:5] ? valid_379 : _GEN_2997; // @[DCache.scala 234:{48,48}]
  wire  _GEN_2999 = 9'h17c == _GEN_4[13:5] ? valid_380 : _GEN_2998; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3000 = 9'h17d == _GEN_4[13:5] ? valid_381 : _GEN_2999; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3001 = 9'h17e == _GEN_4[13:5] ? valid_382 : _GEN_3000; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3002 = 9'h17f == _GEN_4[13:5] ? valid_383 : _GEN_3001; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3003 = 9'h180 == _GEN_4[13:5] ? valid_384 : _GEN_3002; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3004 = 9'h181 == _GEN_4[13:5] ? valid_385 : _GEN_3003; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3005 = 9'h182 == _GEN_4[13:5] ? valid_386 : _GEN_3004; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3006 = 9'h183 == _GEN_4[13:5] ? valid_387 : _GEN_3005; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3007 = 9'h184 == _GEN_4[13:5] ? valid_388 : _GEN_3006; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3008 = 9'h185 == _GEN_4[13:5] ? valid_389 : _GEN_3007; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3009 = 9'h186 == _GEN_4[13:5] ? valid_390 : _GEN_3008; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3010 = 9'h187 == _GEN_4[13:5] ? valid_391 : _GEN_3009; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3011 = 9'h188 == _GEN_4[13:5] ? valid_392 : _GEN_3010; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3012 = 9'h189 == _GEN_4[13:5] ? valid_393 : _GEN_3011; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3013 = 9'h18a == _GEN_4[13:5] ? valid_394 : _GEN_3012; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3014 = 9'h18b == _GEN_4[13:5] ? valid_395 : _GEN_3013; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3015 = 9'h18c == _GEN_4[13:5] ? valid_396 : _GEN_3014; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3016 = 9'h18d == _GEN_4[13:5] ? valid_397 : _GEN_3015; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3017 = 9'h18e == _GEN_4[13:5] ? valid_398 : _GEN_3016; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3018 = 9'h18f == _GEN_4[13:5] ? valid_399 : _GEN_3017; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3019 = 9'h190 == _GEN_4[13:5] ? valid_400 : _GEN_3018; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3020 = 9'h191 == _GEN_4[13:5] ? valid_401 : _GEN_3019; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3021 = 9'h192 == _GEN_4[13:5] ? valid_402 : _GEN_3020; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3022 = 9'h193 == _GEN_4[13:5] ? valid_403 : _GEN_3021; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3023 = 9'h194 == _GEN_4[13:5] ? valid_404 : _GEN_3022; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3024 = 9'h195 == _GEN_4[13:5] ? valid_405 : _GEN_3023; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3025 = 9'h196 == _GEN_4[13:5] ? valid_406 : _GEN_3024; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3026 = 9'h197 == _GEN_4[13:5] ? valid_407 : _GEN_3025; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3027 = 9'h198 == _GEN_4[13:5] ? valid_408 : _GEN_3026; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3028 = 9'h199 == _GEN_4[13:5] ? valid_409 : _GEN_3027; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3029 = 9'h19a == _GEN_4[13:5] ? valid_410 : _GEN_3028; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3030 = 9'h19b == _GEN_4[13:5] ? valid_411 : _GEN_3029; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3031 = 9'h19c == _GEN_4[13:5] ? valid_412 : _GEN_3030; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3032 = 9'h19d == _GEN_4[13:5] ? valid_413 : _GEN_3031; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3033 = 9'h19e == _GEN_4[13:5] ? valid_414 : _GEN_3032; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3034 = 9'h19f == _GEN_4[13:5] ? valid_415 : _GEN_3033; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3035 = 9'h1a0 == _GEN_4[13:5] ? valid_416 : _GEN_3034; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3036 = 9'h1a1 == _GEN_4[13:5] ? valid_417 : _GEN_3035; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3037 = 9'h1a2 == _GEN_4[13:5] ? valid_418 : _GEN_3036; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3038 = 9'h1a3 == _GEN_4[13:5] ? valid_419 : _GEN_3037; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3039 = 9'h1a4 == _GEN_4[13:5] ? valid_420 : _GEN_3038; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3040 = 9'h1a5 == _GEN_4[13:5] ? valid_421 : _GEN_3039; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3041 = 9'h1a6 == _GEN_4[13:5] ? valid_422 : _GEN_3040; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3042 = 9'h1a7 == _GEN_4[13:5] ? valid_423 : _GEN_3041; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3043 = 9'h1a8 == _GEN_4[13:5] ? valid_424 : _GEN_3042; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3044 = 9'h1a9 == _GEN_4[13:5] ? valid_425 : _GEN_3043; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3045 = 9'h1aa == _GEN_4[13:5] ? valid_426 : _GEN_3044; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3046 = 9'h1ab == _GEN_4[13:5] ? valid_427 : _GEN_3045; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3047 = 9'h1ac == _GEN_4[13:5] ? valid_428 : _GEN_3046; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3048 = 9'h1ad == _GEN_4[13:5] ? valid_429 : _GEN_3047; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3049 = 9'h1ae == _GEN_4[13:5] ? valid_430 : _GEN_3048; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3050 = 9'h1af == _GEN_4[13:5] ? valid_431 : _GEN_3049; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3051 = 9'h1b0 == _GEN_4[13:5] ? valid_432 : _GEN_3050; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3052 = 9'h1b1 == _GEN_4[13:5] ? valid_433 : _GEN_3051; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3053 = 9'h1b2 == _GEN_4[13:5] ? valid_434 : _GEN_3052; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3054 = 9'h1b3 == _GEN_4[13:5] ? valid_435 : _GEN_3053; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3055 = 9'h1b4 == _GEN_4[13:5] ? valid_436 : _GEN_3054; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3056 = 9'h1b5 == _GEN_4[13:5] ? valid_437 : _GEN_3055; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3057 = 9'h1b6 == _GEN_4[13:5] ? valid_438 : _GEN_3056; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3058 = 9'h1b7 == _GEN_4[13:5] ? valid_439 : _GEN_3057; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3059 = 9'h1b8 == _GEN_4[13:5] ? valid_440 : _GEN_3058; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3060 = 9'h1b9 == _GEN_4[13:5] ? valid_441 : _GEN_3059; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3061 = 9'h1ba == _GEN_4[13:5] ? valid_442 : _GEN_3060; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3062 = 9'h1bb == _GEN_4[13:5] ? valid_443 : _GEN_3061; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3063 = 9'h1bc == _GEN_4[13:5] ? valid_444 : _GEN_3062; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3064 = 9'h1bd == _GEN_4[13:5] ? valid_445 : _GEN_3063; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3065 = 9'h1be == _GEN_4[13:5] ? valid_446 : _GEN_3064; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3066 = 9'h1bf == _GEN_4[13:5] ? valid_447 : _GEN_3065; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3067 = 9'h1c0 == _GEN_4[13:5] ? valid_448 : _GEN_3066; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3068 = 9'h1c1 == _GEN_4[13:5] ? valid_449 : _GEN_3067; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3069 = 9'h1c2 == _GEN_4[13:5] ? valid_450 : _GEN_3068; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3070 = 9'h1c3 == _GEN_4[13:5] ? valid_451 : _GEN_3069; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3071 = 9'h1c4 == _GEN_4[13:5] ? valid_452 : _GEN_3070; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3072 = 9'h1c5 == _GEN_4[13:5] ? valid_453 : _GEN_3071; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3073 = 9'h1c6 == _GEN_4[13:5] ? valid_454 : _GEN_3072; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3074 = 9'h1c7 == _GEN_4[13:5] ? valid_455 : _GEN_3073; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3075 = 9'h1c8 == _GEN_4[13:5] ? valid_456 : _GEN_3074; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3076 = 9'h1c9 == _GEN_4[13:5] ? valid_457 : _GEN_3075; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3077 = 9'h1ca == _GEN_4[13:5] ? valid_458 : _GEN_3076; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3078 = 9'h1cb == _GEN_4[13:5] ? valid_459 : _GEN_3077; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3079 = 9'h1cc == _GEN_4[13:5] ? valid_460 : _GEN_3078; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3080 = 9'h1cd == _GEN_4[13:5] ? valid_461 : _GEN_3079; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3081 = 9'h1ce == _GEN_4[13:5] ? valid_462 : _GEN_3080; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3082 = 9'h1cf == _GEN_4[13:5] ? valid_463 : _GEN_3081; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3083 = 9'h1d0 == _GEN_4[13:5] ? valid_464 : _GEN_3082; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3084 = 9'h1d1 == _GEN_4[13:5] ? valid_465 : _GEN_3083; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3085 = 9'h1d2 == _GEN_4[13:5] ? valid_466 : _GEN_3084; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3086 = 9'h1d3 == _GEN_4[13:5] ? valid_467 : _GEN_3085; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3087 = 9'h1d4 == _GEN_4[13:5] ? valid_468 : _GEN_3086; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3088 = 9'h1d5 == _GEN_4[13:5] ? valid_469 : _GEN_3087; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3089 = 9'h1d6 == _GEN_4[13:5] ? valid_470 : _GEN_3088; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3090 = 9'h1d7 == _GEN_4[13:5] ? valid_471 : _GEN_3089; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3091 = 9'h1d8 == _GEN_4[13:5] ? valid_472 : _GEN_3090; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3092 = 9'h1d9 == _GEN_4[13:5] ? valid_473 : _GEN_3091; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3093 = 9'h1da == _GEN_4[13:5] ? valid_474 : _GEN_3092; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3094 = 9'h1db == _GEN_4[13:5] ? valid_475 : _GEN_3093; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3095 = 9'h1dc == _GEN_4[13:5] ? valid_476 : _GEN_3094; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3096 = 9'h1dd == _GEN_4[13:5] ? valid_477 : _GEN_3095; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3097 = 9'h1de == _GEN_4[13:5] ? valid_478 : _GEN_3096; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3098 = 9'h1df == _GEN_4[13:5] ? valid_479 : _GEN_3097; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3099 = 9'h1e0 == _GEN_4[13:5] ? valid_480 : _GEN_3098; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3100 = 9'h1e1 == _GEN_4[13:5] ? valid_481 : _GEN_3099; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3101 = 9'h1e2 == _GEN_4[13:5] ? valid_482 : _GEN_3100; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3102 = 9'h1e3 == _GEN_4[13:5] ? valid_483 : _GEN_3101; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3103 = 9'h1e4 == _GEN_4[13:5] ? valid_484 : _GEN_3102; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3104 = 9'h1e5 == _GEN_4[13:5] ? valid_485 : _GEN_3103; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3105 = 9'h1e6 == _GEN_4[13:5] ? valid_486 : _GEN_3104; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3106 = 9'h1e7 == _GEN_4[13:5] ? valid_487 : _GEN_3105; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3107 = 9'h1e8 == _GEN_4[13:5] ? valid_488 : _GEN_3106; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3108 = 9'h1e9 == _GEN_4[13:5] ? valid_489 : _GEN_3107; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3109 = 9'h1ea == _GEN_4[13:5] ? valid_490 : _GEN_3108; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3110 = 9'h1eb == _GEN_4[13:5] ? valid_491 : _GEN_3109; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3111 = 9'h1ec == _GEN_4[13:5] ? valid_492 : _GEN_3110; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3112 = 9'h1ed == _GEN_4[13:5] ? valid_493 : _GEN_3111; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3113 = 9'h1ee == _GEN_4[13:5] ? valid_494 : _GEN_3112; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3114 = 9'h1ef == _GEN_4[13:5] ? valid_495 : _GEN_3113; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3115 = 9'h1f0 == _GEN_4[13:5] ? valid_496 : _GEN_3114; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3116 = 9'h1f1 == _GEN_4[13:5] ? valid_497 : _GEN_3115; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3117 = 9'h1f2 == _GEN_4[13:5] ? valid_498 : _GEN_3116; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3118 = 9'h1f3 == _GEN_4[13:5] ? valid_499 : _GEN_3117; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3119 = 9'h1f4 == _GEN_4[13:5] ? valid_500 : _GEN_3118; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3120 = 9'h1f5 == _GEN_4[13:5] ? valid_501 : _GEN_3119; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3121 = 9'h1f6 == _GEN_4[13:5] ? valid_502 : _GEN_3120; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3122 = 9'h1f7 == _GEN_4[13:5] ? valid_503 : _GEN_3121; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3123 = 9'h1f8 == _GEN_4[13:5] ? valid_504 : _GEN_3122; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3124 = 9'h1f9 == _GEN_4[13:5] ? valid_505 : _GEN_3123; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3125 = 9'h1fa == _GEN_4[13:5] ? valid_506 : _GEN_3124; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3126 = 9'h1fb == _GEN_4[13:5] ? valid_507 : _GEN_3125; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3127 = 9'h1fc == _GEN_4[13:5] ? valid_508 : _GEN_3126; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3128 = 9'h1fd == _GEN_4[13:5] ? valid_509 : _GEN_3127; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3129 = 9'h1fe == _GEN_4[13:5] ? valid_510 : _GEN_3128; // @[DCache.scala 234:{48,48}]
  wire  _GEN_3130 = 9'h1ff == _GEN_4[13:5] ? valid_511 : _GEN_3129; // @[DCache.scala 234:{48,48}]
  wire  probe_hit = _GEN_3130 & _GEN_4[31:14] == probe_out_tag; // @[DCache.scala 234:48]
  reg [8:0] release_addr_aligned_REG; // @[DCache.scala 245:56]
  wire [31:0] release_addr_aligned = {array_out_tag,release_addr_aligned_REG,5'h0}; // @[Cat.scala 33:92]
  wire  _source_T_2 = _T_27 | _probing_T_1; // @[DCache.scala 249:47]
  reg [1:0] source; // @[Counter.scala 61:40]
  wire [1:0] _source_wrap_value_T_1 = source + 2'h1; // @[Counter.scala 77:24]
  wire [2:0] _x1_c_bits_T_opcode = probe_hit ? 3'h5 : 3'h4; // @[DCache.scala 259:33]
  wire [2:0] _x1_c_bits_T_param = probe_hit ? 3'h1 : 3'h5; // @[DCache.scala 259:33]
  wire [255:0] _x1_c_bits_T_data = probe_hit ? probe_out_data : 256'h0; // @[DCache.scala 259:33]
  wire  _io_cache_req_ready_T_3 = ~(probing | _tl_b_bits_r_T); // @[DCache.scala 266:44]
  SRAM array ( // @[DCache.scala 55:21]
    .clock(array_clock),
    .io_en(array_io_en),
    .io_addr(array_io_addr),
    .io_wdata(array_io_wdata),
    .io_wen(array_io_wen),
    .io_rdata(array_io_rdata)
  );
  assign auto_out_a_valid = state == 3'h4; // @[DCache.scala 257:24]
  assign auto_out_a_bits_source = source; // @[Edges.scala 345:17 349:15]
  assign auto_out_a_bits_address = {req_r_addr[31:5],5'h0}; // @[Cat.scala 33:92]
  assign auto_out_b_ready = ~probing & (~lrsc_reserved | lrsc_backoff); // @[DCache.scala 258:26]
  assign auto_out_c_valid = probing | state == 3'h2 & _GEN_535; // @[DCache.scala 260:25]
  assign auto_out_c_bits_opcode = probing ? _x1_c_bits_T_opcode : 3'h7; // @[DCache.scala 259:20]
  assign auto_out_c_bits_param = probing ? _x1_c_bits_T_param : 3'h1; // @[DCache.scala 259:20]
  assign auto_out_c_bits_size = probing ? tl_b_bits_r_size : 3'h5; // @[DCache.scala 259:20]
  assign auto_out_c_bits_source = probing ? tl_b_bits_r_source : source; // @[DCache.scala 259:20]
  assign auto_out_c_bits_address = probing ? tl_b_bits_r_address : release_addr_aligned; // @[DCache.scala 259:20]
  assign auto_out_c_bits_data = probing ? _x1_c_bits_T_data : array_out_data; // @[DCache.scala 259:20]
  assign auto_out_d_ready = state == 3'h3 | state == 3'h5; // @[DCache.scala 261:43]
  assign auto_out_e_valid = state == 3'h6; // @[DCache.scala 263:24]
  assign auto_out_e_bits_sink = tl_d_bits_r_sink; // @[Edges.scala 438:17 439:12]
  assign io_cache_req_ready = state == 3'h0 & ~(probing | _tl_b_bits_r_T); // @[DCache.scala 266:41]
  assign io_cache_resp_valid = (state == 3'h1 & array_hit | _T_11) & _io_cache_req_ready_T_3; // @[DCache.scala 267:77]
  assign io_cache_resp_bits_rdata = is_sc_r ? sc_rdata_64 : rdata_64; // @[DCache.scala 269:25]
  assign array_clock = clock;
  assign array_io_en = _req_r_T | _array_io_en_T_1 | _tl_b_bits_r_T; // @[DCache.scala 70:45]
  assign array_io_addr = _tl_b_bits_r_T ? _GEN_4[13:5] : array_addr[13:5]; // @[DCache.scala 235:19 236:19 71:20]
  assign array_io_wdata = {array_wdata_tag,array_wdata_data}; // @[DCache.scala 72:35]
  assign array_io_wen = _array_io_en_T_1 & _GEN_1571; // @[DCache.scala 164:19 73:20]
  always @(posedge clock) begin
    if (reset) begin // @[Utils.scala 36:20]
      probing <= 1'h0; // @[Utils.scala 36:20]
    end else begin
      probing <= _GEN_2599;
    end
    if (reset) begin // @[DCache.scala 127:30]
      lrsc_reserved <= 1'h0; // @[DCache.scala 127:30]
    end else if (_array_io_en_T_1 & req_r_wen) begin // @[DCache.scala 147:32]
      lrsc_reserved <= 1'h0; // @[DCache.scala 148:19]
    end else if (_tl_b_bits_r_T & auto_out_b_bits_address[31:5] == lrsc_addr) begin // @[DCache.scala 139:73]
      lrsc_reserved <= 1'h0; // @[DCache.scala 140:19]
    end else begin
      lrsc_reserved <= _GEN_536;
    end
    if (reset) begin // @[DCache.scala 129:30]
      lrsc_counter <= 5'h0; // @[DCache.scala 129:30]
    end else if (_array_io_en_T_1 & req_r_wen) begin // @[DCache.scala 147:32]
      lrsc_counter <= 5'h0; // @[DCache.scala 149:19]
    end else if (_tl_b_bits_r_T & auto_out_b_bits_address[31:5] == lrsc_addr) begin // @[DCache.scala 139:73]
      lrsc_counter <= 5'h0; // @[DCache.scala 141:19]
    end else if (lrsc_reserved & ~lrsc_backoff) begin // @[DCache.scala 136:40]
      lrsc_counter <= _lrsc_counter_T_1; // @[DCache.scala 137:18]
    end
    if (reset) begin // @[Reg.scala 35:20]
      tl_b_bits_r_size <= 3'h0; // @[Reg.scala 35:20]
    end else if (_tl_b_bits_r_T) begin // @[Reg.scala 36:18]
      tl_b_bits_r_size <= auto_out_b_bits_size; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      tl_b_bits_r_source <= 2'h0; // @[Reg.scala 35:20]
    end else if (_tl_b_bits_r_T) begin // @[Reg.scala 36:18]
      tl_b_bits_r_source <= auto_out_b_bits_source; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      tl_b_bits_r_address <= 32'h0; // @[Reg.scala 35:20]
    end else if (_tl_b_bits_r_T) begin // @[Reg.scala 36:18]
      tl_b_bits_r_address <= auto_out_b_bits_address; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[DCache.scala 60:118]
      state <= 3'h0; // @[DCache.scala 60:118]
    end else if (3'h0 == state) begin // @[DCache.scala 184:17]
      if (_req_r_T) begin // @[DCache.scala 186:22]
        if (sc_fail) begin // @[DCache.scala 187:21]
          state <= 3'h7;
        end else begin
          state <= 3'h1;
        end
      end
    end else if (3'h1 == state) begin // @[DCache.scala 184:17]
      if (_array_io_en_T_1) begin // @[DCache.scala 191:23]
        state <= 3'h0; // @[DCache.scala 192:15]
      end else begin
        state <= _GEN_2601;
      end
    end else if (3'h2 == state) begin // @[DCache.scala 184:17]
      state <= _GEN_2604;
    end else begin
      state <= _GEN_2614;
    end
    if (reset) begin // @[Reg.scala 35:20]
      tl_d_bits_r_sink <= 6'h0; // @[Reg.scala 35:20]
    end else if (_tl_d_bits_r_T) begin // @[Reg.scala 36:18]
      tl_d_bits_r_sink <= auto_out_d_bits_sink; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      tl_d_bits_r_data <= 256'h0; // @[Reg.scala 35:20]
    end else if (_tl_d_bits_r_T) begin // @[Reg.scala 36:18]
      tl_d_bits_r_data <= auto_out_d_bits_data; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      req_r_addr <= 39'h0; // @[Reg.scala 35:20]
    end else if (_req_r_T) begin // @[Reg.scala 36:18]
      req_r_addr <= io_cache_req_bits_addr; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      req_r_wdata <= 64'h0; // @[Reg.scala 35:20]
    end else if (_req_r_T) begin // @[Reg.scala 36:18]
      req_r_wdata <= io_cache_req_bits_wdata; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      req_r_wmask <= 8'h0; // @[Reg.scala 35:20]
    end else if (_req_r_T) begin // @[Reg.scala 36:18]
      req_r_wmask <= io_cache_req_bits_wmask; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      req_r_wen <= 1'h0; // @[Reg.scala 35:20]
    end else if (_req_r_T) begin // @[Reg.scala 36:18]
      req_r_wen <= io_cache_req_bits_wen; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      req_r_len <= 2'h0; // @[Reg.scala 35:20]
    end else if (_req_r_T) begin // @[Reg.scala 36:18]
      req_r_len <= io_cache_req_bits_len; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      req_r_lrsc <= 1'h0; // @[Reg.scala 35:20]
    end else if (_req_r_T) begin // @[Reg.scala 36:18]
      req_r_lrsc <= io_cache_req_bits_lrsc; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      req_r_amo <= 5'h0; // @[Reg.scala 35:20]
    end else if (_req_r_T) begin // @[Reg.scala 36:18]
      req_r_amo <= io_cache_req_bits_amo; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_0 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h0 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_0 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_0 <= _GEN_2086;
      end
    end else begin
      valid_0 <= _GEN_2086;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_1 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_1 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_1 <= _GEN_2087;
      end
    end else begin
      valid_1 <= _GEN_2087;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_2 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h2 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_2 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_2 <= _GEN_2088;
      end
    end else begin
      valid_2 <= _GEN_2088;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_3 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h3 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_3 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_3 <= _GEN_2089;
      end
    end else begin
      valid_3 <= _GEN_2089;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_4 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h4 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_4 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_4 <= _GEN_2090;
      end
    end else begin
      valid_4 <= _GEN_2090;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_5 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h5 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_5 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_5 <= _GEN_2091;
      end
    end else begin
      valid_5 <= _GEN_2091;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_6 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h6 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_6 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_6 <= _GEN_2092;
      end
    end else begin
      valid_6 <= _GEN_2092;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_7 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h7 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_7 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_7 <= _GEN_2093;
      end
    end else begin
      valid_7 <= _GEN_2093;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_8 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h8 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_8 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_8 <= _GEN_2094;
      end
    end else begin
      valid_8 <= _GEN_2094;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_9 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h9 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_9 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_9 <= _GEN_2095;
      end
    end else begin
      valid_9 <= _GEN_2095;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_10 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'ha == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_10 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_10 <= _GEN_2096;
      end
    end else begin
      valid_10 <= _GEN_2096;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_11 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hb == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_11 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_11 <= _GEN_2097;
      end
    end else begin
      valid_11 <= _GEN_2097;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_12 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hc == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_12 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_12 <= _GEN_2098;
      end
    end else begin
      valid_12 <= _GEN_2098;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_13 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hd == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_13 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_13 <= _GEN_2099;
      end
    end else begin
      valid_13 <= _GEN_2099;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_14 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'he == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_14 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_14 <= _GEN_2100;
      end
    end else begin
      valid_14 <= _GEN_2100;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_15 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hf == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_15 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_15 <= _GEN_2101;
      end
    end else begin
      valid_15 <= _GEN_2101;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_16 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h10 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_16 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_16 <= _GEN_2102;
      end
    end else begin
      valid_16 <= _GEN_2102;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_17 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h11 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_17 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_17 <= _GEN_2103;
      end
    end else begin
      valid_17 <= _GEN_2103;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_18 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h12 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_18 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_18 <= _GEN_2104;
      end
    end else begin
      valid_18 <= _GEN_2104;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_19 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h13 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_19 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_19 <= _GEN_2105;
      end
    end else begin
      valid_19 <= _GEN_2105;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_20 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h14 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_20 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_20 <= _GEN_2106;
      end
    end else begin
      valid_20 <= _GEN_2106;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_21 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h15 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_21 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_21 <= _GEN_2107;
      end
    end else begin
      valid_21 <= _GEN_2107;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_22 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h16 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_22 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_22 <= _GEN_2108;
      end
    end else begin
      valid_22 <= _GEN_2108;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_23 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h17 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_23 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_23 <= _GEN_2109;
      end
    end else begin
      valid_23 <= _GEN_2109;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_24 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h18 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_24 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_24 <= _GEN_2110;
      end
    end else begin
      valid_24 <= _GEN_2110;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_25 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h19 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_25 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_25 <= _GEN_2111;
      end
    end else begin
      valid_25 <= _GEN_2111;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_26 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1a == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_26 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_26 <= _GEN_2112;
      end
    end else begin
      valid_26 <= _GEN_2112;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_27 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1b == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_27 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_27 <= _GEN_2113;
      end
    end else begin
      valid_27 <= _GEN_2113;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_28 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1c == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_28 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_28 <= _GEN_2114;
      end
    end else begin
      valid_28 <= _GEN_2114;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_29 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1d == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_29 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_29 <= _GEN_2115;
      end
    end else begin
      valid_29 <= _GEN_2115;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_30 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1e == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_30 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_30 <= _GEN_2116;
      end
    end else begin
      valid_30 <= _GEN_2116;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_31 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1f == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_31 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_31 <= _GEN_2117;
      end
    end else begin
      valid_31 <= _GEN_2117;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_32 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h20 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_32 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_32 <= _GEN_2118;
      end
    end else begin
      valid_32 <= _GEN_2118;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_33 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h21 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_33 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_33 <= _GEN_2119;
      end
    end else begin
      valid_33 <= _GEN_2119;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_34 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h22 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_34 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_34 <= _GEN_2120;
      end
    end else begin
      valid_34 <= _GEN_2120;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_35 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h23 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_35 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_35 <= _GEN_2121;
      end
    end else begin
      valid_35 <= _GEN_2121;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_36 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h24 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_36 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_36 <= _GEN_2122;
      end
    end else begin
      valid_36 <= _GEN_2122;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_37 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h25 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_37 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_37 <= _GEN_2123;
      end
    end else begin
      valid_37 <= _GEN_2123;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_38 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h26 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_38 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_38 <= _GEN_2124;
      end
    end else begin
      valid_38 <= _GEN_2124;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_39 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h27 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_39 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_39 <= _GEN_2125;
      end
    end else begin
      valid_39 <= _GEN_2125;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_40 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h28 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_40 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_40 <= _GEN_2126;
      end
    end else begin
      valid_40 <= _GEN_2126;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_41 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h29 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_41 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_41 <= _GEN_2127;
      end
    end else begin
      valid_41 <= _GEN_2127;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_42 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h2a == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_42 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_42 <= _GEN_2128;
      end
    end else begin
      valid_42 <= _GEN_2128;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_43 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h2b == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_43 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_43 <= _GEN_2129;
      end
    end else begin
      valid_43 <= _GEN_2129;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_44 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h2c == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_44 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_44 <= _GEN_2130;
      end
    end else begin
      valid_44 <= _GEN_2130;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_45 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h2d == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_45 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_45 <= _GEN_2131;
      end
    end else begin
      valid_45 <= _GEN_2131;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_46 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h2e == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_46 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_46 <= _GEN_2132;
      end
    end else begin
      valid_46 <= _GEN_2132;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_47 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h2f == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_47 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_47 <= _GEN_2133;
      end
    end else begin
      valid_47 <= _GEN_2133;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_48 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h30 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_48 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_48 <= _GEN_2134;
      end
    end else begin
      valid_48 <= _GEN_2134;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_49 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h31 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_49 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_49 <= _GEN_2135;
      end
    end else begin
      valid_49 <= _GEN_2135;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_50 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h32 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_50 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_50 <= _GEN_2136;
      end
    end else begin
      valid_50 <= _GEN_2136;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_51 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h33 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_51 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_51 <= _GEN_2137;
      end
    end else begin
      valid_51 <= _GEN_2137;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_52 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h34 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_52 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_52 <= _GEN_2138;
      end
    end else begin
      valid_52 <= _GEN_2138;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_53 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h35 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_53 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_53 <= _GEN_2139;
      end
    end else begin
      valid_53 <= _GEN_2139;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_54 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h36 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_54 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_54 <= _GEN_2140;
      end
    end else begin
      valid_54 <= _GEN_2140;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_55 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h37 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_55 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_55 <= _GEN_2141;
      end
    end else begin
      valid_55 <= _GEN_2141;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_56 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h38 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_56 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_56 <= _GEN_2142;
      end
    end else begin
      valid_56 <= _GEN_2142;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_57 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h39 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_57 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_57 <= _GEN_2143;
      end
    end else begin
      valid_57 <= _GEN_2143;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_58 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h3a == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_58 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_58 <= _GEN_2144;
      end
    end else begin
      valid_58 <= _GEN_2144;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_59 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h3b == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_59 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_59 <= _GEN_2145;
      end
    end else begin
      valid_59 <= _GEN_2145;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_60 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h3c == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_60 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_60 <= _GEN_2146;
      end
    end else begin
      valid_60 <= _GEN_2146;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_61 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h3d == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_61 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_61 <= _GEN_2147;
      end
    end else begin
      valid_61 <= _GEN_2147;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_62 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h3e == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_62 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_62 <= _GEN_2148;
      end
    end else begin
      valid_62 <= _GEN_2148;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_63 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h3f == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_63 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_63 <= _GEN_2149;
      end
    end else begin
      valid_63 <= _GEN_2149;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_64 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h40 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_64 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_64 <= _GEN_2150;
      end
    end else begin
      valid_64 <= _GEN_2150;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_65 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h41 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_65 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_65 <= _GEN_2151;
      end
    end else begin
      valid_65 <= _GEN_2151;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_66 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h42 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_66 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_66 <= _GEN_2152;
      end
    end else begin
      valid_66 <= _GEN_2152;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_67 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h43 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_67 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_67 <= _GEN_2153;
      end
    end else begin
      valid_67 <= _GEN_2153;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_68 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h44 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_68 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_68 <= _GEN_2154;
      end
    end else begin
      valid_68 <= _GEN_2154;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_69 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h45 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_69 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_69 <= _GEN_2155;
      end
    end else begin
      valid_69 <= _GEN_2155;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_70 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h46 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_70 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_70 <= _GEN_2156;
      end
    end else begin
      valid_70 <= _GEN_2156;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_71 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h47 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_71 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_71 <= _GEN_2157;
      end
    end else begin
      valid_71 <= _GEN_2157;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_72 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h48 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_72 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_72 <= _GEN_2158;
      end
    end else begin
      valid_72 <= _GEN_2158;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_73 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h49 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_73 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_73 <= _GEN_2159;
      end
    end else begin
      valid_73 <= _GEN_2159;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_74 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h4a == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_74 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_74 <= _GEN_2160;
      end
    end else begin
      valid_74 <= _GEN_2160;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_75 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h4b == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_75 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_75 <= _GEN_2161;
      end
    end else begin
      valid_75 <= _GEN_2161;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_76 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h4c == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_76 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_76 <= _GEN_2162;
      end
    end else begin
      valid_76 <= _GEN_2162;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_77 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h4d == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_77 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_77 <= _GEN_2163;
      end
    end else begin
      valid_77 <= _GEN_2163;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_78 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h4e == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_78 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_78 <= _GEN_2164;
      end
    end else begin
      valid_78 <= _GEN_2164;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_79 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h4f == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_79 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_79 <= _GEN_2165;
      end
    end else begin
      valid_79 <= _GEN_2165;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_80 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h50 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_80 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_80 <= _GEN_2166;
      end
    end else begin
      valid_80 <= _GEN_2166;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_81 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h51 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_81 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_81 <= _GEN_2167;
      end
    end else begin
      valid_81 <= _GEN_2167;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_82 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h52 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_82 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_82 <= _GEN_2168;
      end
    end else begin
      valid_82 <= _GEN_2168;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_83 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h53 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_83 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_83 <= _GEN_2169;
      end
    end else begin
      valid_83 <= _GEN_2169;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_84 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h54 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_84 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_84 <= _GEN_2170;
      end
    end else begin
      valid_84 <= _GEN_2170;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_85 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h55 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_85 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_85 <= _GEN_2171;
      end
    end else begin
      valid_85 <= _GEN_2171;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_86 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h56 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_86 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_86 <= _GEN_2172;
      end
    end else begin
      valid_86 <= _GEN_2172;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_87 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h57 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_87 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_87 <= _GEN_2173;
      end
    end else begin
      valid_87 <= _GEN_2173;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_88 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h58 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_88 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_88 <= _GEN_2174;
      end
    end else begin
      valid_88 <= _GEN_2174;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_89 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h59 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_89 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_89 <= _GEN_2175;
      end
    end else begin
      valid_89 <= _GEN_2175;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_90 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h5a == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_90 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_90 <= _GEN_2176;
      end
    end else begin
      valid_90 <= _GEN_2176;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_91 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h5b == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_91 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_91 <= _GEN_2177;
      end
    end else begin
      valid_91 <= _GEN_2177;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_92 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h5c == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_92 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_92 <= _GEN_2178;
      end
    end else begin
      valid_92 <= _GEN_2178;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_93 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h5d == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_93 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_93 <= _GEN_2179;
      end
    end else begin
      valid_93 <= _GEN_2179;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_94 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h5e == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_94 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_94 <= _GEN_2180;
      end
    end else begin
      valid_94 <= _GEN_2180;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_95 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h5f == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_95 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_95 <= _GEN_2181;
      end
    end else begin
      valid_95 <= _GEN_2181;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_96 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h60 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_96 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_96 <= _GEN_2182;
      end
    end else begin
      valid_96 <= _GEN_2182;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_97 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h61 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_97 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_97 <= _GEN_2183;
      end
    end else begin
      valid_97 <= _GEN_2183;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_98 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h62 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_98 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_98 <= _GEN_2184;
      end
    end else begin
      valid_98 <= _GEN_2184;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_99 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h63 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_99 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_99 <= _GEN_2185;
      end
    end else begin
      valid_99 <= _GEN_2185;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_100 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h64 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_100 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_100 <= _GEN_2186;
      end
    end else begin
      valid_100 <= _GEN_2186;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_101 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h65 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_101 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_101 <= _GEN_2187;
      end
    end else begin
      valid_101 <= _GEN_2187;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_102 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h66 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_102 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_102 <= _GEN_2188;
      end
    end else begin
      valid_102 <= _GEN_2188;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_103 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h67 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_103 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_103 <= _GEN_2189;
      end
    end else begin
      valid_103 <= _GEN_2189;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_104 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h68 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_104 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_104 <= _GEN_2190;
      end
    end else begin
      valid_104 <= _GEN_2190;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_105 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h69 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_105 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_105 <= _GEN_2191;
      end
    end else begin
      valid_105 <= _GEN_2191;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_106 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h6a == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_106 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_106 <= _GEN_2192;
      end
    end else begin
      valid_106 <= _GEN_2192;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_107 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h6b == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_107 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_107 <= _GEN_2193;
      end
    end else begin
      valid_107 <= _GEN_2193;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_108 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h6c == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_108 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_108 <= _GEN_2194;
      end
    end else begin
      valid_108 <= _GEN_2194;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_109 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h6d == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_109 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_109 <= _GEN_2195;
      end
    end else begin
      valid_109 <= _GEN_2195;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_110 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h6e == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_110 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_110 <= _GEN_2196;
      end
    end else begin
      valid_110 <= _GEN_2196;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_111 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h6f == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_111 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_111 <= _GEN_2197;
      end
    end else begin
      valid_111 <= _GEN_2197;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_112 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h70 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_112 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_112 <= _GEN_2198;
      end
    end else begin
      valid_112 <= _GEN_2198;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_113 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h71 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_113 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_113 <= _GEN_2199;
      end
    end else begin
      valid_113 <= _GEN_2199;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_114 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h72 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_114 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_114 <= _GEN_2200;
      end
    end else begin
      valid_114 <= _GEN_2200;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_115 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h73 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_115 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_115 <= _GEN_2201;
      end
    end else begin
      valid_115 <= _GEN_2201;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_116 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h74 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_116 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_116 <= _GEN_2202;
      end
    end else begin
      valid_116 <= _GEN_2202;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_117 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h75 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_117 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_117 <= _GEN_2203;
      end
    end else begin
      valid_117 <= _GEN_2203;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_118 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h76 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_118 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_118 <= _GEN_2204;
      end
    end else begin
      valid_118 <= _GEN_2204;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_119 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h77 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_119 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_119 <= _GEN_2205;
      end
    end else begin
      valid_119 <= _GEN_2205;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_120 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h78 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_120 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_120 <= _GEN_2206;
      end
    end else begin
      valid_120 <= _GEN_2206;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_121 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h79 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_121 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_121 <= _GEN_2207;
      end
    end else begin
      valid_121 <= _GEN_2207;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_122 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h7a == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_122 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_122 <= _GEN_2208;
      end
    end else begin
      valid_122 <= _GEN_2208;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_123 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h7b == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_123 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_123 <= _GEN_2209;
      end
    end else begin
      valid_123 <= _GEN_2209;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_124 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h7c == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_124 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_124 <= _GEN_2210;
      end
    end else begin
      valid_124 <= _GEN_2210;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_125 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h7d == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_125 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_125 <= _GEN_2211;
      end
    end else begin
      valid_125 <= _GEN_2211;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_126 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h7e == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_126 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_126 <= _GEN_2212;
      end
    end else begin
      valid_126 <= _GEN_2212;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_127 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h7f == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_127 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_127 <= _GEN_2213;
      end
    end else begin
      valid_127 <= _GEN_2213;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_128 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h80 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_128 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_128 <= _GEN_2214;
      end
    end else begin
      valid_128 <= _GEN_2214;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_129 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h81 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_129 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_129 <= _GEN_2215;
      end
    end else begin
      valid_129 <= _GEN_2215;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_130 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h82 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_130 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_130 <= _GEN_2216;
      end
    end else begin
      valid_130 <= _GEN_2216;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_131 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h83 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_131 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_131 <= _GEN_2217;
      end
    end else begin
      valid_131 <= _GEN_2217;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_132 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h84 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_132 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_132 <= _GEN_2218;
      end
    end else begin
      valid_132 <= _GEN_2218;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_133 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h85 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_133 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_133 <= _GEN_2219;
      end
    end else begin
      valid_133 <= _GEN_2219;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_134 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h86 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_134 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_134 <= _GEN_2220;
      end
    end else begin
      valid_134 <= _GEN_2220;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_135 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h87 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_135 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_135 <= _GEN_2221;
      end
    end else begin
      valid_135 <= _GEN_2221;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_136 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h88 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_136 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_136 <= _GEN_2222;
      end
    end else begin
      valid_136 <= _GEN_2222;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_137 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h89 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_137 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_137 <= _GEN_2223;
      end
    end else begin
      valid_137 <= _GEN_2223;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_138 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h8a == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_138 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_138 <= _GEN_2224;
      end
    end else begin
      valid_138 <= _GEN_2224;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_139 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h8b == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_139 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_139 <= _GEN_2225;
      end
    end else begin
      valid_139 <= _GEN_2225;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_140 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h8c == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_140 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_140 <= _GEN_2226;
      end
    end else begin
      valid_140 <= _GEN_2226;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_141 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h8d == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_141 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_141 <= _GEN_2227;
      end
    end else begin
      valid_141 <= _GEN_2227;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_142 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h8e == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_142 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_142 <= _GEN_2228;
      end
    end else begin
      valid_142 <= _GEN_2228;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_143 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h8f == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_143 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_143 <= _GEN_2229;
      end
    end else begin
      valid_143 <= _GEN_2229;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_144 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h90 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_144 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_144 <= _GEN_2230;
      end
    end else begin
      valid_144 <= _GEN_2230;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_145 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h91 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_145 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_145 <= _GEN_2231;
      end
    end else begin
      valid_145 <= _GEN_2231;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_146 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h92 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_146 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_146 <= _GEN_2232;
      end
    end else begin
      valid_146 <= _GEN_2232;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_147 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h93 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_147 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_147 <= _GEN_2233;
      end
    end else begin
      valid_147 <= _GEN_2233;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_148 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h94 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_148 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_148 <= _GEN_2234;
      end
    end else begin
      valid_148 <= _GEN_2234;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_149 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h95 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_149 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_149 <= _GEN_2235;
      end
    end else begin
      valid_149 <= _GEN_2235;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_150 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h96 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_150 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_150 <= _GEN_2236;
      end
    end else begin
      valid_150 <= _GEN_2236;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_151 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h97 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_151 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_151 <= _GEN_2237;
      end
    end else begin
      valid_151 <= _GEN_2237;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_152 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h98 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_152 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_152 <= _GEN_2238;
      end
    end else begin
      valid_152 <= _GEN_2238;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_153 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h99 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_153 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_153 <= _GEN_2239;
      end
    end else begin
      valid_153 <= _GEN_2239;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_154 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h9a == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_154 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_154 <= _GEN_2240;
      end
    end else begin
      valid_154 <= _GEN_2240;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_155 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h9b == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_155 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_155 <= _GEN_2241;
      end
    end else begin
      valid_155 <= _GEN_2241;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_156 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h9c == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_156 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_156 <= _GEN_2242;
      end
    end else begin
      valid_156 <= _GEN_2242;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_157 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h9d == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_157 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_157 <= _GEN_2243;
      end
    end else begin
      valid_157 <= _GEN_2243;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_158 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h9e == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_158 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_158 <= _GEN_2244;
      end
    end else begin
      valid_158 <= _GEN_2244;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_159 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h9f == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_159 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_159 <= _GEN_2245;
      end
    end else begin
      valid_159 <= _GEN_2245;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_160 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'ha0 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_160 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_160 <= _GEN_2246;
      end
    end else begin
      valid_160 <= _GEN_2246;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_161 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'ha1 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_161 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_161 <= _GEN_2247;
      end
    end else begin
      valid_161 <= _GEN_2247;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_162 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'ha2 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_162 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_162 <= _GEN_2248;
      end
    end else begin
      valid_162 <= _GEN_2248;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_163 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'ha3 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_163 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_163 <= _GEN_2249;
      end
    end else begin
      valid_163 <= _GEN_2249;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_164 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'ha4 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_164 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_164 <= _GEN_2250;
      end
    end else begin
      valid_164 <= _GEN_2250;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_165 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'ha5 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_165 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_165 <= _GEN_2251;
      end
    end else begin
      valid_165 <= _GEN_2251;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_166 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'ha6 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_166 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_166 <= _GEN_2252;
      end
    end else begin
      valid_166 <= _GEN_2252;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_167 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'ha7 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_167 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_167 <= _GEN_2253;
      end
    end else begin
      valid_167 <= _GEN_2253;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_168 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'ha8 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_168 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_168 <= _GEN_2254;
      end
    end else begin
      valid_168 <= _GEN_2254;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_169 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'ha9 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_169 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_169 <= _GEN_2255;
      end
    end else begin
      valid_169 <= _GEN_2255;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_170 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'haa == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_170 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_170 <= _GEN_2256;
      end
    end else begin
      valid_170 <= _GEN_2256;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_171 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hab == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_171 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_171 <= _GEN_2257;
      end
    end else begin
      valid_171 <= _GEN_2257;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_172 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hac == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_172 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_172 <= _GEN_2258;
      end
    end else begin
      valid_172 <= _GEN_2258;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_173 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'had == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_173 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_173 <= _GEN_2259;
      end
    end else begin
      valid_173 <= _GEN_2259;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_174 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hae == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_174 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_174 <= _GEN_2260;
      end
    end else begin
      valid_174 <= _GEN_2260;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_175 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'haf == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_175 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_175 <= _GEN_2261;
      end
    end else begin
      valid_175 <= _GEN_2261;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_176 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hb0 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_176 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_176 <= _GEN_2262;
      end
    end else begin
      valid_176 <= _GEN_2262;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_177 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hb1 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_177 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_177 <= _GEN_2263;
      end
    end else begin
      valid_177 <= _GEN_2263;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_178 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hb2 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_178 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_178 <= _GEN_2264;
      end
    end else begin
      valid_178 <= _GEN_2264;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_179 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hb3 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_179 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_179 <= _GEN_2265;
      end
    end else begin
      valid_179 <= _GEN_2265;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_180 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hb4 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_180 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_180 <= _GEN_2266;
      end
    end else begin
      valid_180 <= _GEN_2266;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_181 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hb5 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_181 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_181 <= _GEN_2267;
      end
    end else begin
      valid_181 <= _GEN_2267;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_182 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hb6 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_182 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_182 <= _GEN_2268;
      end
    end else begin
      valid_182 <= _GEN_2268;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_183 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hb7 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_183 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_183 <= _GEN_2269;
      end
    end else begin
      valid_183 <= _GEN_2269;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_184 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hb8 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_184 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_184 <= _GEN_2270;
      end
    end else begin
      valid_184 <= _GEN_2270;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_185 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hb9 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_185 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_185 <= _GEN_2271;
      end
    end else begin
      valid_185 <= _GEN_2271;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_186 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hba == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_186 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_186 <= _GEN_2272;
      end
    end else begin
      valid_186 <= _GEN_2272;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_187 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hbb == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_187 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_187 <= _GEN_2273;
      end
    end else begin
      valid_187 <= _GEN_2273;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_188 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hbc == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_188 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_188 <= _GEN_2274;
      end
    end else begin
      valid_188 <= _GEN_2274;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_189 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hbd == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_189 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_189 <= _GEN_2275;
      end
    end else begin
      valid_189 <= _GEN_2275;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_190 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hbe == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_190 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_190 <= _GEN_2276;
      end
    end else begin
      valid_190 <= _GEN_2276;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_191 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hbf == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_191 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_191 <= _GEN_2277;
      end
    end else begin
      valid_191 <= _GEN_2277;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_192 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hc0 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_192 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_192 <= _GEN_2278;
      end
    end else begin
      valid_192 <= _GEN_2278;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_193 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hc1 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_193 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_193 <= _GEN_2279;
      end
    end else begin
      valid_193 <= _GEN_2279;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_194 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hc2 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_194 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_194 <= _GEN_2280;
      end
    end else begin
      valid_194 <= _GEN_2280;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_195 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hc3 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_195 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_195 <= _GEN_2281;
      end
    end else begin
      valid_195 <= _GEN_2281;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_196 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hc4 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_196 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_196 <= _GEN_2282;
      end
    end else begin
      valid_196 <= _GEN_2282;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_197 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hc5 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_197 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_197 <= _GEN_2283;
      end
    end else begin
      valid_197 <= _GEN_2283;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_198 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hc6 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_198 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_198 <= _GEN_2284;
      end
    end else begin
      valid_198 <= _GEN_2284;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_199 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hc7 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_199 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_199 <= _GEN_2285;
      end
    end else begin
      valid_199 <= _GEN_2285;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_200 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hc8 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_200 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_200 <= _GEN_2286;
      end
    end else begin
      valid_200 <= _GEN_2286;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_201 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hc9 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_201 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_201 <= _GEN_2287;
      end
    end else begin
      valid_201 <= _GEN_2287;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_202 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hca == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_202 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_202 <= _GEN_2288;
      end
    end else begin
      valid_202 <= _GEN_2288;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_203 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hcb == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_203 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_203 <= _GEN_2289;
      end
    end else begin
      valid_203 <= _GEN_2289;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_204 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hcc == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_204 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_204 <= _GEN_2290;
      end
    end else begin
      valid_204 <= _GEN_2290;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_205 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hcd == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_205 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_205 <= _GEN_2291;
      end
    end else begin
      valid_205 <= _GEN_2291;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_206 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hce == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_206 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_206 <= _GEN_2292;
      end
    end else begin
      valid_206 <= _GEN_2292;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_207 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hcf == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_207 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_207 <= _GEN_2293;
      end
    end else begin
      valid_207 <= _GEN_2293;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_208 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hd0 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_208 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_208 <= _GEN_2294;
      end
    end else begin
      valid_208 <= _GEN_2294;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_209 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hd1 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_209 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_209 <= _GEN_2295;
      end
    end else begin
      valid_209 <= _GEN_2295;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_210 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hd2 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_210 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_210 <= _GEN_2296;
      end
    end else begin
      valid_210 <= _GEN_2296;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_211 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hd3 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_211 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_211 <= _GEN_2297;
      end
    end else begin
      valid_211 <= _GEN_2297;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_212 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hd4 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_212 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_212 <= _GEN_2298;
      end
    end else begin
      valid_212 <= _GEN_2298;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_213 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hd5 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_213 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_213 <= _GEN_2299;
      end
    end else begin
      valid_213 <= _GEN_2299;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_214 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hd6 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_214 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_214 <= _GEN_2300;
      end
    end else begin
      valid_214 <= _GEN_2300;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_215 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hd7 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_215 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_215 <= _GEN_2301;
      end
    end else begin
      valid_215 <= _GEN_2301;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_216 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hd8 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_216 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_216 <= _GEN_2302;
      end
    end else begin
      valid_216 <= _GEN_2302;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_217 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hd9 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_217 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_217 <= _GEN_2303;
      end
    end else begin
      valid_217 <= _GEN_2303;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_218 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hda == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_218 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_218 <= _GEN_2304;
      end
    end else begin
      valid_218 <= _GEN_2304;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_219 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hdb == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_219 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_219 <= _GEN_2305;
      end
    end else begin
      valid_219 <= _GEN_2305;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_220 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hdc == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_220 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_220 <= _GEN_2306;
      end
    end else begin
      valid_220 <= _GEN_2306;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_221 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hdd == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_221 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_221 <= _GEN_2307;
      end
    end else begin
      valid_221 <= _GEN_2307;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_222 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hde == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_222 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_222 <= _GEN_2308;
      end
    end else begin
      valid_222 <= _GEN_2308;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_223 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hdf == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_223 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_223 <= _GEN_2309;
      end
    end else begin
      valid_223 <= _GEN_2309;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_224 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'he0 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_224 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_224 <= _GEN_2310;
      end
    end else begin
      valid_224 <= _GEN_2310;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_225 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'he1 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_225 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_225 <= _GEN_2311;
      end
    end else begin
      valid_225 <= _GEN_2311;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_226 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'he2 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_226 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_226 <= _GEN_2312;
      end
    end else begin
      valid_226 <= _GEN_2312;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_227 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'he3 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_227 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_227 <= _GEN_2313;
      end
    end else begin
      valid_227 <= _GEN_2313;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_228 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'he4 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_228 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_228 <= _GEN_2314;
      end
    end else begin
      valid_228 <= _GEN_2314;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_229 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'he5 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_229 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_229 <= _GEN_2315;
      end
    end else begin
      valid_229 <= _GEN_2315;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_230 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'he6 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_230 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_230 <= _GEN_2316;
      end
    end else begin
      valid_230 <= _GEN_2316;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_231 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'he7 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_231 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_231 <= _GEN_2317;
      end
    end else begin
      valid_231 <= _GEN_2317;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_232 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'he8 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_232 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_232 <= _GEN_2318;
      end
    end else begin
      valid_232 <= _GEN_2318;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_233 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'he9 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_233 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_233 <= _GEN_2319;
      end
    end else begin
      valid_233 <= _GEN_2319;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_234 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hea == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_234 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_234 <= _GEN_2320;
      end
    end else begin
      valid_234 <= _GEN_2320;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_235 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'heb == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_235 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_235 <= _GEN_2321;
      end
    end else begin
      valid_235 <= _GEN_2321;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_236 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hec == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_236 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_236 <= _GEN_2322;
      end
    end else begin
      valid_236 <= _GEN_2322;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_237 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hed == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_237 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_237 <= _GEN_2323;
      end
    end else begin
      valid_237 <= _GEN_2323;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_238 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hee == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_238 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_238 <= _GEN_2324;
      end
    end else begin
      valid_238 <= _GEN_2324;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_239 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hef == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_239 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_239 <= _GEN_2325;
      end
    end else begin
      valid_239 <= _GEN_2325;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_240 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hf0 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_240 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_240 <= _GEN_2326;
      end
    end else begin
      valid_240 <= _GEN_2326;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_241 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hf1 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_241 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_241 <= _GEN_2327;
      end
    end else begin
      valid_241 <= _GEN_2327;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_242 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hf2 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_242 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_242 <= _GEN_2328;
      end
    end else begin
      valid_242 <= _GEN_2328;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_243 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hf3 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_243 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_243 <= _GEN_2329;
      end
    end else begin
      valid_243 <= _GEN_2329;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_244 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hf4 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_244 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_244 <= _GEN_2330;
      end
    end else begin
      valid_244 <= _GEN_2330;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_245 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hf5 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_245 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_245 <= _GEN_2331;
      end
    end else begin
      valid_245 <= _GEN_2331;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_246 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hf6 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_246 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_246 <= _GEN_2332;
      end
    end else begin
      valid_246 <= _GEN_2332;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_247 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hf7 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_247 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_247 <= _GEN_2333;
      end
    end else begin
      valid_247 <= _GEN_2333;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_248 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hf8 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_248 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_248 <= _GEN_2334;
      end
    end else begin
      valid_248 <= _GEN_2334;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_249 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hf9 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_249 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_249 <= _GEN_2335;
      end
    end else begin
      valid_249 <= _GEN_2335;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_250 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hfa == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_250 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_250 <= _GEN_2336;
      end
    end else begin
      valid_250 <= _GEN_2336;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_251 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hfb == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_251 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_251 <= _GEN_2337;
      end
    end else begin
      valid_251 <= _GEN_2337;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_252 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hfc == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_252 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_252 <= _GEN_2338;
      end
    end else begin
      valid_252 <= _GEN_2338;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_253 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hfd == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_253 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_253 <= _GEN_2339;
      end
    end else begin
      valid_253 <= _GEN_2339;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_254 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hfe == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_254 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_254 <= _GEN_2340;
      end
    end else begin
      valid_254 <= _GEN_2340;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_255 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'hff == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_255 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_255 <= _GEN_2341;
      end
    end else begin
      valid_255 <= _GEN_2341;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_256 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h100 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_256 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_256 <= _GEN_2342;
      end
    end else begin
      valid_256 <= _GEN_2342;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_257 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h101 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_257 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_257 <= _GEN_2343;
      end
    end else begin
      valid_257 <= _GEN_2343;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_258 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h102 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_258 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_258 <= _GEN_2344;
      end
    end else begin
      valid_258 <= _GEN_2344;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_259 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h103 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_259 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_259 <= _GEN_2345;
      end
    end else begin
      valid_259 <= _GEN_2345;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_260 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h104 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_260 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_260 <= _GEN_2346;
      end
    end else begin
      valid_260 <= _GEN_2346;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_261 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h105 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_261 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_261 <= _GEN_2347;
      end
    end else begin
      valid_261 <= _GEN_2347;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_262 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h106 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_262 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_262 <= _GEN_2348;
      end
    end else begin
      valid_262 <= _GEN_2348;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_263 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h107 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_263 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_263 <= _GEN_2349;
      end
    end else begin
      valid_263 <= _GEN_2349;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_264 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h108 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_264 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_264 <= _GEN_2350;
      end
    end else begin
      valid_264 <= _GEN_2350;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_265 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h109 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_265 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_265 <= _GEN_2351;
      end
    end else begin
      valid_265 <= _GEN_2351;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_266 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h10a == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_266 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_266 <= _GEN_2352;
      end
    end else begin
      valid_266 <= _GEN_2352;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_267 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h10b == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_267 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_267 <= _GEN_2353;
      end
    end else begin
      valid_267 <= _GEN_2353;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_268 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h10c == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_268 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_268 <= _GEN_2354;
      end
    end else begin
      valid_268 <= _GEN_2354;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_269 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h10d == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_269 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_269 <= _GEN_2355;
      end
    end else begin
      valid_269 <= _GEN_2355;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_270 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h10e == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_270 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_270 <= _GEN_2356;
      end
    end else begin
      valid_270 <= _GEN_2356;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_271 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h10f == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_271 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_271 <= _GEN_2357;
      end
    end else begin
      valid_271 <= _GEN_2357;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_272 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h110 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_272 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_272 <= _GEN_2358;
      end
    end else begin
      valid_272 <= _GEN_2358;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_273 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h111 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_273 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_273 <= _GEN_2359;
      end
    end else begin
      valid_273 <= _GEN_2359;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_274 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h112 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_274 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_274 <= _GEN_2360;
      end
    end else begin
      valid_274 <= _GEN_2360;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_275 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h113 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_275 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_275 <= _GEN_2361;
      end
    end else begin
      valid_275 <= _GEN_2361;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_276 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h114 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_276 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_276 <= _GEN_2362;
      end
    end else begin
      valid_276 <= _GEN_2362;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_277 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h115 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_277 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_277 <= _GEN_2363;
      end
    end else begin
      valid_277 <= _GEN_2363;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_278 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h116 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_278 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_278 <= _GEN_2364;
      end
    end else begin
      valid_278 <= _GEN_2364;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_279 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h117 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_279 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_279 <= _GEN_2365;
      end
    end else begin
      valid_279 <= _GEN_2365;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_280 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h118 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_280 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_280 <= _GEN_2366;
      end
    end else begin
      valid_280 <= _GEN_2366;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_281 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h119 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_281 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_281 <= _GEN_2367;
      end
    end else begin
      valid_281 <= _GEN_2367;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_282 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h11a == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_282 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_282 <= _GEN_2368;
      end
    end else begin
      valid_282 <= _GEN_2368;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_283 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h11b == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_283 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_283 <= _GEN_2369;
      end
    end else begin
      valid_283 <= _GEN_2369;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_284 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h11c == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_284 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_284 <= _GEN_2370;
      end
    end else begin
      valid_284 <= _GEN_2370;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_285 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h11d == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_285 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_285 <= _GEN_2371;
      end
    end else begin
      valid_285 <= _GEN_2371;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_286 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h11e == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_286 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_286 <= _GEN_2372;
      end
    end else begin
      valid_286 <= _GEN_2372;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_287 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h11f == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_287 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_287 <= _GEN_2373;
      end
    end else begin
      valid_287 <= _GEN_2373;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_288 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h120 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_288 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_288 <= _GEN_2374;
      end
    end else begin
      valid_288 <= _GEN_2374;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_289 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h121 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_289 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_289 <= _GEN_2375;
      end
    end else begin
      valid_289 <= _GEN_2375;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_290 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h122 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_290 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_290 <= _GEN_2376;
      end
    end else begin
      valid_290 <= _GEN_2376;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_291 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h123 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_291 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_291 <= _GEN_2377;
      end
    end else begin
      valid_291 <= _GEN_2377;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_292 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h124 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_292 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_292 <= _GEN_2378;
      end
    end else begin
      valid_292 <= _GEN_2378;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_293 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h125 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_293 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_293 <= _GEN_2379;
      end
    end else begin
      valid_293 <= _GEN_2379;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_294 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h126 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_294 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_294 <= _GEN_2380;
      end
    end else begin
      valid_294 <= _GEN_2380;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_295 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h127 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_295 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_295 <= _GEN_2381;
      end
    end else begin
      valid_295 <= _GEN_2381;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_296 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h128 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_296 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_296 <= _GEN_2382;
      end
    end else begin
      valid_296 <= _GEN_2382;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_297 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h129 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_297 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_297 <= _GEN_2383;
      end
    end else begin
      valid_297 <= _GEN_2383;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_298 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h12a == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_298 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_298 <= _GEN_2384;
      end
    end else begin
      valid_298 <= _GEN_2384;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_299 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h12b == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_299 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_299 <= _GEN_2385;
      end
    end else begin
      valid_299 <= _GEN_2385;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_300 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h12c == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_300 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_300 <= _GEN_2386;
      end
    end else begin
      valid_300 <= _GEN_2386;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_301 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h12d == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_301 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_301 <= _GEN_2387;
      end
    end else begin
      valid_301 <= _GEN_2387;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_302 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h12e == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_302 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_302 <= _GEN_2388;
      end
    end else begin
      valid_302 <= _GEN_2388;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_303 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h12f == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_303 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_303 <= _GEN_2389;
      end
    end else begin
      valid_303 <= _GEN_2389;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_304 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h130 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_304 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_304 <= _GEN_2390;
      end
    end else begin
      valid_304 <= _GEN_2390;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_305 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h131 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_305 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_305 <= _GEN_2391;
      end
    end else begin
      valid_305 <= _GEN_2391;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_306 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h132 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_306 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_306 <= _GEN_2392;
      end
    end else begin
      valid_306 <= _GEN_2392;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_307 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h133 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_307 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_307 <= _GEN_2393;
      end
    end else begin
      valid_307 <= _GEN_2393;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_308 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h134 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_308 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_308 <= _GEN_2394;
      end
    end else begin
      valid_308 <= _GEN_2394;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_309 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h135 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_309 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_309 <= _GEN_2395;
      end
    end else begin
      valid_309 <= _GEN_2395;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_310 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h136 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_310 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_310 <= _GEN_2396;
      end
    end else begin
      valid_310 <= _GEN_2396;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_311 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h137 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_311 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_311 <= _GEN_2397;
      end
    end else begin
      valid_311 <= _GEN_2397;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_312 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h138 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_312 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_312 <= _GEN_2398;
      end
    end else begin
      valid_312 <= _GEN_2398;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_313 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h139 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_313 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_313 <= _GEN_2399;
      end
    end else begin
      valid_313 <= _GEN_2399;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_314 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h13a == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_314 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_314 <= _GEN_2400;
      end
    end else begin
      valid_314 <= _GEN_2400;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_315 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h13b == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_315 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_315 <= _GEN_2401;
      end
    end else begin
      valid_315 <= _GEN_2401;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_316 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h13c == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_316 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_316 <= _GEN_2402;
      end
    end else begin
      valid_316 <= _GEN_2402;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_317 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h13d == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_317 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_317 <= _GEN_2403;
      end
    end else begin
      valid_317 <= _GEN_2403;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_318 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h13e == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_318 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_318 <= _GEN_2404;
      end
    end else begin
      valid_318 <= _GEN_2404;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_319 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h13f == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_319 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_319 <= _GEN_2405;
      end
    end else begin
      valid_319 <= _GEN_2405;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_320 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h140 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_320 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_320 <= _GEN_2406;
      end
    end else begin
      valid_320 <= _GEN_2406;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_321 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h141 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_321 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_321 <= _GEN_2407;
      end
    end else begin
      valid_321 <= _GEN_2407;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_322 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h142 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_322 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_322 <= _GEN_2408;
      end
    end else begin
      valid_322 <= _GEN_2408;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_323 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h143 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_323 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_323 <= _GEN_2409;
      end
    end else begin
      valid_323 <= _GEN_2409;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_324 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h144 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_324 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_324 <= _GEN_2410;
      end
    end else begin
      valid_324 <= _GEN_2410;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_325 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h145 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_325 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_325 <= _GEN_2411;
      end
    end else begin
      valid_325 <= _GEN_2411;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_326 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h146 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_326 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_326 <= _GEN_2412;
      end
    end else begin
      valid_326 <= _GEN_2412;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_327 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h147 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_327 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_327 <= _GEN_2413;
      end
    end else begin
      valid_327 <= _GEN_2413;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_328 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h148 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_328 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_328 <= _GEN_2414;
      end
    end else begin
      valid_328 <= _GEN_2414;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_329 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h149 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_329 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_329 <= _GEN_2415;
      end
    end else begin
      valid_329 <= _GEN_2415;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_330 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h14a == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_330 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_330 <= _GEN_2416;
      end
    end else begin
      valid_330 <= _GEN_2416;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_331 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h14b == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_331 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_331 <= _GEN_2417;
      end
    end else begin
      valid_331 <= _GEN_2417;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_332 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h14c == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_332 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_332 <= _GEN_2418;
      end
    end else begin
      valid_332 <= _GEN_2418;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_333 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h14d == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_333 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_333 <= _GEN_2419;
      end
    end else begin
      valid_333 <= _GEN_2419;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_334 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h14e == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_334 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_334 <= _GEN_2420;
      end
    end else begin
      valid_334 <= _GEN_2420;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_335 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h14f == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_335 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_335 <= _GEN_2421;
      end
    end else begin
      valid_335 <= _GEN_2421;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_336 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h150 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_336 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_336 <= _GEN_2422;
      end
    end else begin
      valid_336 <= _GEN_2422;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_337 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h151 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_337 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_337 <= _GEN_2423;
      end
    end else begin
      valid_337 <= _GEN_2423;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_338 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h152 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_338 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_338 <= _GEN_2424;
      end
    end else begin
      valid_338 <= _GEN_2424;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_339 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h153 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_339 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_339 <= _GEN_2425;
      end
    end else begin
      valid_339 <= _GEN_2425;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_340 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h154 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_340 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_340 <= _GEN_2426;
      end
    end else begin
      valid_340 <= _GEN_2426;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_341 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h155 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_341 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_341 <= _GEN_2427;
      end
    end else begin
      valid_341 <= _GEN_2427;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_342 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h156 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_342 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_342 <= _GEN_2428;
      end
    end else begin
      valid_342 <= _GEN_2428;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_343 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h157 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_343 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_343 <= _GEN_2429;
      end
    end else begin
      valid_343 <= _GEN_2429;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_344 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h158 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_344 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_344 <= _GEN_2430;
      end
    end else begin
      valid_344 <= _GEN_2430;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_345 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h159 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_345 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_345 <= _GEN_2431;
      end
    end else begin
      valid_345 <= _GEN_2431;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_346 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h15a == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_346 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_346 <= _GEN_2432;
      end
    end else begin
      valid_346 <= _GEN_2432;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_347 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h15b == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_347 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_347 <= _GEN_2433;
      end
    end else begin
      valid_347 <= _GEN_2433;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_348 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h15c == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_348 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_348 <= _GEN_2434;
      end
    end else begin
      valid_348 <= _GEN_2434;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_349 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h15d == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_349 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_349 <= _GEN_2435;
      end
    end else begin
      valid_349 <= _GEN_2435;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_350 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h15e == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_350 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_350 <= _GEN_2436;
      end
    end else begin
      valid_350 <= _GEN_2436;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_351 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h15f == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_351 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_351 <= _GEN_2437;
      end
    end else begin
      valid_351 <= _GEN_2437;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_352 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h160 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_352 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_352 <= _GEN_2438;
      end
    end else begin
      valid_352 <= _GEN_2438;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_353 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h161 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_353 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_353 <= _GEN_2439;
      end
    end else begin
      valid_353 <= _GEN_2439;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_354 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h162 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_354 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_354 <= _GEN_2440;
      end
    end else begin
      valid_354 <= _GEN_2440;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_355 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h163 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_355 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_355 <= _GEN_2441;
      end
    end else begin
      valid_355 <= _GEN_2441;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_356 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h164 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_356 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_356 <= _GEN_2442;
      end
    end else begin
      valid_356 <= _GEN_2442;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_357 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h165 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_357 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_357 <= _GEN_2443;
      end
    end else begin
      valid_357 <= _GEN_2443;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_358 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h166 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_358 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_358 <= _GEN_2444;
      end
    end else begin
      valid_358 <= _GEN_2444;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_359 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h167 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_359 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_359 <= _GEN_2445;
      end
    end else begin
      valid_359 <= _GEN_2445;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_360 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h168 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_360 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_360 <= _GEN_2446;
      end
    end else begin
      valid_360 <= _GEN_2446;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_361 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h169 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_361 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_361 <= _GEN_2447;
      end
    end else begin
      valid_361 <= _GEN_2447;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_362 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h16a == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_362 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_362 <= _GEN_2448;
      end
    end else begin
      valid_362 <= _GEN_2448;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_363 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h16b == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_363 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_363 <= _GEN_2449;
      end
    end else begin
      valid_363 <= _GEN_2449;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_364 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h16c == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_364 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_364 <= _GEN_2450;
      end
    end else begin
      valid_364 <= _GEN_2450;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_365 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h16d == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_365 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_365 <= _GEN_2451;
      end
    end else begin
      valid_365 <= _GEN_2451;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_366 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h16e == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_366 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_366 <= _GEN_2452;
      end
    end else begin
      valid_366 <= _GEN_2452;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_367 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h16f == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_367 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_367 <= _GEN_2453;
      end
    end else begin
      valid_367 <= _GEN_2453;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_368 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h170 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_368 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_368 <= _GEN_2454;
      end
    end else begin
      valid_368 <= _GEN_2454;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_369 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h171 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_369 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_369 <= _GEN_2455;
      end
    end else begin
      valid_369 <= _GEN_2455;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_370 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h172 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_370 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_370 <= _GEN_2456;
      end
    end else begin
      valid_370 <= _GEN_2456;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_371 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h173 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_371 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_371 <= _GEN_2457;
      end
    end else begin
      valid_371 <= _GEN_2457;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_372 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h174 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_372 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_372 <= _GEN_2458;
      end
    end else begin
      valid_372 <= _GEN_2458;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_373 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h175 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_373 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_373 <= _GEN_2459;
      end
    end else begin
      valid_373 <= _GEN_2459;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_374 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h176 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_374 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_374 <= _GEN_2460;
      end
    end else begin
      valid_374 <= _GEN_2460;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_375 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h177 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_375 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_375 <= _GEN_2461;
      end
    end else begin
      valid_375 <= _GEN_2461;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_376 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h178 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_376 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_376 <= _GEN_2462;
      end
    end else begin
      valid_376 <= _GEN_2462;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_377 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h179 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_377 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_377 <= _GEN_2463;
      end
    end else begin
      valid_377 <= _GEN_2463;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_378 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h17a == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_378 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_378 <= _GEN_2464;
      end
    end else begin
      valid_378 <= _GEN_2464;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_379 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h17b == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_379 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_379 <= _GEN_2465;
      end
    end else begin
      valid_379 <= _GEN_2465;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_380 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h17c == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_380 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_380 <= _GEN_2466;
      end
    end else begin
      valid_380 <= _GEN_2466;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_381 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h17d == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_381 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_381 <= _GEN_2467;
      end
    end else begin
      valid_381 <= _GEN_2467;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_382 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h17e == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_382 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_382 <= _GEN_2468;
      end
    end else begin
      valid_382 <= _GEN_2468;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_383 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h17f == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_383 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_383 <= _GEN_2469;
      end
    end else begin
      valid_383 <= _GEN_2469;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_384 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h180 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_384 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_384 <= _GEN_2470;
      end
    end else begin
      valid_384 <= _GEN_2470;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_385 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h181 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_385 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_385 <= _GEN_2471;
      end
    end else begin
      valid_385 <= _GEN_2471;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_386 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h182 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_386 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_386 <= _GEN_2472;
      end
    end else begin
      valid_386 <= _GEN_2472;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_387 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h183 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_387 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_387 <= _GEN_2473;
      end
    end else begin
      valid_387 <= _GEN_2473;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_388 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h184 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_388 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_388 <= _GEN_2474;
      end
    end else begin
      valid_388 <= _GEN_2474;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_389 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h185 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_389 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_389 <= _GEN_2475;
      end
    end else begin
      valid_389 <= _GEN_2475;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_390 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h186 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_390 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_390 <= _GEN_2476;
      end
    end else begin
      valid_390 <= _GEN_2476;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_391 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h187 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_391 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_391 <= _GEN_2477;
      end
    end else begin
      valid_391 <= _GEN_2477;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_392 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h188 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_392 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_392 <= _GEN_2478;
      end
    end else begin
      valid_392 <= _GEN_2478;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_393 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h189 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_393 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_393 <= _GEN_2479;
      end
    end else begin
      valid_393 <= _GEN_2479;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_394 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h18a == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_394 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_394 <= _GEN_2480;
      end
    end else begin
      valid_394 <= _GEN_2480;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_395 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h18b == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_395 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_395 <= _GEN_2481;
      end
    end else begin
      valid_395 <= _GEN_2481;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_396 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h18c == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_396 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_396 <= _GEN_2482;
      end
    end else begin
      valid_396 <= _GEN_2482;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_397 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h18d == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_397 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_397 <= _GEN_2483;
      end
    end else begin
      valid_397 <= _GEN_2483;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_398 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h18e == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_398 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_398 <= _GEN_2484;
      end
    end else begin
      valid_398 <= _GEN_2484;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_399 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h18f == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_399 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_399 <= _GEN_2485;
      end
    end else begin
      valid_399 <= _GEN_2485;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_400 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h190 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_400 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_400 <= _GEN_2486;
      end
    end else begin
      valid_400 <= _GEN_2486;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_401 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h191 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_401 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_401 <= _GEN_2487;
      end
    end else begin
      valid_401 <= _GEN_2487;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_402 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h192 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_402 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_402 <= _GEN_2488;
      end
    end else begin
      valid_402 <= _GEN_2488;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_403 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h193 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_403 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_403 <= _GEN_2489;
      end
    end else begin
      valid_403 <= _GEN_2489;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_404 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h194 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_404 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_404 <= _GEN_2490;
      end
    end else begin
      valid_404 <= _GEN_2490;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_405 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h195 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_405 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_405 <= _GEN_2491;
      end
    end else begin
      valid_405 <= _GEN_2491;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_406 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h196 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_406 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_406 <= _GEN_2492;
      end
    end else begin
      valid_406 <= _GEN_2492;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_407 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h197 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_407 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_407 <= _GEN_2493;
      end
    end else begin
      valid_407 <= _GEN_2493;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_408 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h198 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_408 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_408 <= _GEN_2494;
      end
    end else begin
      valid_408 <= _GEN_2494;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_409 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h199 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_409 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_409 <= _GEN_2495;
      end
    end else begin
      valid_409 <= _GEN_2495;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_410 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h19a == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_410 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_410 <= _GEN_2496;
      end
    end else begin
      valid_410 <= _GEN_2496;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_411 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h19b == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_411 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_411 <= _GEN_2497;
      end
    end else begin
      valid_411 <= _GEN_2497;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_412 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h19c == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_412 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_412 <= _GEN_2498;
      end
    end else begin
      valid_412 <= _GEN_2498;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_413 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h19d == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_413 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_413 <= _GEN_2499;
      end
    end else begin
      valid_413 <= _GEN_2499;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_414 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h19e == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_414 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_414 <= _GEN_2500;
      end
    end else begin
      valid_414 <= _GEN_2500;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_415 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h19f == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_415 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_415 <= _GEN_2501;
      end
    end else begin
      valid_415 <= _GEN_2501;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_416 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1a0 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_416 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_416 <= _GEN_2502;
      end
    end else begin
      valid_416 <= _GEN_2502;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_417 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1a1 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_417 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_417 <= _GEN_2503;
      end
    end else begin
      valid_417 <= _GEN_2503;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_418 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1a2 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_418 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_418 <= _GEN_2504;
      end
    end else begin
      valid_418 <= _GEN_2504;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_419 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1a3 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_419 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_419 <= _GEN_2505;
      end
    end else begin
      valid_419 <= _GEN_2505;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_420 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1a4 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_420 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_420 <= _GEN_2506;
      end
    end else begin
      valid_420 <= _GEN_2506;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_421 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1a5 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_421 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_421 <= _GEN_2507;
      end
    end else begin
      valid_421 <= _GEN_2507;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_422 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1a6 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_422 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_422 <= _GEN_2508;
      end
    end else begin
      valid_422 <= _GEN_2508;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_423 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1a7 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_423 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_423 <= _GEN_2509;
      end
    end else begin
      valid_423 <= _GEN_2509;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_424 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1a8 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_424 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_424 <= _GEN_2510;
      end
    end else begin
      valid_424 <= _GEN_2510;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_425 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1a9 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_425 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_425 <= _GEN_2511;
      end
    end else begin
      valid_425 <= _GEN_2511;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_426 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1aa == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_426 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_426 <= _GEN_2512;
      end
    end else begin
      valid_426 <= _GEN_2512;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_427 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1ab == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_427 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_427 <= _GEN_2513;
      end
    end else begin
      valid_427 <= _GEN_2513;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_428 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1ac == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_428 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_428 <= _GEN_2514;
      end
    end else begin
      valid_428 <= _GEN_2514;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_429 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1ad == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_429 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_429 <= _GEN_2515;
      end
    end else begin
      valid_429 <= _GEN_2515;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_430 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1ae == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_430 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_430 <= _GEN_2516;
      end
    end else begin
      valid_430 <= _GEN_2516;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_431 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1af == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_431 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_431 <= _GEN_2517;
      end
    end else begin
      valid_431 <= _GEN_2517;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_432 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1b0 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_432 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_432 <= _GEN_2518;
      end
    end else begin
      valid_432 <= _GEN_2518;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_433 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1b1 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_433 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_433 <= _GEN_2519;
      end
    end else begin
      valid_433 <= _GEN_2519;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_434 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1b2 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_434 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_434 <= _GEN_2520;
      end
    end else begin
      valid_434 <= _GEN_2520;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_435 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1b3 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_435 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_435 <= _GEN_2521;
      end
    end else begin
      valid_435 <= _GEN_2521;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_436 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1b4 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_436 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_436 <= _GEN_2522;
      end
    end else begin
      valid_436 <= _GEN_2522;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_437 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1b5 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_437 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_437 <= _GEN_2523;
      end
    end else begin
      valid_437 <= _GEN_2523;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_438 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1b6 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_438 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_438 <= _GEN_2524;
      end
    end else begin
      valid_438 <= _GEN_2524;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_439 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1b7 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_439 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_439 <= _GEN_2525;
      end
    end else begin
      valid_439 <= _GEN_2525;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_440 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1b8 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_440 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_440 <= _GEN_2526;
      end
    end else begin
      valid_440 <= _GEN_2526;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_441 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1b9 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_441 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_441 <= _GEN_2527;
      end
    end else begin
      valid_441 <= _GEN_2527;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_442 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1ba == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_442 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_442 <= _GEN_2528;
      end
    end else begin
      valid_442 <= _GEN_2528;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_443 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1bb == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_443 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_443 <= _GEN_2529;
      end
    end else begin
      valid_443 <= _GEN_2529;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_444 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1bc == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_444 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_444 <= _GEN_2530;
      end
    end else begin
      valid_444 <= _GEN_2530;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_445 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1bd == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_445 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_445 <= _GEN_2531;
      end
    end else begin
      valid_445 <= _GEN_2531;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_446 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1be == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_446 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_446 <= _GEN_2532;
      end
    end else begin
      valid_446 <= _GEN_2532;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_447 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1bf == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_447 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_447 <= _GEN_2533;
      end
    end else begin
      valid_447 <= _GEN_2533;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_448 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1c0 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_448 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_448 <= _GEN_2534;
      end
    end else begin
      valid_448 <= _GEN_2534;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_449 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1c1 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_449 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_449 <= _GEN_2535;
      end
    end else begin
      valid_449 <= _GEN_2535;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_450 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1c2 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_450 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_450 <= _GEN_2536;
      end
    end else begin
      valid_450 <= _GEN_2536;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_451 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1c3 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_451 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_451 <= _GEN_2537;
      end
    end else begin
      valid_451 <= _GEN_2537;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_452 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1c4 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_452 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_452 <= _GEN_2538;
      end
    end else begin
      valid_452 <= _GEN_2538;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_453 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1c5 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_453 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_453 <= _GEN_2539;
      end
    end else begin
      valid_453 <= _GEN_2539;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_454 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1c6 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_454 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_454 <= _GEN_2540;
      end
    end else begin
      valid_454 <= _GEN_2540;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_455 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1c7 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_455 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_455 <= _GEN_2541;
      end
    end else begin
      valid_455 <= _GEN_2541;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_456 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1c8 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_456 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_456 <= _GEN_2542;
      end
    end else begin
      valid_456 <= _GEN_2542;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_457 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1c9 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_457 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_457 <= _GEN_2543;
      end
    end else begin
      valid_457 <= _GEN_2543;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_458 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1ca == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_458 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_458 <= _GEN_2544;
      end
    end else begin
      valid_458 <= _GEN_2544;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_459 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1cb == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_459 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_459 <= _GEN_2545;
      end
    end else begin
      valid_459 <= _GEN_2545;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_460 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1cc == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_460 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_460 <= _GEN_2546;
      end
    end else begin
      valid_460 <= _GEN_2546;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_461 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1cd == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_461 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_461 <= _GEN_2547;
      end
    end else begin
      valid_461 <= _GEN_2547;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_462 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1ce == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_462 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_462 <= _GEN_2548;
      end
    end else begin
      valid_462 <= _GEN_2548;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_463 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1cf == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_463 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_463 <= _GEN_2549;
      end
    end else begin
      valid_463 <= _GEN_2549;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_464 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1d0 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_464 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_464 <= _GEN_2550;
      end
    end else begin
      valid_464 <= _GEN_2550;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_465 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1d1 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_465 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_465 <= _GEN_2551;
      end
    end else begin
      valid_465 <= _GEN_2551;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_466 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1d2 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_466 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_466 <= _GEN_2552;
      end
    end else begin
      valid_466 <= _GEN_2552;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_467 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1d3 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_467 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_467 <= _GEN_2553;
      end
    end else begin
      valid_467 <= _GEN_2553;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_468 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1d4 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_468 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_468 <= _GEN_2554;
      end
    end else begin
      valid_468 <= _GEN_2554;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_469 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1d5 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_469 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_469 <= _GEN_2555;
      end
    end else begin
      valid_469 <= _GEN_2555;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_470 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1d6 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_470 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_470 <= _GEN_2556;
      end
    end else begin
      valid_470 <= _GEN_2556;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_471 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1d7 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_471 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_471 <= _GEN_2557;
      end
    end else begin
      valid_471 <= _GEN_2557;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_472 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1d8 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_472 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_472 <= _GEN_2558;
      end
    end else begin
      valid_472 <= _GEN_2558;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_473 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1d9 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_473 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_473 <= _GEN_2559;
      end
    end else begin
      valid_473 <= _GEN_2559;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_474 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1da == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_474 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_474 <= _GEN_2560;
      end
    end else begin
      valid_474 <= _GEN_2560;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_475 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1db == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_475 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_475 <= _GEN_2561;
      end
    end else begin
      valid_475 <= _GEN_2561;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_476 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1dc == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_476 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_476 <= _GEN_2562;
      end
    end else begin
      valid_476 <= _GEN_2562;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_477 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1dd == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_477 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_477 <= _GEN_2563;
      end
    end else begin
      valid_477 <= _GEN_2563;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_478 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1de == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_478 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_478 <= _GEN_2564;
      end
    end else begin
      valid_478 <= _GEN_2564;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_479 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1df == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_479 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_479 <= _GEN_2565;
      end
    end else begin
      valid_479 <= _GEN_2565;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_480 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1e0 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_480 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_480 <= _GEN_2566;
      end
    end else begin
      valid_480 <= _GEN_2566;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_481 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1e1 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_481 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_481 <= _GEN_2567;
      end
    end else begin
      valid_481 <= _GEN_2567;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_482 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1e2 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_482 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_482 <= _GEN_2568;
      end
    end else begin
      valid_482 <= _GEN_2568;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_483 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1e3 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_483 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_483 <= _GEN_2569;
      end
    end else begin
      valid_483 <= _GEN_2569;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_484 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1e4 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_484 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_484 <= _GEN_2570;
      end
    end else begin
      valid_484 <= _GEN_2570;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_485 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1e5 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_485 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_485 <= _GEN_2571;
      end
    end else begin
      valid_485 <= _GEN_2571;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_486 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1e6 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_486 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_486 <= _GEN_2572;
      end
    end else begin
      valid_486 <= _GEN_2572;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_487 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1e7 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_487 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_487 <= _GEN_2573;
      end
    end else begin
      valid_487 <= _GEN_2573;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_488 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1e8 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_488 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_488 <= _GEN_2574;
      end
    end else begin
      valid_488 <= _GEN_2574;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_489 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1e9 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_489 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_489 <= _GEN_2575;
      end
    end else begin
      valid_489 <= _GEN_2575;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_490 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1ea == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_490 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_490 <= _GEN_2576;
      end
    end else begin
      valid_490 <= _GEN_2576;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_491 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1eb == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_491 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_491 <= _GEN_2577;
      end
    end else begin
      valid_491 <= _GEN_2577;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_492 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1ec == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_492 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_492 <= _GEN_2578;
      end
    end else begin
      valid_492 <= _GEN_2578;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_493 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1ed == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_493 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_493 <= _GEN_2579;
      end
    end else begin
      valid_493 <= _GEN_2579;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_494 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1ee == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_494 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_494 <= _GEN_2580;
      end
    end else begin
      valid_494 <= _GEN_2580;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_495 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1ef == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_495 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_495 <= _GEN_2581;
      end
    end else begin
      valid_495 <= _GEN_2581;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_496 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1f0 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_496 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_496 <= _GEN_2582;
      end
    end else begin
      valid_496 <= _GEN_2582;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_497 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1f1 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_497 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_497 <= _GEN_2583;
      end
    end else begin
      valid_497 <= _GEN_2583;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_498 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1f2 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_498 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_498 <= _GEN_2584;
      end
    end else begin
      valid_498 <= _GEN_2584;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_499 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1f3 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_499 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_499 <= _GEN_2585;
      end
    end else begin
      valid_499 <= _GEN_2585;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_500 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1f4 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_500 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_500 <= _GEN_2586;
      end
    end else begin
      valid_500 <= _GEN_2586;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_501 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1f5 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_501 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_501 <= _GEN_2587;
      end
    end else begin
      valid_501 <= _GEN_2587;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_502 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1f6 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_502 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_502 <= _GEN_2588;
      end
    end else begin
      valid_502 <= _GEN_2588;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_503 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1f7 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_503 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_503 <= _GEN_2589;
      end
    end else begin
      valid_503 <= _GEN_2589;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_504 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1f8 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_504 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_504 <= _GEN_2590;
      end
    end else begin
      valid_504 <= _GEN_2590;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_505 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1f9 == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_505 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_505 <= _GEN_2591;
      end
    end else begin
      valid_505 <= _GEN_2591;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_506 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1fa == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_506 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_506 <= _GEN_2592;
      end
    end else begin
      valid_506 <= _GEN_2592;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_507 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1fb == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_507 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_507 <= _GEN_2593;
      end
    end else begin
      valid_507 <= _GEN_2593;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_508 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1fc == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_508 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_508 <= _GEN_2594;
      end
    end else begin
      valid_508 <= _GEN_2594;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_509 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1fd == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_509 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_509 <= _GEN_2595;
      end
    end else begin
      valid_509 <= _GEN_2595;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_510 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1fe == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_510 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_510 <= _GEN_2596;
      end
    end else begin
      valid_510 <= _GEN_2596;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_511 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (9'h1ff == _GEN_4[13:5]) begin // @[DCache.scala 241:33]
        valid_511 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_511 <= _GEN_2597;
      end
    end else begin
      valid_511 <= _GEN_2597;
    end
    array_out_REG <= io_cache_req_ready & io_cache_req_valid; // @[Decoupled.scala 51:35]
    if (reset) begin // @[Reg.scala 35:20]
      array_out_r <= 274'h0; // @[Reg.scala 35:20]
    end else if (array_out_REG) begin // @[Utils.scala 50:8]
      array_out_r <= array_io_rdata;
    end
    if (reset) begin // @[DCache.scala 128:30]
      lrsc_addr <= 27'h0; // @[DCache.scala 128:30]
    end else if (_array_io_en_T_1 & is_lr_r) begin // @[DCache.scala 132:30]
      lrsc_addr <= req_r_addr[31:5]; // @[DCache.scala 134:19]
    end
    if (reset) begin // @[Reg.scala 35:20]
      sc_fail_r <= 1'h0; // @[Reg.scala 35:20]
    end else if (_req_r_T) begin // @[Reg.scala 36:18]
      sc_fail_r <= sc_fail; // @[Reg.scala 36:22]
    end
    probe_out_REG <= tl_b_ready & auto_out_b_valid; // @[Decoupled.scala 51:35]
    if (reset) begin // @[Reg.scala 35:20]
      probe_out_r <= 274'h0; // @[Reg.scala 35:20]
    end else if (probe_out_REG) begin // @[Reg.scala 36:18]
      probe_out_r <= array_io_rdata; // @[Reg.scala 36:22]
    end
    release_addr_aligned_REG <= array_io_addr; // @[DCache.scala 245:56]
    if (reset) begin // @[Counter.scala 61:40]
      source <= 2'h0; // @[Counter.scala 61:40]
    end else if (_source_T_2) begin // @[Counter.scala 118:16]
      source <= _source_wrap_value_T_1; // @[Counter.scala 77:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  probing = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  lrsc_reserved = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  lrsc_counter = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  tl_b_bits_r_size = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  tl_b_bits_r_source = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  tl_b_bits_r_address = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  state = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  tl_d_bits_r_sink = _RAND_7[5:0];
  _RAND_8 = {8{`RANDOM}};
  tl_d_bits_r_data = _RAND_8[255:0];
  _RAND_9 = {2{`RANDOM}};
  req_r_addr = _RAND_9[38:0];
  _RAND_10 = {2{`RANDOM}};
  req_r_wdata = _RAND_10[63:0];
  _RAND_11 = {1{`RANDOM}};
  req_r_wmask = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  req_r_wen = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  req_r_len = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  req_r_lrsc = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  req_r_amo = _RAND_15[4:0];
  _RAND_16 = {1{`RANDOM}};
  valid_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  valid_1 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  valid_2 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  valid_3 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  valid_4 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  valid_5 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  valid_6 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  valid_7 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  valid_8 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  valid_9 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  valid_10 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  valid_11 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  valid_12 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  valid_13 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  valid_14 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  valid_15 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  valid_16 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  valid_17 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  valid_18 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  valid_19 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  valid_20 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  valid_21 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  valid_22 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  valid_23 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  valid_24 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  valid_25 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  valid_26 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  valid_27 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  valid_28 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  valid_29 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  valid_30 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  valid_31 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  valid_32 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  valid_33 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  valid_34 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  valid_35 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  valid_36 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  valid_37 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  valid_38 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  valid_39 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  valid_40 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  valid_41 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  valid_42 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  valid_43 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  valid_44 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  valid_45 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  valid_46 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  valid_47 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  valid_48 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  valid_49 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  valid_50 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  valid_51 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  valid_52 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  valid_53 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  valid_54 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  valid_55 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  valid_56 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  valid_57 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  valid_58 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  valid_59 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  valid_60 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  valid_61 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  valid_62 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  valid_63 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  valid_64 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  valid_65 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  valid_66 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  valid_67 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  valid_68 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  valid_69 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  valid_70 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  valid_71 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  valid_72 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  valid_73 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  valid_74 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  valid_75 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  valid_76 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  valid_77 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  valid_78 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  valid_79 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  valid_80 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  valid_81 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  valid_82 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  valid_83 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  valid_84 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  valid_85 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  valid_86 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  valid_87 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  valid_88 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  valid_89 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  valid_90 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  valid_91 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  valid_92 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  valid_93 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  valid_94 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  valid_95 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  valid_96 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  valid_97 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  valid_98 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  valid_99 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  valid_100 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  valid_101 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  valid_102 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  valid_103 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  valid_104 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  valid_105 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  valid_106 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  valid_107 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  valid_108 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  valid_109 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  valid_110 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  valid_111 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  valid_112 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  valid_113 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  valid_114 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  valid_115 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  valid_116 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  valid_117 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  valid_118 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  valid_119 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  valid_120 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  valid_121 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  valid_122 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  valid_123 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  valid_124 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  valid_125 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  valid_126 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  valid_127 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  valid_128 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  valid_129 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  valid_130 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  valid_131 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  valid_132 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  valid_133 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  valid_134 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  valid_135 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  valid_136 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  valid_137 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  valid_138 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  valid_139 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  valid_140 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  valid_141 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  valid_142 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  valid_143 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  valid_144 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  valid_145 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  valid_146 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  valid_147 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  valid_148 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  valid_149 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  valid_150 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  valid_151 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  valid_152 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  valid_153 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  valid_154 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  valid_155 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  valid_156 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  valid_157 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  valid_158 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  valid_159 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  valid_160 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  valid_161 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  valid_162 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  valid_163 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  valid_164 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  valid_165 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  valid_166 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  valid_167 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  valid_168 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  valid_169 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  valid_170 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  valid_171 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  valid_172 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  valid_173 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  valid_174 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  valid_175 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  valid_176 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  valid_177 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  valid_178 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  valid_179 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  valid_180 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  valid_181 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  valid_182 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  valid_183 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  valid_184 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  valid_185 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  valid_186 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  valid_187 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  valid_188 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  valid_189 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  valid_190 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  valid_191 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  valid_192 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  valid_193 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  valid_194 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  valid_195 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  valid_196 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  valid_197 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  valid_198 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  valid_199 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  valid_200 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  valid_201 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  valid_202 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  valid_203 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  valid_204 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  valid_205 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  valid_206 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  valid_207 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  valid_208 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  valid_209 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  valid_210 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  valid_211 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  valid_212 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  valid_213 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  valid_214 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  valid_215 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  valid_216 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  valid_217 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  valid_218 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  valid_219 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  valid_220 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  valid_221 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  valid_222 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  valid_223 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  valid_224 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  valid_225 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  valid_226 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  valid_227 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  valid_228 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  valid_229 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  valid_230 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  valid_231 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  valid_232 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  valid_233 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  valid_234 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  valid_235 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  valid_236 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  valid_237 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  valid_238 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  valid_239 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  valid_240 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  valid_241 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  valid_242 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  valid_243 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  valid_244 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  valid_245 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  valid_246 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  valid_247 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  valid_248 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  valid_249 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  valid_250 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  valid_251 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  valid_252 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  valid_253 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  valid_254 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  valid_255 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  valid_256 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  valid_257 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  valid_258 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  valid_259 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  valid_260 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  valid_261 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  valid_262 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  valid_263 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  valid_264 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  valid_265 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  valid_266 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  valid_267 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  valid_268 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  valid_269 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  valid_270 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  valid_271 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  valid_272 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  valid_273 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  valid_274 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  valid_275 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  valid_276 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  valid_277 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  valid_278 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  valid_279 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  valid_280 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  valid_281 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  valid_282 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  valid_283 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  valid_284 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  valid_285 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  valid_286 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  valid_287 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  valid_288 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  valid_289 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  valid_290 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  valid_291 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  valid_292 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  valid_293 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  valid_294 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  valid_295 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  valid_296 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  valid_297 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  valid_298 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  valid_299 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  valid_300 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  valid_301 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  valid_302 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  valid_303 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  valid_304 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  valid_305 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  valid_306 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  valid_307 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  valid_308 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  valid_309 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  valid_310 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  valid_311 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  valid_312 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  valid_313 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  valid_314 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  valid_315 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  valid_316 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  valid_317 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  valid_318 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  valid_319 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  valid_320 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  valid_321 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  valid_322 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  valid_323 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  valid_324 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  valid_325 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  valid_326 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  valid_327 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  valid_328 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  valid_329 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  valid_330 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  valid_331 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  valid_332 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  valid_333 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  valid_334 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  valid_335 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  valid_336 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  valid_337 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  valid_338 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  valid_339 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  valid_340 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  valid_341 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  valid_342 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  valid_343 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  valid_344 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  valid_345 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  valid_346 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  valid_347 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  valid_348 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  valid_349 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  valid_350 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  valid_351 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  valid_352 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  valid_353 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  valid_354 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  valid_355 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  valid_356 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  valid_357 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  valid_358 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  valid_359 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  valid_360 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  valid_361 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  valid_362 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  valid_363 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  valid_364 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  valid_365 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  valid_366 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  valid_367 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  valid_368 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  valid_369 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  valid_370 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  valid_371 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  valid_372 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  valid_373 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  valid_374 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  valid_375 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  valid_376 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  valid_377 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  valid_378 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  valid_379 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  valid_380 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  valid_381 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  valid_382 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  valid_383 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  valid_384 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  valid_385 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  valid_386 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  valid_387 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  valid_388 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  valid_389 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  valid_390 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  valid_391 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  valid_392 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  valid_393 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  valid_394 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  valid_395 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  valid_396 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  valid_397 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  valid_398 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  valid_399 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  valid_400 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  valid_401 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  valid_402 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  valid_403 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  valid_404 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  valid_405 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  valid_406 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  valid_407 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  valid_408 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  valid_409 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  valid_410 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  valid_411 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  valid_412 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  valid_413 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  valid_414 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  valid_415 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  valid_416 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  valid_417 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  valid_418 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  valid_419 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  valid_420 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  valid_421 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  valid_422 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  valid_423 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  valid_424 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  valid_425 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  valid_426 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  valid_427 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  valid_428 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  valid_429 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  valid_430 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  valid_431 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  valid_432 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  valid_433 = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  valid_434 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  valid_435 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  valid_436 = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  valid_437 = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  valid_438 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  valid_439 = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  valid_440 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  valid_441 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  valid_442 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  valid_443 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  valid_444 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  valid_445 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  valid_446 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  valid_447 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  valid_448 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  valid_449 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  valid_450 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  valid_451 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  valid_452 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  valid_453 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  valid_454 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  valid_455 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  valid_456 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  valid_457 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  valid_458 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  valid_459 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  valid_460 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  valid_461 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  valid_462 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  valid_463 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  valid_464 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  valid_465 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  valid_466 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  valid_467 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  valid_468 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  valid_469 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  valid_470 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  valid_471 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  valid_472 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  valid_473 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  valid_474 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  valid_475 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  valid_476 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  valid_477 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  valid_478 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  valid_479 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  valid_480 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  valid_481 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  valid_482 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  valid_483 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  valid_484 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  valid_485 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  valid_486 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  valid_487 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  valid_488 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  valid_489 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  valid_490 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  valid_491 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  valid_492 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  valid_493 = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  valid_494 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  valid_495 = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  valid_496 = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  valid_497 = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  valid_498 = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  valid_499 = _RAND_515[0:0];
  _RAND_516 = {1{`RANDOM}};
  valid_500 = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  valid_501 = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  valid_502 = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  valid_503 = _RAND_519[0:0];
  _RAND_520 = {1{`RANDOM}};
  valid_504 = _RAND_520[0:0];
  _RAND_521 = {1{`RANDOM}};
  valid_505 = _RAND_521[0:0];
  _RAND_522 = {1{`RANDOM}};
  valid_506 = _RAND_522[0:0];
  _RAND_523 = {1{`RANDOM}};
  valid_507 = _RAND_523[0:0];
  _RAND_524 = {1{`RANDOM}};
  valid_508 = _RAND_524[0:0];
  _RAND_525 = {1{`RANDOM}};
  valid_509 = _RAND_525[0:0];
  _RAND_526 = {1{`RANDOM}};
  valid_510 = _RAND_526[0:0];
  _RAND_527 = {1{`RANDOM}};
  valid_511 = _RAND_527[0:0];
  _RAND_528 = {1{`RANDOM}};
  array_out_REG = _RAND_528[0:0];
  _RAND_529 = {9{`RANDOM}};
  array_out_r = _RAND_529[273:0];
  _RAND_530 = {1{`RANDOM}};
  lrsc_addr = _RAND_530[26:0];
  _RAND_531 = {1{`RANDOM}};
  sc_fail_r = _RAND_531[0:0];
  _RAND_532 = {1{`RANDOM}};
  probe_out_REG = _RAND_532[0:0];
  _RAND_533 = {9{`RANDOM}};
  probe_out_r = _RAND_533[273:0];
  _RAND_534 = {1{`RANDOM}};
  release_addr_aligned_REG = _RAND_534[8:0];
  _RAND_535 = {1{`RANDOM}};
  source = _RAND_535[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Uncache(
  input         clock,
  input         reset,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_opcode,
  output [2:0]  auto_out_a_bits_size,
  output [1:0]  auto_out_a_bits_source,
  output [31:0] auto_out_a_bits_address,
  output [7:0]  auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [63:0] auto_out_d_bits_data,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [38:0] io_in_req_bits_addr,
  input  [63:0] io_in_req_bits_wdata,
  input  [7:0]  io_in_req_bits_wmask,
  input         io_in_req_bits_wen,
  input  [1:0]  io_in_req_bits_len,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [63:0] io_in_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  _source_T = auto_out_a_ready & io_in_req_valid; // @[Decoupled.scala 51:35]
  reg [1:0] source; // @[Counter.scala 61:40]
  wire [1:0] _source_wrap_value_T_1 = source + 2'h1; // @[Counter.scala 77:24]
  wire [2:0] _get_bits_a_mask_sizeOH_T = {{1'd0}, io_in_req_bits_len}; // @[Misc.scala 201:34]
  wire [1:0] get_bits_a_mask_sizeOH_shiftAmount = _get_bits_a_mask_sizeOH_T[1:0]; // @[OneHot.scala 63:49]
  wire [3:0] _get_bits_a_mask_sizeOH_T_1 = 4'h1 << get_bits_a_mask_sizeOH_shiftAmount; // @[OneHot.scala 64:12]
  wire [2:0] get_bits_a_mask_sizeOH = _get_bits_a_mask_sizeOH_T_1[2:0] | 3'h1; // @[Misc.scala 201:81]
  wire  _get_bits_a_mask_T = io_in_req_bits_len >= 2'h3; // @[Misc.scala 205:21]
  wire  get_bits_a_mask_size = get_bits_a_mask_sizeOH[2]; // @[Misc.scala 208:26]
  wire  get_bits_a_mask_bit = io_in_req_bits_addr[2]; // @[Misc.scala 209:26]
  wire  get_bits_a_mask_nbit = ~get_bits_a_mask_bit; // @[Misc.scala 210:20]
  wire  get_bits_a_mask_acc = _get_bits_a_mask_T | get_bits_a_mask_size & get_bits_a_mask_nbit; // @[Misc.scala 214:29]
  wire  get_bits_a_mask_acc_1 = _get_bits_a_mask_T | get_bits_a_mask_size & get_bits_a_mask_bit; // @[Misc.scala 214:29]
  wire  get_bits_a_mask_size_1 = get_bits_a_mask_sizeOH[1]; // @[Misc.scala 208:26]
  wire  get_bits_a_mask_bit_1 = io_in_req_bits_addr[1]; // @[Misc.scala 209:26]
  wire  get_bits_a_mask_nbit_1 = ~get_bits_a_mask_bit_1; // @[Misc.scala 210:20]
  wire  get_bits_a_mask_eq_2 = get_bits_a_mask_nbit & get_bits_a_mask_nbit_1; // @[Misc.scala 213:27]
  wire  get_bits_a_mask_acc_2 = get_bits_a_mask_acc | get_bits_a_mask_size_1 & get_bits_a_mask_eq_2; // @[Misc.scala 214:29]
  wire  get_bits_a_mask_eq_3 = get_bits_a_mask_nbit & get_bits_a_mask_bit_1; // @[Misc.scala 213:27]
  wire  get_bits_a_mask_acc_3 = get_bits_a_mask_acc | get_bits_a_mask_size_1 & get_bits_a_mask_eq_3; // @[Misc.scala 214:29]
  wire  get_bits_a_mask_eq_4 = get_bits_a_mask_bit & get_bits_a_mask_nbit_1; // @[Misc.scala 213:27]
  wire  get_bits_a_mask_acc_4 = get_bits_a_mask_acc_1 | get_bits_a_mask_size_1 & get_bits_a_mask_eq_4; // @[Misc.scala 214:29]
  wire  get_bits_a_mask_eq_5 = get_bits_a_mask_bit & get_bits_a_mask_bit_1; // @[Misc.scala 213:27]
  wire  get_bits_a_mask_acc_5 = get_bits_a_mask_acc_1 | get_bits_a_mask_size_1 & get_bits_a_mask_eq_5; // @[Misc.scala 214:29]
  wire  get_bits_a_mask_size_2 = get_bits_a_mask_sizeOH[0]; // @[Misc.scala 208:26]
  wire  get_bits_a_mask_bit_2 = io_in_req_bits_addr[0]; // @[Misc.scala 209:26]
  wire  get_bits_a_mask_nbit_2 = ~get_bits_a_mask_bit_2; // @[Misc.scala 210:20]
  wire  get_bits_a_mask_eq_6 = get_bits_a_mask_eq_2 & get_bits_a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  get_bits_a_mask_acc_6 = get_bits_a_mask_acc_2 | get_bits_a_mask_size_2 & get_bits_a_mask_eq_6; // @[Misc.scala 214:29]
  wire  get_bits_a_mask_eq_7 = get_bits_a_mask_eq_2 & get_bits_a_mask_bit_2; // @[Misc.scala 213:27]
  wire  get_bits_a_mask_acc_7 = get_bits_a_mask_acc_2 | get_bits_a_mask_size_2 & get_bits_a_mask_eq_7; // @[Misc.scala 214:29]
  wire  get_bits_a_mask_eq_8 = get_bits_a_mask_eq_3 & get_bits_a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  get_bits_a_mask_acc_8 = get_bits_a_mask_acc_3 | get_bits_a_mask_size_2 & get_bits_a_mask_eq_8; // @[Misc.scala 214:29]
  wire  get_bits_a_mask_eq_9 = get_bits_a_mask_eq_3 & get_bits_a_mask_bit_2; // @[Misc.scala 213:27]
  wire  get_bits_a_mask_acc_9 = get_bits_a_mask_acc_3 | get_bits_a_mask_size_2 & get_bits_a_mask_eq_9; // @[Misc.scala 214:29]
  wire  get_bits_a_mask_eq_10 = get_bits_a_mask_eq_4 & get_bits_a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  get_bits_a_mask_acc_10 = get_bits_a_mask_acc_4 | get_bits_a_mask_size_2 & get_bits_a_mask_eq_10; // @[Misc.scala 214:29]
  wire  get_bits_a_mask_eq_11 = get_bits_a_mask_eq_4 & get_bits_a_mask_bit_2; // @[Misc.scala 213:27]
  wire  get_bits_a_mask_acc_11 = get_bits_a_mask_acc_4 | get_bits_a_mask_size_2 & get_bits_a_mask_eq_11; // @[Misc.scala 214:29]
  wire  get_bits_a_mask_eq_12 = get_bits_a_mask_eq_5 & get_bits_a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  get_bits_a_mask_acc_12 = get_bits_a_mask_acc_5 | get_bits_a_mask_size_2 & get_bits_a_mask_eq_12; // @[Misc.scala 214:29]
  wire  get_bits_a_mask_eq_13 = get_bits_a_mask_eq_5 & get_bits_a_mask_bit_2; // @[Misc.scala 213:27]
  wire  get_bits_a_mask_acc_13 = get_bits_a_mask_acc_5 | get_bits_a_mask_size_2 & get_bits_a_mask_eq_13; // @[Misc.scala 214:29]
  wire [7:0] get_bits_mask = {get_bits_a_mask_acc_13,get_bits_a_mask_acc_12,get_bits_a_mask_acc_11,
    get_bits_a_mask_acc_10,get_bits_a_mask_acc_9,get_bits_a_mask_acc_8,get_bits_a_mask_acc_7,get_bits_a_mask_acc_6}; // @[Cat.scala 33:92]
  wire [31:0] put_bits_address = io_in_req_bits_addr[31:0]; // @[Edges.scala 483:17 488:15]
  assign auto_out_a_valid = io_in_req_valid; // @[Nodes.scala 1212:84 Bus.scala 140:14]
  assign auto_out_a_bits_opcode = io_in_req_bits_wen ? 3'h1 : 3'h4; // @[Bus.scala 150:25]
  assign auto_out_a_bits_size = io_in_req_bits_wen ? _get_bits_a_mask_sizeOH_T : _get_bits_a_mask_sizeOH_T; // @[Bus.scala 150:25]
  assign auto_out_a_bits_source = source; // @[Bus.scala 150:25]
  assign auto_out_a_bits_address = io_in_req_bits_wen ? put_bits_address : put_bits_address; // @[Bus.scala 150:25]
  assign auto_out_a_bits_mask = io_in_req_bits_wen ? io_in_req_bits_wmask : get_bits_mask; // @[Bus.scala 150:25]
  assign auto_out_a_bits_data = io_in_req_bits_wen ? io_in_req_bits_wdata : 64'h0; // @[Bus.scala 150:25]
  assign auto_out_d_ready = io_in_resp_ready; // @[Nodes.scala 1212:84 Bus.scala 143:14]
  assign io_in_req_ready = auto_out_a_ready; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign io_in_resp_valid = auto_out_d_valid; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign io_in_resp_bits_rdata = auto_out_d_bits_data; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  always @(posedge clock) begin
    if (reset) begin // @[Counter.scala 61:40]
      source <= 2'h0; // @[Counter.scala 61:40]
    end else if (_source_T) begin // @[Counter.scala 118:16]
      source <= _source_wrap_value_T_1; // @[Counter.scala 77:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  source = _RAND_0[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLXbar(
  input          clock,
  input          reset,
  output         auto_in_2_a_ready,
  input          auto_in_2_a_valid,
  input  [1:0]   auto_in_2_a_bits_source,
  input  [31:0]  auto_in_2_a_bits_address,
  input          auto_in_2_b_ready,
  output         auto_in_2_b_valid,
  output [2:0]   auto_in_2_b_bits_size,
  output [1:0]   auto_in_2_b_bits_source,
  output [31:0]  auto_in_2_b_bits_address,
  output         auto_in_2_c_ready,
  input          auto_in_2_c_valid,
  input  [2:0]   auto_in_2_c_bits_opcode,
  input  [2:0]   auto_in_2_c_bits_param,
  input  [2:0]   auto_in_2_c_bits_size,
  input  [1:0]   auto_in_2_c_bits_source,
  input  [31:0]  auto_in_2_c_bits_address,
  input  [255:0] auto_in_2_c_bits_data,
  input          auto_in_2_d_ready,
  output         auto_in_2_d_valid,
  output [5:0]   auto_in_2_d_bits_sink,
  output [255:0] auto_in_2_d_bits_data,
  output         auto_in_2_e_ready,
  input          auto_in_2_e_valid,
  input  [5:0]   auto_in_2_e_bits_sink,
  output         auto_in_1_a_ready,
  input          auto_in_1_a_valid,
  input  [2:0]   auto_in_1_a_bits_opcode,
  input  [2:0]   auto_in_1_a_bits_size,
  input  [1:0]   auto_in_1_a_bits_source,
  input  [31:0]  auto_in_1_a_bits_address,
  input  [31:0]  auto_in_1_a_bits_mask,
  input  [255:0] auto_in_1_a_bits_data,
  input          auto_in_1_d_ready,
  output         auto_in_1_d_valid,
  output [2:0]   auto_in_1_d_bits_opcode,
  output [2:0]   auto_in_1_d_bits_size,
  output [1:0]   auto_in_1_d_bits_source,
  output [255:0] auto_in_1_d_bits_data,
  output         auto_in_0_a_ready,
  input          auto_in_0_a_valid,
  input  [1:0]   auto_in_0_a_bits_source,
  input  [31:0]  auto_in_0_a_bits_address,
  input          auto_in_0_d_ready,
  output         auto_in_0_d_valid,
  output [255:0] auto_in_0_d_bits_data,
  input          auto_out_a_ready,
  output         auto_out_a_valid,
  output [2:0]   auto_out_a_bits_opcode,
  output [2:0]   auto_out_a_bits_param,
  output [2:0]   auto_out_a_bits_size,
  output [3:0]   auto_out_a_bits_source,
  output [31:0]  auto_out_a_bits_address,
  output [31:0]  auto_out_a_bits_mask,
  output [255:0] auto_out_a_bits_data,
  output         auto_out_b_ready,
  input          auto_out_b_valid,
  input  [2:0]   auto_out_b_bits_size,
  input  [3:0]   auto_out_b_bits_source,
  input  [31:0]  auto_out_b_bits_address,
  input          auto_out_c_ready,
  output         auto_out_c_valid,
  output [2:0]   auto_out_c_bits_opcode,
  output [2:0]   auto_out_c_bits_param,
  output [2:0]   auto_out_c_bits_size,
  output [3:0]   auto_out_c_bits_source,
  output [31:0]  auto_out_c_bits_address,
  output [255:0] auto_out_c_bits_data,
  output         auto_out_d_ready,
  input          auto_out_d_valid,
  input  [2:0]   auto_out_d_bits_opcode,
  input  [2:0]   auto_out_d_bits_size,
  input  [3:0]   auto_out_d_bits_source,
  input  [5:0]   auto_out_d_bits_sink,
  input  [255:0] auto_out_d_bits_data,
  input          auto_out_e_ready,
  output         auto_out_e_valid,
  output [5:0]   auto_out_e_bits_sink
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire [3:0] _GEN_0 = {{2'd0}, auto_in_0_a_bits_source}; // @[Xbar.scala 240:55]
  wire [3:0] in_0_a_bits_source = _GEN_0 | 4'h8; // @[Xbar.scala 240:55]
  wire [2:0] _GEN_1 = {{1'd0}, auto_in_1_a_bits_source}; // @[Xbar.scala 240:55]
  wire [2:0] _in_1_a_bits_source_T = _GEN_1 | 3'h4; // @[Xbar.scala 240:55]
  wire  requestBOI_0_2 = auto_out_b_bits_source[3:2] == 2'h0; // @[Parameters.scala 54:32]
  wire  requestDOI_0_0 = auto_out_d_bits_source[3:2] == 2'h2; // @[Parameters.scala 54:32]
  wire  requestDOI_0_1 = auto_out_d_bits_source[3:2] == 2'h1; // @[Parameters.scala 54:32]
  wire  requestDOI_0_2 = auto_out_d_bits_source[3:2] == 2'h0; // @[Parameters.scala 54:32]
  reg  beatsLeft; // @[Arbiter.scala 88:30]
  wire  idle = ~beatsLeft; // @[Arbiter.scala 89:28]
  wire  latch = idle & auto_out_a_ready; // @[Arbiter.scala 90:24]
  wire [2:0] _readys_T = {auto_in_2_a_valid,auto_in_1_a_valid,auto_in_0_a_valid}; // @[Cat.scala 33:92]
  wire [2:0] _GEN_2 = {{1'd0}, _readys_T[2:1]}; // @[package.scala 254:43]
  wire [2:0] _readys_T_2 = _readys_T | _GEN_2; // @[package.scala 254:43]
  wire [2:0] _GEN_3 = {{2'd0}, _readys_T_2[2]}; // @[package.scala 254:43]
  wire [2:0] _readys_T_4 = _readys_T_2 | _GEN_3; // @[package.scala 254:43]
  wire [2:0] _readys_T_7 = {{1'd0}, _readys_T_4[2:1]}; // @[Arbiter.scala 19:90]
  wire [2:0] _readys_T_8 = ~_readys_T_7; // @[Arbiter.scala 19:62]
  wire  readys_0 = _readys_T_8[0]; // @[Arbiter.scala 96:86]
  wire  readys_1 = _readys_T_8[1]; // @[Arbiter.scala 96:86]
  wire  readys_2 = _readys_T_8[2]; // @[Arbiter.scala 96:86]
  wire  earlyWinner_0 = readys_0 & auto_in_0_a_valid; // @[Arbiter.scala 98:79]
  wire  earlyWinner_1 = readys_1 & auto_in_1_a_valid; // @[Arbiter.scala 98:79]
  wire  earlyWinner_2 = readys_2 & auto_in_2_a_valid; // @[Arbiter.scala 98:79]
  wire  prefixOR_2 = earlyWinner_0 | earlyWinner_1; // @[Arbiter.scala 105:53]
  wire  _prefixOR_T = prefixOR_2 | earlyWinner_2; // @[Arbiter.scala 105:53]
  wire  _T_13 = ~reset; // @[Arbiter.scala 106:13]
  wire  _T_16 = auto_in_0_a_valid | auto_in_1_a_valid | auto_in_2_a_valid; // @[Arbiter.scala 108:36]
  wire  _T_17 = ~(auto_in_0_a_valid | auto_in_1_a_valid | auto_in_2_a_valid); // @[Arbiter.scala 108:15]
  reg  state_0; // @[Arbiter.scala 117:26]
  wire  muxStateEarly_0 = idle ? earlyWinner_0 : state_0; // @[Arbiter.scala 118:30]
  reg  state_1; // @[Arbiter.scala 117:26]
  wire  muxStateEarly_1 = idle ? earlyWinner_1 : state_1; // @[Arbiter.scala 118:30]
  reg  state_2; // @[Arbiter.scala 117:26]
  wire  muxStateEarly_2 = idle ? earlyWinner_2 : state_2; // @[Arbiter.scala 118:30]
  wire  _out_0_a_earlyValid_T_6 = state_0 & auto_in_0_a_valid | state_1 & auto_in_1_a_valid | state_2 &
    auto_in_2_a_valid; // @[Mux.scala 27:73]
  wire  out_3_0_a_earlyValid = idle ? _T_16 : _out_0_a_earlyValid_T_6; // @[Arbiter.scala 126:29]
  wire  _beatsLeft_T_2 = auto_out_a_ready & out_3_0_a_earlyValid; // @[ReadyValidCancel.scala 49:33]
  wire  allowed_0 = idle ? readys_0 : state_0; // @[Arbiter.scala 122:24]
  wire  allowed_1 = idle ? readys_1 : state_1; // @[Arbiter.scala 122:24]
  wire  allowed_2 = idle ? readys_2 : state_2; // @[Arbiter.scala 122:24]
  wire [31:0] _T_43 = muxStateEarly_0 ? 32'hffffffff : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _T_44 = muxStateEarly_1 ? auto_in_1_a_bits_mask : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _T_45 = muxStateEarly_2 ? 32'hffffffff : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _T_46 = _T_43 | _T_44; // @[Mux.scala 27:73]
  wire [31:0] _T_48 = muxStateEarly_0 ? auto_in_0_a_bits_address : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _T_49 = muxStateEarly_1 ? auto_in_1_a_bits_address : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _T_50 = muxStateEarly_2 ? auto_in_2_a_bits_address : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _T_51 = _T_48 | _T_49; // @[Mux.scala 27:73]
  wire [3:0] _T_53 = muxStateEarly_0 ? in_0_a_bits_source : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] in_1_a_bits_source = {{1'd0}, _in_1_a_bits_source_T}; // @[Xbar.scala 234:18 240:29]
  wire [3:0] _T_54 = muxStateEarly_1 ? in_1_a_bits_source : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] in_2_a_bits_source = {{2'd0}, auto_in_2_a_bits_source}; // @[Xbar.scala 234:18 240:29]
  wire [3:0] _T_55 = muxStateEarly_2 ? in_2_a_bits_source : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_56 = _T_53 | _T_54; // @[Mux.scala 27:73]
  wire [2:0] _T_58 = muxStateEarly_0 ? 3'h5 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_59 = muxStateEarly_1 ? auto_in_1_a_bits_size : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_60 = muxStateEarly_2 ? 3'h5 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_61 = _T_58 | _T_59; // @[Mux.scala 27:73]
  wire [2:0] _T_68 = muxStateEarly_0 ? 3'h4 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_69 = muxStateEarly_1 ? auto_in_1_a_bits_opcode : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_70 = muxStateEarly_2 ? 3'h6 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_71 = _T_68 | _T_69; // @[Mux.scala 27:73]
  assign auto_in_2_a_ready = auto_out_a_ready & allowed_2; // @[Arbiter.scala 124:31]
  assign auto_in_2_b_valid = auto_out_b_valid & requestBOI_0_2; // @[Xbar.scala 182:40]
  assign auto_in_2_b_bits_size = auto_out_b_bits_size; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_2_b_bits_source = auto_out_b_bits_source[1:0]; // @[Xbar.scala 231:69]
  assign auto_in_2_b_bits_address = auto_out_b_bits_address; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_2_c_ready = auto_out_c_ready; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_2_d_valid = auto_out_d_valid & requestDOI_0_2; // @[Xbar.scala 182:40]
  assign auto_in_2_d_bits_sink = auto_out_d_bits_sink; // @[Xbar.scala 326:53]
  assign auto_in_2_d_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_2_e_ready = auto_out_e_ready; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_1_a_ready = auto_out_a_ready & allowed_1; // @[Arbiter.scala 124:31]
  assign auto_in_1_d_valid = auto_out_d_valid & requestDOI_0_1; // @[Xbar.scala 182:40]
  assign auto_in_1_d_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_1_d_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_1_d_bits_source = auto_out_d_bits_source[1:0]; // @[Xbar.scala 231:69]
  assign auto_in_1_d_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_0_a_ready = auto_out_a_ready & allowed_0; // @[Arbiter.scala 124:31]
  assign auto_in_0_d_valid = auto_out_d_valid & requestDOI_0_0; // @[Xbar.scala 182:40]
  assign auto_in_0_d_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_out_a_valid = idle ? _T_16 : _out_0_a_earlyValid_T_6; // @[Arbiter.scala 126:29]
  assign auto_out_a_bits_opcode = _T_71 | _T_70; // @[Mux.scala 27:73]
  assign auto_out_a_bits_param = muxStateEarly_2 ? 3'h1 : 3'h0; // @[Mux.scala 27:73]
  assign auto_out_a_bits_size = _T_61 | _T_60; // @[Mux.scala 27:73]
  assign auto_out_a_bits_source = _T_56 | _T_55; // @[Mux.scala 27:73]
  assign auto_out_a_bits_address = _T_51 | _T_50; // @[Mux.scala 27:73]
  assign auto_out_a_bits_mask = _T_46 | _T_45; // @[Mux.scala 27:73]
  assign auto_out_a_bits_data = muxStateEarly_1 ? auto_in_1_a_bits_data : 256'h0; // @[Mux.scala 27:73]
  assign auto_out_b_ready = requestBOI_0_2 & auto_in_2_b_ready; // @[Mux.scala 27:73]
  assign auto_out_c_valid = auto_in_2_c_valid; // @[ReadyValidCancel.scala 21:38]
  assign auto_out_c_bits_opcode = auto_in_2_c_bits_opcode; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_c_bits_param = auto_in_2_c_bits_param; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_c_bits_size = auto_in_2_c_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_c_bits_source = {{2'd0}, auto_in_2_c_bits_source}; // @[Xbar.scala 234:18 262:29]
  assign auto_out_c_bits_address = auto_in_2_c_bits_address; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_c_bits_data = auto_in_2_c_bits_data; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_d_ready = requestDOI_0_0 & auto_in_0_d_ready | requestDOI_0_1 & auto_in_1_d_ready | requestDOI_0_2 &
    auto_in_2_d_ready; // @[Mux.scala 27:73]
  assign auto_out_e_valid = auto_in_2_e_valid; // @[ReadyValidCancel.scala 21:38]
  assign auto_out_e_bits_sink = auto_in_2_e_bits_sink; // @[Xbar.scala 231:69]
  always @(posedge clock) begin
    if (reset) begin // @[Arbiter.scala 88:30]
      beatsLeft <= 1'h0; // @[Arbiter.scala 88:30]
    end else if (latch) begin // @[Arbiter.scala 114:23]
      beatsLeft <= 1'h0;
    end else begin
      beatsLeft <= beatsLeft - _beatsLeft_T_2;
    end
    if (reset) begin // @[Arbiter.scala 117:26]
      state_0 <= 1'h0; // @[Arbiter.scala 117:26]
    end else if (idle) begin // @[Arbiter.scala 118:30]
      state_0 <= earlyWinner_0;
    end
    if (reset) begin // @[Arbiter.scala 117:26]
      state_1 <= 1'h0; // @[Arbiter.scala 117:26]
    end else if (idle) begin // @[Arbiter.scala 118:30]
      state_1 <= earlyWinner_1;
    end
    if (reset) begin // @[Arbiter.scala 117:26]
      state_2 <= 1'h0; // @[Arbiter.scala 117:26]
    end else if (idle) begin // @[Arbiter.scala 118:30]
      state_2 <= earlyWinner_2;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~((~earlyWinner_0 | ~earlyWinner_1) & (~prefixOR_2 | ~earlyWinner_2))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:106 assert((prefixOR zip earlyWinner) map { case (p,w) => !p || !w } reduce {_ && _})\n"
            ); // @[Arbiter.scala 106:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~((~earlyWinner_0 | ~earlyWinner_1) & (~prefixOR_2 | ~earlyWinner_2))) begin
          $fatal; // @[Arbiter.scala 106:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & ~(~(auto_in_0_a_valid | auto_in_1_a_valid | auto_in_2_a_valid) | _prefixOR_T)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:108 assert (!earlyValids.reduce(_||_) || earlyWinner.reduce(_||_))\n"
            ); // @[Arbiter.scala 108:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_13 & ~(~(auto_in_0_a_valid | auto_in_1_a_valid | auto_in_2_a_valid) | _prefixOR_T)) begin
          $fatal; // @[Arbiter.scala 108:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & ~(_T_17 | _T_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:109 assert (!validQuals .reduce(_||_) || validQuals .reduce(_||_))\n"
            ); // @[Arbiter.scala 109:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_13 & ~(_T_17 | _T_16)) begin
          $fatal; // @[Arbiter.scala 109:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  beatsLeft = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  state_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  state_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  state_2 = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Repeater(
  input          clock,
  input          reset,
  input          io_repeat,
  output         io_enq_ready,
  input          io_enq_valid,
  input  [2:0]   io_enq_bits_opcode,
  input  [2:0]   io_enq_bits_size,
  input  [1:0]   io_enq_bits_source,
  input  [255:0] io_enq_bits_data,
  input          io_deq_ready,
  output         io_deq_valid,
  output [2:0]   io_deq_bits_opcode,
  output [2:0]   io_deq_bits_size,
  output [1:0]   io_deq_bits_source,
  output [255:0] io_deq_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [255:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg  full; // @[Repeater.scala 19:21]
  reg [2:0] saved_opcode; // @[Repeater.scala 20:18]
  reg [2:0] saved_size; // @[Repeater.scala 20:18]
  reg [1:0] saved_source; // @[Repeater.scala 20:18]
  reg [255:0] saved_data; // @[Repeater.scala 20:18]
  wire  _T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  _GEN_0 = _T & io_repeat | full; // @[Repeater.scala 19:21 28:{38,45}]
  wire  _T_2 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  assign io_enq_ready = io_deq_ready & ~full; // @[Repeater.scala 24:32]
  assign io_deq_valid = io_enq_valid | full; // @[Repeater.scala 23:32]
  assign io_deq_bits_opcode = full ? saved_opcode : io_enq_bits_opcode; // @[Repeater.scala 25:21]
  assign io_deq_bits_size = full ? saved_size : io_enq_bits_size; // @[Repeater.scala 25:21]
  assign io_deq_bits_source = full ? saved_source : io_enq_bits_source; // @[Repeater.scala 25:21]
  assign io_deq_bits_data = full ? saved_data : io_enq_bits_data; // @[Repeater.scala 25:21]
  always @(posedge clock) begin
    if (reset) begin // @[Repeater.scala 19:21]
      full <= 1'h0; // @[Repeater.scala 19:21]
    end else if (_T_2 & ~io_repeat) begin // @[Repeater.scala 29:38]
      full <= 1'h0; // @[Repeater.scala 29:45]
    end else begin
      full <= _GEN_0;
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_opcode <= io_enq_bits_opcode; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_size <= io_enq_bits_size; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_source <= io_enq_bits_source; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_data <= io_enq_bits_data; // @[Repeater.scala 28:62]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  full = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  saved_opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  saved_size = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  saved_source = _RAND_3[1:0];
  _RAND_4 = {8{`RANDOM}};
  saved_data = _RAND_4[255:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLWidthWidget(
  input          clock,
  input          reset,
  output         auto_in_a_ready,
  input          auto_in_a_valid,
  input  [2:0]   auto_in_a_bits_opcode,
  input  [2:0]   auto_in_a_bits_size,
  input  [1:0]   auto_in_a_bits_source,
  input  [31:0]  auto_in_a_bits_address,
  input  [7:0]   auto_in_a_bits_mask,
  input  [63:0]  auto_in_a_bits_data,
  input          auto_in_d_ready,
  output         auto_in_d_valid,
  output [63:0]  auto_in_d_bits_data,
  input          auto_out_a_ready,
  output         auto_out_a_valid,
  output [2:0]   auto_out_a_bits_opcode,
  output [2:0]   auto_out_a_bits_size,
  output [1:0]   auto_out_a_bits_source,
  output [31:0]  auto_out_a_bits_address,
  output [31:0]  auto_out_a_bits_mask,
  output [255:0] auto_out_a_bits_data,
  output         auto_out_d_ready,
  input          auto_out_d_valid,
  input  [2:0]   auto_out_d_bits_opcode,
  input  [2:0]   auto_out_d_bits_size,
  input  [1:0]   auto_out_d_bits_source,
  input  [255:0] auto_out_d_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
`endif // RANDOMIZE_REG_INIT
  wire  repeated_repeater_clock; // @[Repeater.scala 35:26]
  wire  repeated_repeater_reset; // @[Repeater.scala 35:26]
  wire  repeated_repeater_io_repeat; // @[Repeater.scala 35:26]
  wire  repeated_repeater_io_enq_ready; // @[Repeater.scala 35:26]
  wire  repeated_repeater_io_enq_valid; // @[Repeater.scala 35:26]
  wire [2:0] repeated_repeater_io_enq_bits_opcode; // @[Repeater.scala 35:26]
  wire [2:0] repeated_repeater_io_enq_bits_size; // @[Repeater.scala 35:26]
  wire [1:0] repeated_repeater_io_enq_bits_source; // @[Repeater.scala 35:26]
  wire [255:0] repeated_repeater_io_enq_bits_data; // @[Repeater.scala 35:26]
  wire  repeated_repeater_io_deq_ready; // @[Repeater.scala 35:26]
  wire  repeated_repeater_io_deq_valid; // @[Repeater.scala 35:26]
  wire [2:0] repeated_repeater_io_deq_bits_opcode; // @[Repeater.scala 35:26]
  wire [2:0] repeated_repeater_io_deq_bits_size; // @[Repeater.scala 35:26]
  wire [1:0] repeated_repeater_io_deq_bits_source; // @[Repeater.scala 35:26]
  wire [255:0] repeated_repeater_io_deq_bits_data; // @[Repeater.scala 35:26]
  wire  hasData = ~auto_in_a_bits_opcode[2]; // @[Edges.scala 91:28]
  wire [11:0] _limit_T_1 = 12'h1f << auto_in_a_bits_size; // @[package.scala 235:71]
  wire [4:0] _limit_T_3 = ~_limit_T_1[4:0]; // @[package.scala 235:46]
  wire [1:0] limit = _limit_T_3[4:3]; // @[WidthWidget.scala 33:47]
  reg [1:0] count; // @[WidthWidget.scala 35:27]
  wire  last = count == limit | ~hasData; // @[WidthWidget.scala 37:36]
  wire [1:0] _enable_T_1 = count & limit; // @[WidthWidget.scala 38:63]
  wire  enable_0 = ~(|_enable_T_1); // @[WidthWidget.scala 38:47]
  wire [1:0] _enable_T_3 = count ^ 2'h1; // @[WidthWidget.scala 38:56]
  wire [1:0] _enable_T_4 = _enable_T_3 & limit; // @[WidthWidget.scala 38:63]
  wire  enable_1 = ~(|_enable_T_4); // @[WidthWidget.scala 38:47]
  wire [1:0] _enable_T_6 = count ^ 2'h2; // @[WidthWidget.scala 38:56]
  wire [1:0] _enable_T_7 = _enable_T_6 & limit; // @[WidthWidget.scala 38:63]
  wire  enable_2 = ~(|_enable_T_7); // @[WidthWidget.scala 38:47]
  wire  _bundleIn_0_a_ready_T = ~last; // @[WidthWidget.scala 71:32]
  wire  bundleIn_0_a_ready = auto_out_a_ready | ~last; // @[WidthWidget.scala 71:29]
  wire  _T = bundleIn_0_a_ready & auto_in_a_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _count_T_1 = count + 2'h1; // @[WidthWidget.scala 45:24]
  reg  x1_a_bits_data_rdata_written_once; // @[WidthWidget.scala 57:41]
  wire  x1_a_bits_data_masked_enable_0 = enable_0 | ~x1_a_bits_data_rdata_written_once; // @[WidthWidget.scala 58:42]
  wire  x1_a_bits_data_masked_enable_1 = enable_1 | ~x1_a_bits_data_rdata_written_once; // @[WidthWidget.scala 58:42]
  wire  x1_a_bits_data_masked_enable_2 = enable_2 | ~x1_a_bits_data_rdata_written_once; // @[WidthWidget.scala 58:42]
  reg [63:0] x1_a_bits_data_rdata_0; // @[WidthWidget.scala 61:24]
  reg [63:0] x1_a_bits_data_rdata_1; // @[WidthWidget.scala 61:24]
  reg [63:0] x1_a_bits_data_rdata_2; // @[WidthWidget.scala 61:24]
  wire [63:0] x1_a_bits_data_mdata_0 = x1_a_bits_data_masked_enable_0 ? auto_in_a_bits_data : x1_a_bits_data_rdata_0; // @[WidthWidget.scala 63:88]
  wire [63:0] x1_a_bits_data_mdata_1 = x1_a_bits_data_masked_enable_1 ? auto_in_a_bits_data : x1_a_bits_data_rdata_1; // @[WidthWidget.scala 63:88]
  wire [63:0] x1_a_bits_data_mdata_2 = x1_a_bits_data_masked_enable_2 ? auto_in_a_bits_data : x1_a_bits_data_rdata_2; // @[WidthWidget.scala 63:88]
  wire  _GEN_4 = _T & _bundleIn_0_a_ready_T | x1_a_bits_data_rdata_written_once; // @[WidthWidget.scala 64:35 65:30 57:41]
  wire [127:0] x1_a_bits_data_lo = {x1_a_bits_data_mdata_1,x1_a_bits_data_mdata_0}; // @[Cat.scala 33:92]
  wire [127:0] x1_a_bits_data_hi = {auto_in_a_bits_data,x1_a_bits_data_mdata_2}; // @[Cat.scala 33:92]
  wire [4:0] _x1_a_bits_mask_sizeOH_T = {{2'd0}, auto_in_a_bits_size}; // @[Misc.scala 201:34]
  wire [2:0] x1_a_bits_mask_sizeOH_shiftAmount = _x1_a_bits_mask_sizeOH_T[2:0]; // @[OneHot.scala 63:49]
  wire [7:0] _x1_a_bits_mask_sizeOH_T_1 = 8'h1 << x1_a_bits_mask_sizeOH_shiftAmount; // @[OneHot.scala 64:12]
  wire [4:0] x1_a_bits_mask_sizeOH = _x1_a_bits_mask_sizeOH_T_1[4:0] | 5'h1; // @[Misc.scala 201:81]
  wire  _x1_a_bits_mask_T = auto_in_a_bits_size >= 3'h5; // @[Misc.scala 205:21]
  wire  x1_a_bits_mask_size = x1_a_bits_mask_sizeOH[4]; // @[Misc.scala 208:26]
  wire  x1_a_bits_mask_bit = auto_in_a_bits_address[4]; // @[Misc.scala 209:26]
  wire  x1_a_bits_mask_nbit = ~x1_a_bits_mask_bit; // @[Misc.scala 210:20]
  wire  x1_a_bits_mask_acc = _x1_a_bits_mask_T | x1_a_bits_mask_size & x1_a_bits_mask_nbit; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_acc_1 = _x1_a_bits_mask_T | x1_a_bits_mask_size & x1_a_bits_mask_bit; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_size_1 = x1_a_bits_mask_sizeOH[3]; // @[Misc.scala 208:26]
  wire  x1_a_bits_mask_bit_1 = auto_in_a_bits_address[3]; // @[Misc.scala 209:26]
  wire  x1_a_bits_mask_nbit_1 = ~x1_a_bits_mask_bit_1; // @[Misc.scala 210:20]
  wire  x1_a_bits_mask_eq_2 = x1_a_bits_mask_nbit & x1_a_bits_mask_nbit_1; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_2 = x1_a_bits_mask_acc | x1_a_bits_mask_size_1 & x1_a_bits_mask_eq_2; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_3 = x1_a_bits_mask_nbit & x1_a_bits_mask_bit_1; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_3 = x1_a_bits_mask_acc | x1_a_bits_mask_size_1 & x1_a_bits_mask_eq_3; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_4 = x1_a_bits_mask_bit & x1_a_bits_mask_nbit_1; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_4 = x1_a_bits_mask_acc_1 | x1_a_bits_mask_size_1 & x1_a_bits_mask_eq_4; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_5 = x1_a_bits_mask_bit & x1_a_bits_mask_bit_1; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_5 = x1_a_bits_mask_acc_1 | x1_a_bits_mask_size_1 & x1_a_bits_mask_eq_5; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_size_2 = x1_a_bits_mask_sizeOH[2]; // @[Misc.scala 208:26]
  wire  x1_a_bits_mask_bit_2 = auto_in_a_bits_address[2]; // @[Misc.scala 209:26]
  wire  x1_a_bits_mask_nbit_2 = ~x1_a_bits_mask_bit_2; // @[Misc.scala 210:20]
  wire  x1_a_bits_mask_eq_6 = x1_a_bits_mask_eq_2 & x1_a_bits_mask_nbit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_6 = x1_a_bits_mask_acc_2 | x1_a_bits_mask_size_2 & x1_a_bits_mask_eq_6; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_7 = x1_a_bits_mask_eq_2 & x1_a_bits_mask_bit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_7 = x1_a_bits_mask_acc_2 | x1_a_bits_mask_size_2 & x1_a_bits_mask_eq_7; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_8 = x1_a_bits_mask_eq_3 & x1_a_bits_mask_nbit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_8 = x1_a_bits_mask_acc_3 | x1_a_bits_mask_size_2 & x1_a_bits_mask_eq_8; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_9 = x1_a_bits_mask_eq_3 & x1_a_bits_mask_bit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_9 = x1_a_bits_mask_acc_3 | x1_a_bits_mask_size_2 & x1_a_bits_mask_eq_9; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_10 = x1_a_bits_mask_eq_4 & x1_a_bits_mask_nbit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_10 = x1_a_bits_mask_acc_4 | x1_a_bits_mask_size_2 & x1_a_bits_mask_eq_10; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_11 = x1_a_bits_mask_eq_4 & x1_a_bits_mask_bit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_11 = x1_a_bits_mask_acc_4 | x1_a_bits_mask_size_2 & x1_a_bits_mask_eq_11; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_12 = x1_a_bits_mask_eq_5 & x1_a_bits_mask_nbit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_12 = x1_a_bits_mask_acc_5 | x1_a_bits_mask_size_2 & x1_a_bits_mask_eq_12; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_13 = x1_a_bits_mask_eq_5 & x1_a_bits_mask_bit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_13 = x1_a_bits_mask_acc_5 | x1_a_bits_mask_size_2 & x1_a_bits_mask_eq_13; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_size_3 = x1_a_bits_mask_sizeOH[1]; // @[Misc.scala 208:26]
  wire  x1_a_bits_mask_bit_3 = auto_in_a_bits_address[1]; // @[Misc.scala 209:26]
  wire  x1_a_bits_mask_nbit_3 = ~x1_a_bits_mask_bit_3; // @[Misc.scala 210:20]
  wire  x1_a_bits_mask_eq_14 = x1_a_bits_mask_eq_6 & x1_a_bits_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_14 = x1_a_bits_mask_acc_6 | x1_a_bits_mask_size_3 & x1_a_bits_mask_eq_14; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_15 = x1_a_bits_mask_eq_6 & x1_a_bits_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_15 = x1_a_bits_mask_acc_6 | x1_a_bits_mask_size_3 & x1_a_bits_mask_eq_15; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_16 = x1_a_bits_mask_eq_7 & x1_a_bits_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_16 = x1_a_bits_mask_acc_7 | x1_a_bits_mask_size_3 & x1_a_bits_mask_eq_16; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_17 = x1_a_bits_mask_eq_7 & x1_a_bits_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_17 = x1_a_bits_mask_acc_7 | x1_a_bits_mask_size_3 & x1_a_bits_mask_eq_17; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_18 = x1_a_bits_mask_eq_8 & x1_a_bits_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_18 = x1_a_bits_mask_acc_8 | x1_a_bits_mask_size_3 & x1_a_bits_mask_eq_18; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_19 = x1_a_bits_mask_eq_8 & x1_a_bits_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_19 = x1_a_bits_mask_acc_8 | x1_a_bits_mask_size_3 & x1_a_bits_mask_eq_19; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_20 = x1_a_bits_mask_eq_9 & x1_a_bits_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_20 = x1_a_bits_mask_acc_9 | x1_a_bits_mask_size_3 & x1_a_bits_mask_eq_20; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_21 = x1_a_bits_mask_eq_9 & x1_a_bits_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_21 = x1_a_bits_mask_acc_9 | x1_a_bits_mask_size_3 & x1_a_bits_mask_eq_21; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_22 = x1_a_bits_mask_eq_10 & x1_a_bits_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_22 = x1_a_bits_mask_acc_10 | x1_a_bits_mask_size_3 & x1_a_bits_mask_eq_22; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_23 = x1_a_bits_mask_eq_10 & x1_a_bits_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_23 = x1_a_bits_mask_acc_10 | x1_a_bits_mask_size_3 & x1_a_bits_mask_eq_23; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_24 = x1_a_bits_mask_eq_11 & x1_a_bits_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_24 = x1_a_bits_mask_acc_11 | x1_a_bits_mask_size_3 & x1_a_bits_mask_eq_24; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_25 = x1_a_bits_mask_eq_11 & x1_a_bits_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_25 = x1_a_bits_mask_acc_11 | x1_a_bits_mask_size_3 & x1_a_bits_mask_eq_25; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_26 = x1_a_bits_mask_eq_12 & x1_a_bits_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_26 = x1_a_bits_mask_acc_12 | x1_a_bits_mask_size_3 & x1_a_bits_mask_eq_26; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_27 = x1_a_bits_mask_eq_12 & x1_a_bits_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_27 = x1_a_bits_mask_acc_12 | x1_a_bits_mask_size_3 & x1_a_bits_mask_eq_27; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_28 = x1_a_bits_mask_eq_13 & x1_a_bits_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_28 = x1_a_bits_mask_acc_13 | x1_a_bits_mask_size_3 & x1_a_bits_mask_eq_28; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_29 = x1_a_bits_mask_eq_13 & x1_a_bits_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_29 = x1_a_bits_mask_acc_13 | x1_a_bits_mask_size_3 & x1_a_bits_mask_eq_29; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_size_4 = x1_a_bits_mask_sizeOH[0]; // @[Misc.scala 208:26]
  wire  x1_a_bits_mask_bit_4 = auto_in_a_bits_address[0]; // @[Misc.scala 209:26]
  wire  x1_a_bits_mask_nbit_4 = ~x1_a_bits_mask_bit_4; // @[Misc.scala 210:20]
  wire  x1_a_bits_mask_eq_30 = x1_a_bits_mask_eq_14 & x1_a_bits_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_30 = x1_a_bits_mask_acc_14 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_30; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_31 = x1_a_bits_mask_eq_14 & x1_a_bits_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_31 = x1_a_bits_mask_acc_14 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_31; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_32 = x1_a_bits_mask_eq_15 & x1_a_bits_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_32 = x1_a_bits_mask_acc_15 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_32; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_33 = x1_a_bits_mask_eq_15 & x1_a_bits_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_33 = x1_a_bits_mask_acc_15 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_33; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_34 = x1_a_bits_mask_eq_16 & x1_a_bits_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_34 = x1_a_bits_mask_acc_16 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_34; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_35 = x1_a_bits_mask_eq_16 & x1_a_bits_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_35 = x1_a_bits_mask_acc_16 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_35; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_36 = x1_a_bits_mask_eq_17 & x1_a_bits_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_36 = x1_a_bits_mask_acc_17 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_36; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_37 = x1_a_bits_mask_eq_17 & x1_a_bits_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_37 = x1_a_bits_mask_acc_17 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_37; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_38 = x1_a_bits_mask_eq_18 & x1_a_bits_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_38 = x1_a_bits_mask_acc_18 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_38; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_39 = x1_a_bits_mask_eq_18 & x1_a_bits_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_39 = x1_a_bits_mask_acc_18 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_39; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_40 = x1_a_bits_mask_eq_19 & x1_a_bits_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_40 = x1_a_bits_mask_acc_19 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_40; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_41 = x1_a_bits_mask_eq_19 & x1_a_bits_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_41 = x1_a_bits_mask_acc_19 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_41; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_42 = x1_a_bits_mask_eq_20 & x1_a_bits_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_42 = x1_a_bits_mask_acc_20 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_42; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_43 = x1_a_bits_mask_eq_20 & x1_a_bits_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_43 = x1_a_bits_mask_acc_20 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_43; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_44 = x1_a_bits_mask_eq_21 & x1_a_bits_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_44 = x1_a_bits_mask_acc_21 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_44; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_45 = x1_a_bits_mask_eq_21 & x1_a_bits_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_45 = x1_a_bits_mask_acc_21 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_45; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_46 = x1_a_bits_mask_eq_22 & x1_a_bits_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_46 = x1_a_bits_mask_acc_22 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_46; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_47 = x1_a_bits_mask_eq_22 & x1_a_bits_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_47 = x1_a_bits_mask_acc_22 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_47; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_48 = x1_a_bits_mask_eq_23 & x1_a_bits_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_48 = x1_a_bits_mask_acc_23 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_48; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_49 = x1_a_bits_mask_eq_23 & x1_a_bits_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_49 = x1_a_bits_mask_acc_23 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_49; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_50 = x1_a_bits_mask_eq_24 & x1_a_bits_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_50 = x1_a_bits_mask_acc_24 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_50; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_51 = x1_a_bits_mask_eq_24 & x1_a_bits_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_51 = x1_a_bits_mask_acc_24 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_51; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_52 = x1_a_bits_mask_eq_25 & x1_a_bits_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_52 = x1_a_bits_mask_acc_25 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_52; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_53 = x1_a_bits_mask_eq_25 & x1_a_bits_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_53 = x1_a_bits_mask_acc_25 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_53; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_54 = x1_a_bits_mask_eq_26 & x1_a_bits_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_54 = x1_a_bits_mask_acc_26 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_54; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_55 = x1_a_bits_mask_eq_26 & x1_a_bits_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_55 = x1_a_bits_mask_acc_26 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_55; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_56 = x1_a_bits_mask_eq_27 & x1_a_bits_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_56 = x1_a_bits_mask_acc_27 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_56; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_57 = x1_a_bits_mask_eq_27 & x1_a_bits_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_57 = x1_a_bits_mask_acc_27 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_57; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_58 = x1_a_bits_mask_eq_28 & x1_a_bits_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_58 = x1_a_bits_mask_acc_28 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_58; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_59 = x1_a_bits_mask_eq_28 & x1_a_bits_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_59 = x1_a_bits_mask_acc_28 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_59; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_60 = x1_a_bits_mask_eq_29 & x1_a_bits_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_60 = x1_a_bits_mask_acc_29 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_60; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_61 = x1_a_bits_mask_eq_29 & x1_a_bits_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_61 = x1_a_bits_mask_acc_29 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_61; // @[Misc.scala 214:29]
  wire [7:0] x1_a_bits_mask_lo_lo = {x1_a_bits_mask_acc_37,x1_a_bits_mask_acc_36,x1_a_bits_mask_acc_35,
    x1_a_bits_mask_acc_34,x1_a_bits_mask_acc_33,x1_a_bits_mask_acc_32,x1_a_bits_mask_acc_31,x1_a_bits_mask_acc_30}; // @[Cat.scala 33:92]
  wire [15:0] x1_a_bits_mask_lo = {x1_a_bits_mask_acc_45,x1_a_bits_mask_acc_44,x1_a_bits_mask_acc_43,
    x1_a_bits_mask_acc_42,x1_a_bits_mask_acc_41,x1_a_bits_mask_acc_40,x1_a_bits_mask_acc_39,x1_a_bits_mask_acc_38,
    x1_a_bits_mask_lo_lo}; // @[Cat.scala 33:92]
  wire [7:0] x1_a_bits_mask_hi_lo = {x1_a_bits_mask_acc_53,x1_a_bits_mask_acc_52,x1_a_bits_mask_acc_51,
    x1_a_bits_mask_acc_50,x1_a_bits_mask_acc_49,x1_a_bits_mask_acc_48,x1_a_bits_mask_acc_47,x1_a_bits_mask_acc_46}; // @[Cat.scala 33:92]
  wire [31:0] _x1_a_bits_mask_T_1 = {x1_a_bits_mask_acc_61,x1_a_bits_mask_acc_60,x1_a_bits_mask_acc_59,
    x1_a_bits_mask_acc_58,x1_a_bits_mask_acc_57,x1_a_bits_mask_acc_56,x1_a_bits_mask_acc_55,x1_a_bits_mask_acc_54,
    x1_a_bits_mask_hi_lo,x1_a_bits_mask_lo}; // @[Cat.scala 33:92]
  reg  x1_a_bits_mask_rdata_written_once; // @[WidthWidget.scala 57:41]
  wire  x1_a_bits_mask_masked_enable_0 = enable_0 | ~x1_a_bits_mask_rdata_written_once; // @[WidthWidget.scala 58:42]
  wire  x1_a_bits_mask_masked_enable_1 = enable_1 | ~x1_a_bits_mask_rdata_written_once; // @[WidthWidget.scala 58:42]
  wire  x1_a_bits_mask_masked_enable_2 = enable_2 | ~x1_a_bits_mask_rdata_written_once; // @[WidthWidget.scala 58:42]
  reg [7:0] x1_a_bits_mask_rdata_0; // @[WidthWidget.scala 61:24]
  reg [7:0] x1_a_bits_mask_rdata_1; // @[WidthWidget.scala 61:24]
  reg [7:0] x1_a_bits_mask_rdata_2; // @[WidthWidget.scala 61:24]
  wire [7:0] x1_a_bits_mask_mdata_0 = x1_a_bits_mask_masked_enable_0 ? auto_in_a_bits_mask : x1_a_bits_mask_rdata_0; // @[WidthWidget.scala 63:88]
  wire [7:0] x1_a_bits_mask_mdata_1 = x1_a_bits_mask_masked_enable_1 ? auto_in_a_bits_mask : x1_a_bits_mask_rdata_1; // @[WidthWidget.scala 63:88]
  wire [7:0] x1_a_bits_mask_mdata_2 = x1_a_bits_mask_masked_enable_2 ? auto_in_a_bits_mask : x1_a_bits_mask_rdata_2; // @[WidthWidget.scala 63:88]
  wire  _GEN_8 = _T & _bundleIn_0_a_ready_T | x1_a_bits_mask_rdata_written_once; // @[WidthWidget.scala 64:35 65:30 57:41]
  wire [31:0] _x1_a_bits_mask_T_5 = {auto_in_a_bits_mask,x1_a_bits_mask_mdata_2,x1_a_bits_mask_mdata_1,
    x1_a_bits_mask_mdata_0}; // @[Cat.scala 33:92]
  wire [31:0] _x1_a_bits_mask_T_7 = hasData ? _x1_a_bits_mask_T_5 : 32'hffffffff; // @[WidthWidget.scala 80:93]
  wire [255:0] cated_bits_data = {repeated_repeater_io_deq_bits_data[255:64],auto_out_d_bits_data[63:0]}; // @[Cat.scala 33:92]
  wire [2:0] cated_bits_opcode = repeated_repeater_io_deq_bits_opcode; // @[WidthWidget.scala 156:25 157:15]
  wire  repeat_hasData = cated_bits_opcode[0]; // @[Edges.scala 105:36]
  wire [2:0] cated_bits_size = repeated_repeater_io_deq_bits_size; // @[WidthWidget.scala 156:25 157:15]
  wire [11:0] _repeat_limit_T_1 = 12'h1f << cated_bits_size; // @[package.scala 235:71]
  wire [4:0] _repeat_limit_T_3 = ~_repeat_limit_T_1[4:0]; // @[package.scala 235:46]
  wire [1:0] repeat_limit = _repeat_limit_T_3[4:3]; // @[WidthWidget.scala 98:47]
  reg [1:0] repeat_count; // @[WidthWidget.scala 100:26]
  wire  repeat_first = repeat_count == 2'h0; // @[WidthWidget.scala 101:25]
  wire  repeat_last = repeat_count == repeat_limit | ~repeat_hasData; // @[WidthWidget.scala 102:35]
  wire  cated_valid = repeated_repeater_io_deq_valid; // @[WidthWidget.scala 156:25 157:15]
  wire  _repeat_T = auto_in_d_ready & cated_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _repeat_count_T_1 = repeat_count + 2'h1; // @[WidthWidget.scala 105:24]
  reg [1:0] repeat_sel_sel_sources_0; // @[WidthWidget.scala 181:27]
  reg [1:0] repeat_sel_sel_sources_1; // @[WidthWidget.scala 181:27]
  reg [1:0] repeat_sel_sel_sources_2; // @[WidthWidget.scala 181:27]
  reg [1:0] repeat_sel_sel_sources_3; // @[WidthWidget.scala 181:27]
  wire [1:0] repeat_sel_sel_a_sel = auto_in_a_bits_address[4:3]; // @[WidthWidget.scala 182:38]
  wire [1:0] cated_bits_source = repeated_repeater_io_deq_bits_source; // @[WidthWidget.scala 156:25 157:15]
  wire  repeat_sel_sel_bypass = auto_in_a_valid & auto_in_a_bits_source == cated_bits_source; // @[WidthWidget.scala 190:33]
  wire [1:0] _GEN_23 = 2'h1 == cated_bits_source ? repeat_sel_sel_sources_1 : repeat_sel_sel_sources_0; // @[WidthWidget.scala 192:{17,17}]
  wire [1:0] _GEN_24 = 2'h2 == cated_bits_source ? repeat_sel_sel_sources_2 : _GEN_23; // @[WidthWidget.scala 192:{17,17}]
  wire [1:0] _GEN_25 = 2'h3 == cated_bits_source ? repeat_sel_sel_sources_3 : _GEN_24; // @[WidthWidget.scala 192:{17,17}]
  wire [1:0] repeat_sel_sel = repeat_sel_sel_bypass ? repeat_sel_sel_a_sel : _GEN_25; // @[WidthWidget.scala 192:17]
  reg [1:0] repeat_sel_hold_r; // @[Reg.scala 19:16]
  wire [1:0] _GEN_26 = repeat_first ? repeat_sel_sel : repeat_sel_hold_r; // @[Reg.scala 19:16 20:{18,22}]
  wire [1:0] _repeat_sel_T = ~repeat_limit; // @[WidthWidget.scala 117:18]
  wire [1:0] repeat_sel = _GEN_26 & _repeat_sel_T; // @[WidthWidget.scala 117:16]
  wire [1:0] repeat_index = repeat_sel | repeat_count; // @[WidthWidget.scala 121:24]
  wire [63:0] repeat_bundleIn_0_d_bits_data_mux_0 = cated_bits_data[63:0]; // @[WidthWidget.scala 123:55]
  wire [63:0] repeat_bundleIn_0_d_bits_data_mux_1 = cated_bits_data[127:64]; // @[WidthWidget.scala 123:55]
  wire [63:0] repeat_bundleIn_0_d_bits_data_mux_2 = cated_bits_data[191:128]; // @[WidthWidget.scala 123:55]
  wire [63:0] repeat_bundleIn_0_d_bits_data_mux_3 = cated_bits_data[255:192]; // @[WidthWidget.scala 123:55]
  wire [63:0] _GEN_28 = 2'h1 == repeat_index ? repeat_bundleIn_0_d_bits_data_mux_1 : repeat_bundleIn_0_d_bits_data_mux_0
    ; // @[WidthWidget.scala 132:{30,30}]
  wire [63:0] _GEN_29 = 2'h2 == repeat_index ? repeat_bundleIn_0_d_bits_data_mux_2 : _GEN_28; // @[WidthWidget.scala 132:{30,30}]
  Repeater repeated_repeater ( // @[Repeater.scala 35:26]
    .clock(repeated_repeater_clock),
    .reset(repeated_repeater_reset),
    .io_repeat(repeated_repeater_io_repeat),
    .io_enq_ready(repeated_repeater_io_enq_ready),
    .io_enq_valid(repeated_repeater_io_enq_valid),
    .io_enq_bits_opcode(repeated_repeater_io_enq_bits_opcode),
    .io_enq_bits_size(repeated_repeater_io_enq_bits_size),
    .io_enq_bits_source(repeated_repeater_io_enq_bits_source),
    .io_enq_bits_data(repeated_repeater_io_enq_bits_data),
    .io_deq_ready(repeated_repeater_io_deq_ready),
    .io_deq_valid(repeated_repeater_io_deq_valid),
    .io_deq_bits_opcode(repeated_repeater_io_deq_bits_opcode),
    .io_deq_bits_size(repeated_repeater_io_deq_bits_size),
    .io_deq_bits_source(repeated_repeater_io_deq_bits_source),
    .io_deq_bits_data(repeated_repeater_io_deq_bits_data)
  );
  assign auto_in_a_ready = auto_out_a_ready | ~last; // @[WidthWidget.scala 71:29]
  assign auto_in_d_valid = repeated_repeater_io_deq_valid; // @[WidthWidget.scala 156:25 157:15]
  assign auto_in_d_bits_data = 2'h3 == repeat_index ? repeat_bundleIn_0_d_bits_data_mux_3 : _GEN_29; // @[WidthWidget.scala 132:{30,30}]
  assign auto_out_a_valid = auto_in_a_valid & last; // @[WidthWidget.scala 72:29]
  assign auto_out_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_a_bits_mask = _x1_a_bits_mask_T_1 & _x1_a_bits_mask_T_7; // @[WidthWidget.scala 80:88]
  assign auto_out_a_bits_data = {x1_a_bits_data_hi,x1_a_bits_data_lo}; // @[Cat.scala 33:92]
  assign auto_out_d_ready = repeated_repeater_io_enq_ready; // @[Nodes.scala 1212:84 Repeater.scala 37:21]
  assign repeated_repeater_clock = clock;
  assign repeated_repeater_reset = reset;
  assign repeated_repeater_io_repeat = ~repeat_last; // @[WidthWidget.scala 143:7]
  assign repeated_repeater_io_enq_valid = auto_out_d_valid; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign repeated_repeater_io_enq_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign repeated_repeater_io_enq_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign repeated_repeater_io_enq_bits_source = auto_out_d_bits_source; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign repeated_repeater_io_enq_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign repeated_repeater_io_deq_ready = auto_in_d_ready; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  always @(posedge clock) begin
    if (reset) begin // @[WidthWidget.scala 35:27]
      count <= 2'h0; // @[WidthWidget.scala 35:27]
    end else if (_T) begin // @[WidthWidget.scala 44:24]
      if (last) begin // @[WidthWidget.scala 47:21]
        count <= 2'h0; // @[WidthWidget.scala 48:17]
      end else begin
        count <= _count_T_1; // @[WidthWidget.scala 45:15]
      end
    end
    if (reset) begin // @[WidthWidget.scala 57:41]
      x1_a_bits_data_rdata_written_once <= 1'h0; // @[WidthWidget.scala 57:41]
    end else begin
      x1_a_bits_data_rdata_written_once <= _GEN_4;
    end
    if (_T & _bundleIn_0_a_ready_T) begin // @[WidthWidget.scala 64:35]
      if (x1_a_bits_data_masked_enable_0) begin // @[WidthWidget.scala 63:88]
        x1_a_bits_data_rdata_0 <= auto_in_a_bits_data;
      end
    end
    if (_T & _bundleIn_0_a_ready_T) begin // @[WidthWidget.scala 64:35]
      if (x1_a_bits_data_masked_enable_1) begin // @[WidthWidget.scala 63:88]
        x1_a_bits_data_rdata_1 <= auto_in_a_bits_data;
      end
    end
    if (_T & _bundleIn_0_a_ready_T) begin // @[WidthWidget.scala 64:35]
      if (x1_a_bits_data_masked_enable_2) begin // @[WidthWidget.scala 63:88]
        x1_a_bits_data_rdata_2 <= auto_in_a_bits_data;
      end
    end
    if (reset) begin // @[WidthWidget.scala 57:41]
      x1_a_bits_mask_rdata_written_once <= 1'h0; // @[WidthWidget.scala 57:41]
    end else begin
      x1_a_bits_mask_rdata_written_once <= _GEN_8;
    end
    if (_T & _bundleIn_0_a_ready_T) begin // @[WidthWidget.scala 64:35]
      if (x1_a_bits_mask_masked_enable_0) begin // @[WidthWidget.scala 63:88]
        x1_a_bits_mask_rdata_0 <= auto_in_a_bits_mask;
      end
    end
    if (_T & _bundleIn_0_a_ready_T) begin // @[WidthWidget.scala 64:35]
      if (x1_a_bits_mask_masked_enable_1) begin // @[WidthWidget.scala 63:88]
        x1_a_bits_mask_rdata_1 <= auto_in_a_bits_mask;
      end
    end
    if (_T & _bundleIn_0_a_ready_T) begin // @[WidthWidget.scala 64:35]
      if (x1_a_bits_mask_masked_enable_2) begin // @[WidthWidget.scala 63:88]
        x1_a_bits_mask_rdata_2 <= auto_in_a_bits_mask;
      end
    end
    if (reset) begin // @[WidthWidget.scala 100:26]
      repeat_count <= 2'h0; // @[WidthWidget.scala 100:26]
    end else if (_repeat_T) begin // @[WidthWidget.scala 104:25]
      if (repeat_last) begin // @[WidthWidget.scala 106:21]
        repeat_count <= 2'h0; // @[WidthWidget.scala 106:29]
      end else begin
        repeat_count <= _repeat_count_T_1; // @[WidthWidget.scala 105:15]
      end
    end
    if (_T) begin // @[WidthWidget.scala 183:28]
      if (2'h0 == auto_in_a_bits_source) begin // @[WidthWidget.scala 184:37]
        repeat_sel_sel_sources_0 <= repeat_sel_sel_a_sel; // @[WidthWidget.scala 184:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 183:28]
      if (2'h1 == auto_in_a_bits_source) begin // @[WidthWidget.scala 184:37]
        repeat_sel_sel_sources_1 <= repeat_sel_sel_a_sel; // @[WidthWidget.scala 184:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 183:28]
      if (2'h2 == auto_in_a_bits_source) begin // @[WidthWidget.scala 184:37]
        repeat_sel_sel_sources_2 <= repeat_sel_sel_a_sel; // @[WidthWidget.scala 184:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 183:28]
      if (2'h3 == auto_in_a_bits_source) begin // @[WidthWidget.scala 184:37]
        repeat_sel_sel_sources_3 <= repeat_sel_sel_a_sel; // @[WidthWidget.scala 184:37]
      end
    end
    if (repeat_first) begin // @[Reg.scala 20:18]
      if (repeat_sel_sel_bypass) begin // @[WidthWidget.scala 192:17]
        repeat_sel_hold_r <= repeat_sel_sel_a_sel;
      end else if (2'h3 == cated_bits_source) begin // @[WidthWidget.scala 192:17]
        repeat_sel_hold_r <= repeat_sel_sel_sources_3; // @[WidthWidget.scala 192:17]
      end else if (2'h2 == cated_bits_source) begin // @[WidthWidget.scala 192:17]
        repeat_sel_hold_r <= repeat_sel_sel_sources_2; // @[WidthWidget.scala 192:17]
      end else begin
        repeat_sel_hold_r <= _GEN_23;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  x1_a_bits_data_rdata_written_once = _RAND_1[0:0];
  _RAND_2 = {2{`RANDOM}};
  x1_a_bits_data_rdata_0 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  x1_a_bits_data_rdata_1 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  x1_a_bits_data_rdata_2 = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  x1_a_bits_mask_rdata_written_once = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  x1_a_bits_mask_rdata_0 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  x1_a_bits_mask_rdata_1 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  x1_a_bits_mask_rdata_2 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  repeat_count = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  repeat_sel_sel_sources_0 = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  repeat_sel_sel_sources_1 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  repeat_sel_sel_sources_2 = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  repeat_sel_sel_sources_3 = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  repeat_sel_hold_r = _RAND_14[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MaxPeriodFibonacciLFSR(
  input   clock,
  input   reset,
  output  io_out_0,
  output  io_out_1,
  output  io_out_2,
  output  io_out_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg  state_0; // @[PRNG.scala 55:49]
  reg  state_1; // @[PRNG.scala 55:49]
  reg  state_2; // @[PRNG.scala 55:49]
  reg  state_3; // @[PRNG.scala 55:49]
  wire  _T = state_3 ^ state_2; // @[LFSR.scala 15:41]
  assign io_out_0 = state_0; // @[PRNG.scala 78:10]
  assign io_out_1 = state_1; // @[PRNG.scala 78:10]
  assign io_out_2 = state_2; // @[PRNG.scala 78:10]
  assign io_out_3 = state_3; // @[PRNG.scala 78:10]
  always @(posedge clock) begin
    state_0 <= reset | _T; // @[PRNG.scala 55:{49,49}]
    if (reset) begin // @[PRNG.scala 55:49]
      state_1 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_1 <= state_0;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_2 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_2 <= state_1;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_3 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_3 <= state_2;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  state_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  state_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  state_3 = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BPU(
  input         clock,
  input         reset,
  input  [63:0] io_pc,
  input  [63:0] io_jmp_packet_target,
  input         io_jmp_packet_bp_update,
  input         io_jmp_packet_bp_taken,
  input  [63:0] io_jmp_packet_bp_pc,
  output [63:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [63:0] _RAND_513;
  reg [63:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [63:0] _RAND_516;
  reg [63:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [63:0] _RAND_519;
  reg [63:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [63:0] _RAND_522;
  reg [63:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [63:0] _RAND_525;
  reg [63:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [63:0] _RAND_528;
  reg [63:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [63:0] _RAND_531;
  reg [63:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [63:0] _RAND_534;
  reg [63:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [63:0] _RAND_537;
  reg [63:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [63:0] _RAND_540;
  reg [63:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [63:0] _RAND_543;
  reg [63:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [63:0] _RAND_546;
  reg [63:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [63:0] _RAND_549;
  reg [63:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [63:0] _RAND_552;
  reg [63:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [63:0] _RAND_555;
  reg [63:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [63:0] _RAND_558;
  reg [63:0] _RAND_559;
  reg [31:0] _RAND_560;
`endif // RANDOMIZE_REG_INIT
  wire  btb_replace_idx_prng_clock; // @[PRNG.scala 91:22]
  wire  btb_replace_idx_prng_reset; // @[PRNG.scala 91:22]
  wire  btb_replace_idx_prng_io_out_0; // @[PRNG.scala 91:22]
  wire  btb_replace_idx_prng_io_out_1; // @[PRNG.scala 91:22]
  wire  btb_replace_idx_prng_io_out_2; // @[PRNG.scala 91:22]
  wire  btb_replace_idx_prng_io_out_3; // @[PRNG.scala 91:22]
  reg [8:0] ghr; // @[BPU.scala 26:20]
  reg [1:0] pht_0; // @[BPU.scala 27:20]
  reg [1:0] pht_1; // @[BPU.scala 27:20]
  reg [1:0] pht_2; // @[BPU.scala 27:20]
  reg [1:0] pht_3; // @[BPU.scala 27:20]
  reg [1:0] pht_4; // @[BPU.scala 27:20]
  reg [1:0] pht_5; // @[BPU.scala 27:20]
  reg [1:0] pht_6; // @[BPU.scala 27:20]
  reg [1:0] pht_7; // @[BPU.scala 27:20]
  reg [1:0] pht_8; // @[BPU.scala 27:20]
  reg [1:0] pht_9; // @[BPU.scala 27:20]
  reg [1:0] pht_10; // @[BPU.scala 27:20]
  reg [1:0] pht_11; // @[BPU.scala 27:20]
  reg [1:0] pht_12; // @[BPU.scala 27:20]
  reg [1:0] pht_13; // @[BPU.scala 27:20]
  reg [1:0] pht_14; // @[BPU.scala 27:20]
  reg [1:0] pht_15; // @[BPU.scala 27:20]
  reg [1:0] pht_16; // @[BPU.scala 27:20]
  reg [1:0] pht_17; // @[BPU.scala 27:20]
  reg [1:0] pht_18; // @[BPU.scala 27:20]
  reg [1:0] pht_19; // @[BPU.scala 27:20]
  reg [1:0] pht_20; // @[BPU.scala 27:20]
  reg [1:0] pht_21; // @[BPU.scala 27:20]
  reg [1:0] pht_22; // @[BPU.scala 27:20]
  reg [1:0] pht_23; // @[BPU.scala 27:20]
  reg [1:0] pht_24; // @[BPU.scala 27:20]
  reg [1:0] pht_25; // @[BPU.scala 27:20]
  reg [1:0] pht_26; // @[BPU.scala 27:20]
  reg [1:0] pht_27; // @[BPU.scala 27:20]
  reg [1:0] pht_28; // @[BPU.scala 27:20]
  reg [1:0] pht_29; // @[BPU.scala 27:20]
  reg [1:0] pht_30; // @[BPU.scala 27:20]
  reg [1:0] pht_31; // @[BPU.scala 27:20]
  reg [1:0] pht_32; // @[BPU.scala 27:20]
  reg [1:0] pht_33; // @[BPU.scala 27:20]
  reg [1:0] pht_34; // @[BPU.scala 27:20]
  reg [1:0] pht_35; // @[BPU.scala 27:20]
  reg [1:0] pht_36; // @[BPU.scala 27:20]
  reg [1:0] pht_37; // @[BPU.scala 27:20]
  reg [1:0] pht_38; // @[BPU.scala 27:20]
  reg [1:0] pht_39; // @[BPU.scala 27:20]
  reg [1:0] pht_40; // @[BPU.scala 27:20]
  reg [1:0] pht_41; // @[BPU.scala 27:20]
  reg [1:0] pht_42; // @[BPU.scala 27:20]
  reg [1:0] pht_43; // @[BPU.scala 27:20]
  reg [1:0] pht_44; // @[BPU.scala 27:20]
  reg [1:0] pht_45; // @[BPU.scala 27:20]
  reg [1:0] pht_46; // @[BPU.scala 27:20]
  reg [1:0] pht_47; // @[BPU.scala 27:20]
  reg [1:0] pht_48; // @[BPU.scala 27:20]
  reg [1:0] pht_49; // @[BPU.scala 27:20]
  reg [1:0] pht_50; // @[BPU.scala 27:20]
  reg [1:0] pht_51; // @[BPU.scala 27:20]
  reg [1:0] pht_52; // @[BPU.scala 27:20]
  reg [1:0] pht_53; // @[BPU.scala 27:20]
  reg [1:0] pht_54; // @[BPU.scala 27:20]
  reg [1:0] pht_55; // @[BPU.scala 27:20]
  reg [1:0] pht_56; // @[BPU.scala 27:20]
  reg [1:0] pht_57; // @[BPU.scala 27:20]
  reg [1:0] pht_58; // @[BPU.scala 27:20]
  reg [1:0] pht_59; // @[BPU.scala 27:20]
  reg [1:0] pht_60; // @[BPU.scala 27:20]
  reg [1:0] pht_61; // @[BPU.scala 27:20]
  reg [1:0] pht_62; // @[BPU.scala 27:20]
  reg [1:0] pht_63; // @[BPU.scala 27:20]
  reg [1:0] pht_64; // @[BPU.scala 27:20]
  reg [1:0] pht_65; // @[BPU.scala 27:20]
  reg [1:0] pht_66; // @[BPU.scala 27:20]
  reg [1:0] pht_67; // @[BPU.scala 27:20]
  reg [1:0] pht_68; // @[BPU.scala 27:20]
  reg [1:0] pht_69; // @[BPU.scala 27:20]
  reg [1:0] pht_70; // @[BPU.scala 27:20]
  reg [1:0] pht_71; // @[BPU.scala 27:20]
  reg [1:0] pht_72; // @[BPU.scala 27:20]
  reg [1:0] pht_73; // @[BPU.scala 27:20]
  reg [1:0] pht_74; // @[BPU.scala 27:20]
  reg [1:0] pht_75; // @[BPU.scala 27:20]
  reg [1:0] pht_76; // @[BPU.scala 27:20]
  reg [1:0] pht_77; // @[BPU.scala 27:20]
  reg [1:0] pht_78; // @[BPU.scala 27:20]
  reg [1:0] pht_79; // @[BPU.scala 27:20]
  reg [1:0] pht_80; // @[BPU.scala 27:20]
  reg [1:0] pht_81; // @[BPU.scala 27:20]
  reg [1:0] pht_82; // @[BPU.scala 27:20]
  reg [1:0] pht_83; // @[BPU.scala 27:20]
  reg [1:0] pht_84; // @[BPU.scala 27:20]
  reg [1:0] pht_85; // @[BPU.scala 27:20]
  reg [1:0] pht_86; // @[BPU.scala 27:20]
  reg [1:0] pht_87; // @[BPU.scala 27:20]
  reg [1:0] pht_88; // @[BPU.scala 27:20]
  reg [1:0] pht_89; // @[BPU.scala 27:20]
  reg [1:0] pht_90; // @[BPU.scala 27:20]
  reg [1:0] pht_91; // @[BPU.scala 27:20]
  reg [1:0] pht_92; // @[BPU.scala 27:20]
  reg [1:0] pht_93; // @[BPU.scala 27:20]
  reg [1:0] pht_94; // @[BPU.scala 27:20]
  reg [1:0] pht_95; // @[BPU.scala 27:20]
  reg [1:0] pht_96; // @[BPU.scala 27:20]
  reg [1:0] pht_97; // @[BPU.scala 27:20]
  reg [1:0] pht_98; // @[BPU.scala 27:20]
  reg [1:0] pht_99; // @[BPU.scala 27:20]
  reg [1:0] pht_100; // @[BPU.scala 27:20]
  reg [1:0] pht_101; // @[BPU.scala 27:20]
  reg [1:0] pht_102; // @[BPU.scala 27:20]
  reg [1:0] pht_103; // @[BPU.scala 27:20]
  reg [1:0] pht_104; // @[BPU.scala 27:20]
  reg [1:0] pht_105; // @[BPU.scala 27:20]
  reg [1:0] pht_106; // @[BPU.scala 27:20]
  reg [1:0] pht_107; // @[BPU.scala 27:20]
  reg [1:0] pht_108; // @[BPU.scala 27:20]
  reg [1:0] pht_109; // @[BPU.scala 27:20]
  reg [1:0] pht_110; // @[BPU.scala 27:20]
  reg [1:0] pht_111; // @[BPU.scala 27:20]
  reg [1:0] pht_112; // @[BPU.scala 27:20]
  reg [1:0] pht_113; // @[BPU.scala 27:20]
  reg [1:0] pht_114; // @[BPU.scala 27:20]
  reg [1:0] pht_115; // @[BPU.scala 27:20]
  reg [1:0] pht_116; // @[BPU.scala 27:20]
  reg [1:0] pht_117; // @[BPU.scala 27:20]
  reg [1:0] pht_118; // @[BPU.scala 27:20]
  reg [1:0] pht_119; // @[BPU.scala 27:20]
  reg [1:0] pht_120; // @[BPU.scala 27:20]
  reg [1:0] pht_121; // @[BPU.scala 27:20]
  reg [1:0] pht_122; // @[BPU.scala 27:20]
  reg [1:0] pht_123; // @[BPU.scala 27:20]
  reg [1:0] pht_124; // @[BPU.scala 27:20]
  reg [1:0] pht_125; // @[BPU.scala 27:20]
  reg [1:0] pht_126; // @[BPU.scala 27:20]
  reg [1:0] pht_127; // @[BPU.scala 27:20]
  reg [1:0] pht_128; // @[BPU.scala 27:20]
  reg [1:0] pht_129; // @[BPU.scala 27:20]
  reg [1:0] pht_130; // @[BPU.scala 27:20]
  reg [1:0] pht_131; // @[BPU.scala 27:20]
  reg [1:0] pht_132; // @[BPU.scala 27:20]
  reg [1:0] pht_133; // @[BPU.scala 27:20]
  reg [1:0] pht_134; // @[BPU.scala 27:20]
  reg [1:0] pht_135; // @[BPU.scala 27:20]
  reg [1:0] pht_136; // @[BPU.scala 27:20]
  reg [1:0] pht_137; // @[BPU.scala 27:20]
  reg [1:0] pht_138; // @[BPU.scala 27:20]
  reg [1:0] pht_139; // @[BPU.scala 27:20]
  reg [1:0] pht_140; // @[BPU.scala 27:20]
  reg [1:0] pht_141; // @[BPU.scala 27:20]
  reg [1:0] pht_142; // @[BPU.scala 27:20]
  reg [1:0] pht_143; // @[BPU.scala 27:20]
  reg [1:0] pht_144; // @[BPU.scala 27:20]
  reg [1:0] pht_145; // @[BPU.scala 27:20]
  reg [1:0] pht_146; // @[BPU.scala 27:20]
  reg [1:0] pht_147; // @[BPU.scala 27:20]
  reg [1:0] pht_148; // @[BPU.scala 27:20]
  reg [1:0] pht_149; // @[BPU.scala 27:20]
  reg [1:0] pht_150; // @[BPU.scala 27:20]
  reg [1:0] pht_151; // @[BPU.scala 27:20]
  reg [1:0] pht_152; // @[BPU.scala 27:20]
  reg [1:0] pht_153; // @[BPU.scala 27:20]
  reg [1:0] pht_154; // @[BPU.scala 27:20]
  reg [1:0] pht_155; // @[BPU.scala 27:20]
  reg [1:0] pht_156; // @[BPU.scala 27:20]
  reg [1:0] pht_157; // @[BPU.scala 27:20]
  reg [1:0] pht_158; // @[BPU.scala 27:20]
  reg [1:0] pht_159; // @[BPU.scala 27:20]
  reg [1:0] pht_160; // @[BPU.scala 27:20]
  reg [1:0] pht_161; // @[BPU.scala 27:20]
  reg [1:0] pht_162; // @[BPU.scala 27:20]
  reg [1:0] pht_163; // @[BPU.scala 27:20]
  reg [1:0] pht_164; // @[BPU.scala 27:20]
  reg [1:0] pht_165; // @[BPU.scala 27:20]
  reg [1:0] pht_166; // @[BPU.scala 27:20]
  reg [1:0] pht_167; // @[BPU.scala 27:20]
  reg [1:0] pht_168; // @[BPU.scala 27:20]
  reg [1:0] pht_169; // @[BPU.scala 27:20]
  reg [1:0] pht_170; // @[BPU.scala 27:20]
  reg [1:0] pht_171; // @[BPU.scala 27:20]
  reg [1:0] pht_172; // @[BPU.scala 27:20]
  reg [1:0] pht_173; // @[BPU.scala 27:20]
  reg [1:0] pht_174; // @[BPU.scala 27:20]
  reg [1:0] pht_175; // @[BPU.scala 27:20]
  reg [1:0] pht_176; // @[BPU.scala 27:20]
  reg [1:0] pht_177; // @[BPU.scala 27:20]
  reg [1:0] pht_178; // @[BPU.scala 27:20]
  reg [1:0] pht_179; // @[BPU.scala 27:20]
  reg [1:0] pht_180; // @[BPU.scala 27:20]
  reg [1:0] pht_181; // @[BPU.scala 27:20]
  reg [1:0] pht_182; // @[BPU.scala 27:20]
  reg [1:0] pht_183; // @[BPU.scala 27:20]
  reg [1:0] pht_184; // @[BPU.scala 27:20]
  reg [1:0] pht_185; // @[BPU.scala 27:20]
  reg [1:0] pht_186; // @[BPU.scala 27:20]
  reg [1:0] pht_187; // @[BPU.scala 27:20]
  reg [1:0] pht_188; // @[BPU.scala 27:20]
  reg [1:0] pht_189; // @[BPU.scala 27:20]
  reg [1:0] pht_190; // @[BPU.scala 27:20]
  reg [1:0] pht_191; // @[BPU.scala 27:20]
  reg [1:0] pht_192; // @[BPU.scala 27:20]
  reg [1:0] pht_193; // @[BPU.scala 27:20]
  reg [1:0] pht_194; // @[BPU.scala 27:20]
  reg [1:0] pht_195; // @[BPU.scala 27:20]
  reg [1:0] pht_196; // @[BPU.scala 27:20]
  reg [1:0] pht_197; // @[BPU.scala 27:20]
  reg [1:0] pht_198; // @[BPU.scala 27:20]
  reg [1:0] pht_199; // @[BPU.scala 27:20]
  reg [1:0] pht_200; // @[BPU.scala 27:20]
  reg [1:0] pht_201; // @[BPU.scala 27:20]
  reg [1:0] pht_202; // @[BPU.scala 27:20]
  reg [1:0] pht_203; // @[BPU.scala 27:20]
  reg [1:0] pht_204; // @[BPU.scala 27:20]
  reg [1:0] pht_205; // @[BPU.scala 27:20]
  reg [1:0] pht_206; // @[BPU.scala 27:20]
  reg [1:0] pht_207; // @[BPU.scala 27:20]
  reg [1:0] pht_208; // @[BPU.scala 27:20]
  reg [1:0] pht_209; // @[BPU.scala 27:20]
  reg [1:0] pht_210; // @[BPU.scala 27:20]
  reg [1:0] pht_211; // @[BPU.scala 27:20]
  reg [1:0] pht_212; // @[BPU.scala 27:20]
  reg [1:0] pht_213; // @[BPU.scala 27:20]
  reg [1:0] pht_214; // @[BPU.scala 27:20]
  reg [1:0] pht_215; // @[BPU.scala 27:20]
  reg [1:0] pht_216; // @[BPU.scala 27:20]
  reg [1:0] pht_217; // @[BPU.scala 27:20]
  reg [1:0] pht_218; // @[BPU.scala 27:20]
  reg [1:0] pht_219; // @[BPU.scala 27:20]
  reg [1:0] pht_220; // @[BPU.scala 27:20]
  reg [1:0] pht_221; // @[BPU.scala 27:20]
  reg [1:0] pht_222; // @[BPU.scala 27:20]
  reg [1:0] pht_223; // @[BPU.scala 27:20]
  reg [1:0] pht_224; // @[BPU.scala 27:20]
  reg [1:0] pht_225; // @[BPU.scala 27:20]
  reg [1:0] pht_226; // @[BPU.scala 27:20]
  reg [1:0] pht_227; // @[BPU.scala 27:20]
  reg [1:0] pht_228; // @[BPU.scala 27:20]
  reg [1:0] pht_229; // @[BPU.scala 27:20]
  reg [1:0] pht_230; // @[BPU.scala 27:20]
  reg [1:0] pht_231; // @[BPU.scala 27:20]
  reg [1:0] pht_232; // @[BPU.scala 27:20]
  reg [1:0] pht_233; // @[BPU.scala 27:20]
  reg [1:0] pht_234; // @[BPU.scala 27:20]
  reg [1:0] pht_235; // @[BPU.scala 27:20]
  reg [1:0] pht_236; // @[BPU.scala 27:20]
  reg [1:0] pht_237; // @[BPU.scala 27:20]
  reg [1:0] pht_238; // @[BPU.scala 27:20]
  reg [1:0] pht_239; // @[BPU.scala 27:20]
  reg [1:0] pht_240; // @[BPU.scala 27:20]
  reg [1:0] pht_241; // @[BPU.scala 27:20]
  reg [1:0] pht_242; // @[BPU.scala 27:20]
  reg [1:0] pht_243; // @[BPU.scala 27:20]
  reg [1:0] pht_244; // @[BPU.scala 27:20]
  reg [1:0] pht_245; // @[BPU.scala 27:20]
  reg [1:0] pht_246; // @[BPU.scala 27:20]
  reg [1:0] pht_247; // @[BPU.scala 27:20]
  reg [1:0] pht_248; // @[BPU.scala 27:20]
  reg [1:0] pht_249; // @[BPU.scala 27:20]
  reg [1:0] pht_250; // @[BPU.scala 27:20]
  reg [1:0] pht_251; // @[BPU.scala 27:20]
  reg [1:0] pht_252; // @[BPU.scala 27:20]
  reg [1:0] pht_253; // @[BPU.scala 27:20]
  reg [1:0] pht_254; // @[BPU.scala 27:20]
  reg [1:0] pht_255; // @[BPU.scala 27:20]
  reg [1:0] pht_256; // @[BPU.scala 27:20]
  reg [1:0] pht_257; // @[BPU.scala 27:20]
  reg [1:0] pht_258; // @[BPU.scala 27:20]
  reg [1:0] pht_259; // @[BPU.scala 27:20]
  reg [1:0] pht_260; // @[BPU.scala 27:20]
  reg [1:0] pht_261; // @[BPU.scala 27:20]
  reg [1:0] pht_262; // @[BPU.scala 27:20]
  reg [1:0] pht_263; // @[BPU.scala 27:20]
  reg [1:0] pht_264; // @[BPU.scala 27:20]
  reg [1:0] pht_265; // @[BPU.scala 27:20]
  reg [1:0] pht_266; // @[BPU.scala 27:20]
  reg [1:0] pht_267; // @[BPU.scala 27:20]
  reg [1:0] pht_268; // @[BPU.scala 27:20]
  reg [1:0] pht_269; // @[BPU.scala 27:20]
  reg [1:0] pht_270; // @[BPU.scala 27:20]
  reg [1:0] pht_271; // @[BPU.scala 27:20]
  reg [1:0] pht_272; // @[BPU.scala 27:20]
  reg [1:0] pht_273; // @[BPU.scala 27:20]
  reg [1:0] pht_274; // @[BPU.scala 27:20]
  reg [1:0] pht_275; // @[BPU.scala 27:20]
  reg [1:0] pht_276; // @[BPU.scala 27:20]
  reg [1:0] pht_277; // @[BPU.scala 27:20]
  reg [1:0] pht_278; // @[BPU.scala 27:20]
  reg [1:0] pht_279; // @[BPU.scala 27:20]
  reg [1:0] pht_280; // @[BPU.scala 27:20]
  reg [1:0] pht_281; // @[BPU.scala 27:20]
  reg [1:0] pht_282; // @[BPU.scala 27:20]
  reg [1:0] pht_283; // @[BPU.scala 27:20]
  reg [1:0] pht_284; // @[BPU.scala 27:20]
  reg [1:0] pht_285; // @[BPU.scala 27:20]
  reg [1:0] pht_286; // @[BPU.scala 27:20]
  reg [1:0] pht_287; // @[BPU.scala 27:20]
  reg [1:0] pht_288; // @[BPU.scala 27:20]
  reg [1:0] pht_289; // @[BPU.scala 27:20]
  reg [1:0] pht_290; // @[BPU.scala 27:20]
  reg [1:0] pht_291; // @[BPU.scala 27:20]
  reg [1:0] pht_292; // @[BPU.scala 27:20]
  reg [1:0] pht_293; // @[BPU.scala 27:20]
  reg [1:0] pht_294; // @[BPU.scala 27:20]
  reg [1:0] pht_295; // @[BPU.scala 27:20]
  reg [1:0] pht_296; // @[BPU.scala 27:20]
  reg [1:0] pht_297; // @[BPU.scala 27:20]
  reg [1:0] pht_298; // @[BPU.scala 27:20]
  reg [1:0] pht_299; // @[BPU.scala 27:20]
  reg [1:0] pht_300; // @[BPU.scala 27:20]
  reg [1:0] pht_301; // @[BPU.scala 27:20]
  reg [1:0] pht_302; // @[BPU.scala 27:20]
  reg [1:0] pht_303; // @[BPU.scala 27:20]
  reg [1:0] pht_304; // @[BPU.scala 27:20]
  reg [1:0] pht_305; // @[BPU.scala 27:20]
  reg [1:0] pht_306; // @[BPU.scala 27:20]
  reg [1:0] pht_307; // @[BPU.scala 27:20]
  reg [1:0] pht_308; // @[BPU.scala 27:20]
  reg [1:0] pht_309; // @[BPU.scala 27:20]
  reg [1:0] pht_310; // @[BPU.scala 27:20]
  reg [1:0] pht_311; // @[BPU.scala 27:20]
  reg [1:0] pht_312; // @[BPU.scala 27:20]
  reg [1:0] pht_313; // @[BPU.scala 27:20]
  reg [1:0] pht_314; // @[BPU.scala 27:20]
  reg [1:0] pht_315; // @[BPU.scala 27:20]
  reg [1:0] pht_316; // @[BPU.scala 27:20]
  reg [1:0] pht_317; // @[BPU.scala 27:20]
  reg [1:0] pht_318; // @[BPU.scala 27:20]
  reg [1:0] pht_319; // @[BPU.scala 27:20]
  reg [1:0] pht_320; // @[BPU.scala 27:20]
  reg [1:0] pht_321; // @[BPU.scala 27:20]
  reg [1:0] pht_322; // @[BPU.scala 27:20]
  reg [1:0] pht_323; // @[BPU.scala 27:20]
  reg [1:0] pht_324; // @[BPU.scala 27:20]
  reg [1:0] pht_325; // @[BPU.scala 27:20]
  reg [1:0] pht_326; // @[BPU.scala 27:20]
  reg [1:0] pht_327; // @[BPU.scala 27:20]
  reg [1:0] pht_328; // @[BPU.scala 27:20]
  reg [1:0] pht_329; // @[BPU.scala 27:20]
  reg [1:0] pht_330; // @[BPU.scala 27:20]
  reg [1:0] pht_331; // @[BPU.scala 27:20]
  reg [1:0] pht_332; // @[BPU.scala 27:20]
  reg [1:0] pht_333; // @[BPU.scala 27:20]
  reg [1:0] pht_334; // @[BPU.scala 27:20]
  reg [1:0] pht_335; // @[BPU.scala 27:20]
  reg [1:0] pht_336; // @[BPU.scala 27:20]
  reg [1:0] pht_337; // @[BPU.scala 27:20]
  reg [1:0] pht_338; // @[BPU.scala 27:20]
  reg [1:0] pht_339; // @[BPU.scala 27:20]
  reg [1:0] pht_340; // @[BPU.scala 27:20]
  reg [1:0] pht_341; // @[BPU.scala 27:20]
  reg [1:0] pht_342; // @[BPU.scala 27:20]
  reg [1:0] pht_343; // @[BPU.scala 27:20]
  reg [1:0] pht_344; // @[BPU.scala 27:20]
  reg [1:0] pht_345; // @[BPU.scala 27:20]
  reg [1:0] pht_346; // @[BPU.scala 27:20]
  reg [1:0] pht_347; // @[BPU.scala 27:20]
  reg [1:0] pht_348; // @[BPU.scala 27:20]
  reg [1:0] pht_349; // @[BPU.scala 27:20]
  reg [1:0] pht_350; // @[BPU.scala 27:20]
  reg [1:0] pht_351; // @[BPU.scala 27:20]
  reg [1:0] pht_352; // @[BPU.scala 27:20]
  reg [1:0] pht_353; // @[BPU.scala 27:20]
  reg [1:0] pht_354; // @[BPU.scala 27:20]
  reg [1:0] pht_355; // @[BPU.scala 27:20]
  reg [1:0] pht_356; // @[BPU.scala 27:20]
  reg [1:0] pht_357; // @[BPU.scala 27:20]
  reg [1:0] pht_358; // @[BPU.scala 27:20]
  reg [1:0] pht_359; // @[BPU.scala 27:20]
  reg [1:0] pht_360; // @[BPU.scala 27:20]
  reg [1:0] pht_361; // @[BPU.scala 27:20]
  reg [1:0] pht_362; // @[BPU.scala 27:20]
  reg [1:0] pht_363; // @[BPU.scala 27:20]
  reg [1:0] pht_364; // @[BPU.scala 27:20]
  reg [1:0] pht_365; // @[BPU.scala 27:20]
  reg [1:0] pht_366; // @[BPU.scala 27:20]
  reg [1:0] pht_367; // @[BPU.scala 27:20]
  reg [1:0] pht_368; // @[BPU.scala 27:20]
  reg [1:0] pht_369; // @[BPU.scala 27:20]
  reg [1:0] pht_370; // @[BPU.scala 27:20]
  reg [1:0] pht_371; // @[BPU.scala 27:20]
  reg [1:0] pht_372; // @[BPU.scala 27:20]
  reg [1:0] pht_373; // @[BPU.scala 27:20]
  reg [1:0] pht_374; // @[BPU.scala 27:20]
  reg [1:0] pht_375; // @[BPU.scala 27:20]
  reg [1:0] pht_376; // @[BPU.scala 27:20]
  reg [1:0] pht_377; // @[BPU.scala 27:20]
  reg [1:0] pht_378; // @[BPU.scala 27:20]
  reg [1:0] pht_379; // @[BPU.scala 27:20]
  reg [1:0] pht_380; // @[BPU.scala 27:20]
  reg [1:0] pht_381; // @[BPU.scala 27:20]
  reg [1:0] pht_382; // @[BPU.scala 27:20]
  reg [1:0] pht_383; // @[BPU.scala 27:20]
  reg [1:0] pht_384; // @[BPU.scala 27:20]
  reg [1:0] pht_385; // @[BPU.scala 27:20]
  reg [1:0] pht_386; // @[BPU.scala 27:20]
  reg [1:0] pht_387; // @[BPU.scala 27:20]
  reg [1:0] pht_388; // @[BPU.scala 27:20]
  reg [1:0] pht_389; // @[BPU.scala 27:20]
  reg [1:0] pht_390; // @[BPU.scala 27:20]
  reg [1:0] pht_391; // @[BPU.scala 27:20]
  reg [1:0] pht_392; // @[BPU.scala 27:20]
  reg [1:0] pht_393; // @[BPU.scala 27:20]
  reg [1:0] pht_394; // @[BPU.scala 27:20]
  reg [1:0] pht_395; // @[BPU.scala 27:20]
  reg [1:0] pht_396; // @[BPU.scala 27:20]
  reg [1:0] pht_397; // @[BPU.scala 27:20]
  reg [1:0] pht_398; // @[BPU.scala 27:20]
  reg [1:0] pht_399; // @[BPU.scala 27:20]
  reg [1:0] pht_400; // @[BPU.scala 27:20]
  reg [1:0] pht_401; // @[BPU.scala 27:20]
  reg [1:0] pht_402; // @[BPU.scala 27:20]
  reg [1:0] pht_403; // @[BPU.scala 27:20]
  reg [1:0] pht_404; // @[BPU.scala 27:20]
  reg [1:0] pht_405; // @[BPU.scala 27:20]
  reg [1:0] pht_406; // @[BPU.scala 27:20]
  reg [1:0] pht_407; // @[BPU.scala 27:20]
  reg [1:0] pht_408; // @[BPU.scala 27:20]
  reg [1:0] pht_409; // @[BPU.scala 27:20]
  reg [1:0] pht_410; // @[BPU.scala 27:20]
  reg [1:0] pht_411; // @[BPU.scala 27:20]
  reg [1:0] pht_412; // @[BPU.scala 27:20]
  reg [1:0] pht_413; // @[BPU.scala 27:20]
  reg [1:0] pht_414; // @[BPU.scala 27:20]
  reg [1:0] pht_415; // @[BPU.scala 27:20]
  reg [1:0] pht_416; // @[BPU.scala 27:20]
  reg [1:0] pht_417; // @[BPU.scala 27:20]
  reg [1:0] pht_418; // @[BPU.scala 27:20]
  reg [1:0] pht_419; // @[BPU.scala 27:20]
  reg [1:0] pht_420; // @[BPU.scala 27:20]
  reg [1:0] pht_421; // @[BPU.scala 27:20]
  reg [1:0] pht_422; // @[BPU.scala 27:20]
  reg [1:0] pht_423; // @[BPU.scala 27:20]
  reg [1:0] pht_424; // @[BPU.scala 27:20]
  reg [1:0] pht_425; // @[BPU.scala 27:20]
  reg [1:0] pht_426; // @[BPU.scala 27:20]
  reg [1:0] pht_427; // @[BPU.scala 27:20]
  reg [1:0] pht_428; // @[BPU.scala 27:20]
  reg [1:0] pht_429; // @[BPU.scala 27:20]
  reg [1:0] pht_430; // @[BPU.scala 27:20]
  reg [1:0] pht_431; // @[BPU.scala 27:20]
  reg [1:0] pht_432; // @[BPU.scala 27:20]
  reg [1:0] pht_433; // @[BPU.scala 27:20]
  reg [1:0] pht_434; // @[BPU.scala 27:20]
  reg [1:0] pht_435; // @[BPU.scala 27:20]
  reg [1:0] pht_436; // @[BPU.scala 27:20]
  reg [1:0] pht_437; // @[BPU.scala 27:20]
  reg [1:0] pht_438; // @[BPU.scala 27:20]
  reg [1:0] pht_439; // @[BPU.scala 27:20]
  reg [1:0] pht_440; // @[BPU.scala 27:20]
  reg [1:0] pht_441; // @[BPU.scala 27:20]
  reg [1:0] pht_442; // @[BPU.scala 27:20]
  reg [1:0] pht_443; // @[BPU.scala 27:20]
  reg [1:0] pht_444; // @[BPU.scala 27:20]
  reg [1:0] pht_445; // @[BPU.scala 27:20]
  reg [1:0] pht_446; // @[BPU.scala 27:20]
  reg [1:0] pht_447; // @[BPU.scala 27:20]
  reg [1:0] pht_448; // @[BPU.scala 27:20]
  reg [1:0] pht_449; // @[BPU.scala 27:20]
  reg [1:0] pht_450; // @[BPU.scala 27:20]
  reg [1:0] pht_451; // @[BPU.scala 27:20]
  reg [1:0] pht_452; // @[BPU.scala 27:20]
  reg [1:0] pht_453; // @[BPU.scala 27:20]
  reg [1:0] pht_454; // @[BPU.scala 27:20]
  reg [1:0] pht_455; // @[BPU.scala 27:20]
  reg [1:0] pht_456; // @[BPU.scala 27:20]
  reg [1:0] pht_457; // @[BPU.scala 27:20]
  reg [1:0] pht_458; // @[BPU.scala 27:20]
  reg [1:0] pht_459; // @[BPU.scala 27:20]
  reg [1:0] pht_460; // @[BPU.scala 27:20]
  reg [1:0] pht_461; // @[BPU.scala 27:20]
  reg [1:0] pht_462; // @[BPU.scala 27:20]
  reg [1:0] pht_463; // @[BPU.scala 27:20]
  reg [1:0] pht_464; // @[BPU.scala 27:20]
  reg [1:0] pht_465; // @[BPU.scala 27:20]
  reg [1:0] pht_466; // @[BPU.scala 27:20]
  reg [1:0] pht_467; // @[BPU.scala 27:20]
  reg [1:0] pht_468; // @[BPU.scala 27:20]
  reg [1:0] pht_469; // @[BPU.scala 27:20]
  reg [1:0] pht_470; // @[BPU.scala 27:20]
  reg [1:0] pht_471; // @[BPU.scala 27:20]
  reg [1:0] pht_472; // @[BPU.scala 27:20]
  reg [1:0] pht_473; // @[BPU.scala 27:20]
  reg [1:0] pht_474; // @[BPU.scala 27:20]
  reg [1:0] pht_475; // @[BPU.scala 27:20]
  reg [1:0] pht_476; // @[BPU.scala 27:20]
  reg [1:0] pht_477; // @[BPU.scala 27:20]
  reg [1:0] pht_478; // @[BPU.scala 27:20]
  reg [1:0] pht_479; // @[BPU.scala 27:20]
  reg [1:0] pht_480; // @[BPU.scala 27:20]
  reg [1:0] pht_481; // @[BPU.scala 27:20]
  reg [1:0] pht_482; // @[BPU.scala 27:20]
  reg [1:0] pht_483; // @[BPU.scala 27:20]
  reg [1:0] pht_484; // @[BPU.scala 27:20]
  reg [1:0] pht_485; // @[BPU.scala 27:20]
  reg [1:0] pht_486; // @[BPU.scala 27:20]
  reg [1:0] pht_487; // @[BPU.scala 27:20]
  reg [1:0] pht_488; // @[BPU.scala 27:20]
  reg [1:0] pht_489; // @[BPU.scala 27:20]
  reg [1:0] pht_490; // @[BPU.scala 27:20]
  reg [1:0] pht_491; // @[BPU.scala 27:20]
  reg [1:0] pht_492; // @[BPU.scala 27:20]
  reg [1:0] pht_493; // @[BPU.scala 27:20]
  reg [1:0] pht_494; // @[BPU.scala 27:20]
  reg [1:0] pht_495; // @[BPU.scala 27:20]
  reg [1:0] pht_496; // @[BPU.scala 27:20]
  reg [1:0] pht_497; // @[BPU.scala 27:20]
  reg [1:0] pht_498; // @[BPU.scala 27:20]
  reg [1:0] pht_499; // @[BPU.scala 27:20]
  reg [1:0] pht_500; // @[BPU.scala 27:20]
  reg [1:0] pht_501; // @[BPU.scala 27:20]
  reg [1:0] pht_502; // @[BPU.scala 27:20]
  reg [1:0] pht_503; // @[BPU.scala 27:20]
  reg [1:0] pht_504; // @[BPU.scala 27:20]
  reg [1:0] pht_505; // @[BPU.scala 27:20]
  reg [1:0] pht_506; // @[BPU.scala 27:20]
  reg [1:0] pht_507; // @[BPU.scala 27:20]
  reg [1:0] pht_508; // @[BPU.scala 27:20]
  reg [1:0] pht_509; // @[BPU.scala 27:20]
  reg [1:0] pht_510; // @[BPU.scala 27:20]
  reg [1:0] pht_511; // @[BPU.scala 27:20]
  reg [36:0] btb_0_tag; // @[BPU.scala 28:20]
  reg [36:0] btb_0_target; // @[BPU.scala 28:20]
  reg  btb_0_valid; // @[BPU.scala 28:20]
  reg [36:0] btb_1_tag; // @[BPU.scala 28:20]
  reg [36:0] btb_1_target; // @[BPU.scala 28:20]
  reg  btb_1_valid; // @[BPU.scala 28:20]
  reg [36:0] btb_2_tag; // @[BPU.scala 28:20]
  reg [36:0] btb_2_target; // @[BPU.scala 28:20]
  reg  btb_2_valid; // @[BPU.scala 28:20]
  reg [36:0] btb_3_tag; // @[BPU.scala 28:20]
  reg [36:0] btb_3_target; // @[BPU.scala 28:20]
  reg  btb_3_valid; // @[BPU.scala 28:20]
  reg [36:0] btb_4_tag; // @[BPU.scala 28:20]
  reg [36:0] btb_4_target; // @[BPU.scala 28:20]
  reg  btb_4_valid; // @[BPU.scala 28:20]
  reg [36:0] btb_5_tag; // @[BPU.scala 28:20]
  reg [36:0] btb_5_target; // @[BPU.scala 28:20]
  reg  btb_5_valid; // @[BPU.scala 28:20]
  reg [36:0] btb_6_tag; // @[BPU.scala 28:20]
  reg [36:0] btb_6_target; // @[BPU.scala 28:20]
  reg  btb_6_valid; // @[BPU.scala 28:20]
  reg [36:0] btb_7_tag; // @[BPU.scala 28:20]
  reg [36:0] btb_7_target; // @[BPU.scala 28:20]
  reg  btb_7_valid; // @[BPU.scala 28:20]
  reg [36:0] btb_8_tag; // @[BPU.scala 28:20]
  reg [36:0] btb_8_target; // @[BPU.scala 28:20]
  reg  btb_8_valid; // @[BPU.scala 28:20]
  reg [36:0] btb_9_tag; // @[BPU.scala 28:20]
  reg [36:0] btb_9_target; // @[BPU.scala 28:20]
  reg  btb_9_valid; // @[BPU.scala 28:20]
  reg [36:0] btb_10_tag; // @[BPU.scala 28:20]
  reg [36:0] btb_10_target; // @[BPU.scala 28:20]
  reg  btb_10_valid; // @[BPU.scala 28:20]
  reg [36:0] btb_11_tag; // @[BPU.scala 28:20]
  reg [36:0] btb_11_target; // @[BPU.scala 28:20]
  reg  btb_11_valid; // @[BPU.scala 28:20]
  reg [36:0] btb_12_tag; // @[BPU.scala 28:20]
  reg [36:0] btb_12_target; // @[BPU.scala 28:20]
  reg  btb_12_valid; // @[BPU.scala 28:20]
  reg [36:0] btb_13_tag; // @[BPU.scala 28:20]
  reg [36:0] btb_13_target; // @[BPU.scala 28:20]
  reg  btb_13_valid; // @[BPU.scala 28:20]
  reg [36:0] btb_14_tag; // @[BPU.scala 28:20]
  reg [36:0] btb_14_target; // @[BPU.scala 28:20]
  reg  btb_14_valid; // @[BPU.scala 28:20]
  reg [36:0] btb_15_tag; // @[BPU.scala 28:20]
  reg [36:0] btb_15_target; // @[BPU.scala 28:20]
  reg  btb_15_valid; // @[BPU.scala 28:20]
  wire [8:0] pht_ridx = io_pc[10:2] ^ ghr; // @[BPU.scala 31:40]
  wire [1:0] _GEN_1 = 9'h1 == pht_ridx ? pht_1 : pht_0; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_2 = 9'h2 == pht_ridx ? pht_2 : _GEN_1; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_3 = 9'h3 == pht_ridx ? pht_3 : _GEN_2; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_4 = 9'h4 == pht_ridx ? pht_4 : _GEN_3; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_5 = 9'h5 == pht_ridx ? pht_5 : _GEN_4; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_6 = 9'h6 == pht_ridx ? pht_6 : _GEN_5; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_7 = 9'h7 == pht_ridx ? pht_7 : _GEN_6; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_8 = 9'h8 == pht_ridx ? pht_8 : _GEN_7; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_9 = 9'h9 == pht_ridx ? pht_9 : _GEN_8; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_10 = 9'ha == pht_ridx ? pht_10 : _GEN_9; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_11 = 9'hb == pht_ridx ? pht_11 : _GEN_10; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_12 = 9'hc == pht_ridx ? pht_12 : _GEN_11; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_13 = 9'hd == pht_ridx ? pht_13 : _GEN_12; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_14 = 9'he == pht_ridx ? pht_14 : _GEN_13; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_15 = 9'hf == pht_ridx ? pht_15 : _GEN_14; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_16 = 9'h10 == pht_ridx ? pht_16 : _GEN_15; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_17 = 9'h11 == pht_ridx ? pht_17 : _GEN_16; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_18 = 9'h12 == pht_ridx ? pht_18 : _GEN_17; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_19 = 9'h13 == pht_ridx ? pht_19 : _GEN_18; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_20 = 9'h14 == pht_ridx ? pht_20 : _GEN_19; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_21 = 9'h15 == pht_ridx ? pht_21 : _GEN_20; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_22 = 9'h16 == pht_ridx ? pht_22 : _GEN_21; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_23 = 9'h17 == pht_ridx ? pht_23 : _GEN_22; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_24 = 9'h18 == pht_ridx ? pht_24 : _GEN_23; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_25 = 9'h19 == pht_ridx ? pht_25 : _GEN_24; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_26 = 9'h1a == pht_ridx ? pht_26 : _GEN_25; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_27 = 9'h1b == pht_ridx ? pht_27 : _GEN_26; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_28 = 9'h1c == pht_ridx ? pht_28 : _GEN_27; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_29 = 9'h1d == pht_ridx ? pht_29 : _GEN_28; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_30 = 9'h1e == pht_ridx ? pht_30 : _GEN_29; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_31 = 9'h1f == pht_ridx ? pht_31 : _GEN_30; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_32 = 9'h20 == pht_ridx ? pht_32 : _GEN_31; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_33 = 9'h21 == pht_ridx ? pht_33 : _GEN_32; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_34 = 9'h22 == pht_ridx ? pht_34 : _GEN_33; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_35 = 9'h23 == pht_ridx ? pht_35 : _GEN_34; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_36 = 9'h24 == pht_ridx ? pht_36 : _GEN_35; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_37 = 9'h25 == pht_ridx ? pht_37 : _GEN_36; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_38 = 9'h26 == pht_ridx ? pht_38 : _GEN_37; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_39 = 9'h27 == pht_ridx ? pht_39 : _GEN_38; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_40 = 9'h28 == pht_ridx ? pht_40 : _GEN_39; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_41 = 9'h29 == pht_ridx ? pht_41 : _GEN_40; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_42 = 9'h2a == pht_ridx ? pht_42 : _GEN_41; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_43 = 9'h2b == pht_ridx ? pht_43 : _GEN_42; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_44 = 9'h2c == pht_ridx ? pht_44 : _GEN_43; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_45 = 9'h2d == pht_ridx ? pht_45 : _GEN_44; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_46 = 9'h2e == pht_ridx ? pht_46 : _GEN_45; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_47 = 9'h2f == pht_ridx ? pht_47 : _GEN_46; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_48 = 9'h30 == pht_ridx ? pht_48 : _GEN_47; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_49 = 9'h31 == pht_ridx ? pht_49 : _GEN_48; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_50 = 9'h32 == pht_ridx ? pht_50 : _GEN_49; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_51 = 9'h33 == pht_ridx ? pht_51 : _GEN_50; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_52 = 9'h34 == pht_ridx ? pht_52 : _GEN_51; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_53 = 9'h35 == pht_ridx ? pht_53 : _GEN_52; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_54 = 9'h36 == pht_ridx ? pht_54 : _GEN_53; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_55 = 9'h37 == pht_ridx ? pht_55 : _GEN_54; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_56 = 9'h38 == pht_ridx ? pht_56 : _GEN_55; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_57 = 9'h39 == pht_ridx ? pht_57 : _GEN_56; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_58 = 9'h3a == pht_ridx ? pht_58 : _GEN_57; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_59 = 9'h3b == pht_ridx ? pht_59 : _GEN_58; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_60 = 9'h3c == pht_ridx ? pht_60 : _GEN_59; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_61 = 9'h3d == pht_ridx ? pht_61 : _GEN_60; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_62 = 9'h3e == pht_ridx ? pht_62 : _GEN_61; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_63 = 9'h3f == pht_ridx ? pht_63 : _GEN_62; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_64 = 9'h40 == pht_ridx ? pht_64 : _GEN_63; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_65 = 9'h41 == pht_ridx ? pht_65 : _GEN_64; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_66 = 9'h42 == pht_ridx ? pht_66 : _GEN_65; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_67 = 9'h43 == pht_ridx ? pht_67 : _GEN_66; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_68 = 9'h44 == pht_ridx ? pht_68 : _GEN_67; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_69 = 9'h45 == pht_ridx ? pht_69 : _GEN_68; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_70 = 9'h46 == pht_ridx ? pht_70 : _GEN_69; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_71 = 9'h47 == pht_ridx ? pht_71 : _GEN_70; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_72 = 9'h48 == pht_ridx ? pht_72 : _GEN_71; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_73 = 9'h49 == pht_ridx ? pht_73 : _GEN_72; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_74 = 9'h4a == pht_ridx ? pht_74 : _GEN_73; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_75 = 9'h4b == pht_ridx ? pht_75 : _GEN_74; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_76 = 9'h4c == pht_ridx ? pht_76 : _GEN_75; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_77 = 9'h4d == pht_ridx ? pht_77 : _GEN_76; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_78 = 9'h4e == pht_ridx ? pht_78 : _GEN_77; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_79 = 9'h4f == pht_ridx ? pht_79 : _GEN_78; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_80 = 9'h50 == pht_ridx ? pht_80 : _GEN_79; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_81 = 9'h51 == pht_ridx ? pht_81 : _GEN_80; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_82 = 9'h52 == pht_ridx ? pht_82 : _GEN_81; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_83 = 9'h53 == pht_ridx ? pht_83 : _GEN_82; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_84 = 9'h54 == pht_ridx ? pht_84 : _GEN_83; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_85 = 9'h55 == pht_ridx ? pht_85 : _GEN_84; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_86 = 9'h56 == pht_ridx ? pht_86 : _GEN_85; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_87 = 9'h57 == pht_ridx ? pht_87 : _GEN_86; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_88 = 9'h58 == pht_ridx ? pht_88 : _GEN_87; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_89 = 9'h59 == pht_ridx ? pht_89 : _GEN_88; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_90 = 9'h5a == pht_ridx ? pht_90 : _GEN_89; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_91 = 9'h5b == pht_ridx ? pht_91 : _GEN_90; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_92 = 9'h5c == pht_ridx ? pht_92 : _GEN_91; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_93 = 9'h5d == pht_ridx ? pht_93 : _GEN_92; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_94 = 9'h5e == pht_ridx ? pht_94 : _GEN_93; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_95 = 9'h5f == pht_ridx ? pht_95 : _GEN_94; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_96 = 9'h60 == pht_ridx ? pht_96 : _GEN_95; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_97 = 9'h61 == pht_ridx ? pht_97 : _GEN_96; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_98 = 9'h62 == pht_ridx ? pht_98 : _GEN_97; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_99 = 9'h63 == pht_ridx ? pht_99 : _GEN_98; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_100 = 9'h64 == pht_ridx ? pht_100 : _GEN_99; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_101 = 9'h65 == pht_ridx ? pht_101 : _GEN_100; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_102 = 9'h66 == pht_ridx ? pht_102 : _GEN_101; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_103 = 9'h67 == pht_ridx ? pht_103 : _GEN_102; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_104 = 9'h68 == pht_ridx ? pht_104 : _GEN_103; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_105 = 9'h69 == pht_ridx ? pht_105 : _GEN_104; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_106 = 9'h6a == pht_ridx ? pht_106 : _GEN_105; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_107 = 9'h6b == pht_ridx ? pht_107 : _GEN_106; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_108 = 9'h6c == pht_ridx ? pht_108 : _GEN_107; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_109 = 9'h6d == pht_ridx ? pht_109 : _GEN_108; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_110 = 9'h6e == pht_ridx ? pht_110 : _GEN_109; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_111 = 9'h6f == pht_ridx ? pht_111 : _GEN_110; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_112 = 9'h70 == pht_ridx ? pht_112 : _GEN_111; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_113 = 9'h71 == pht_ridx ? pht_113 : _GEN_112; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_114 = 9'h72 == pht_ridx ? pht_114 : _GEN_113; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_115 = 9'h73 == pht_ridx ? pht_115 : _GEN_114; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_116 = 9'h74 == pht_ridx ? pht_116 : _GEN_115; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_117 = 9'h75 == pht_ridx ? pht_117 : _GEN_116; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_118 = 9'h76 == pht_ridx ? pht_118 : _GEN_117; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_119 = 9'h77 == pht_ridx ? pht_119 : _GEN_118; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_120 = 9'h78 == pht_ridx ? pht_120 : _GEN_119; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_121 = 9'h79 == pht_ridx ? pht_121 : _GEN_120; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_122 = 9'h7a == pht_ridx ? pht_122 : _GEN_121; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_123 = 9'h7b == pht_ridx ? pht_123 : _GEN_122; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_124 = 9'h7c == pht_ridx ? pht_124 : _GEN_123; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_125 = 9'h7d == pht_ridx ? pht_125 : _GEN_124; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_126 = 9'h7e == pht_ridx ? pht_126 : _GEN_125; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_127 = 9'h7f == pht_ridx ? pht_127 : _GEN_126; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_128 = 9'h80 == pht_ridx ? pht_128 : _GEN_127; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_129 = 9'h81 == pht_ridx ? pht_129 : _GEN_128; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_130 = 9'h82 == pht_ridx ? pht_130 : _GEN_129; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_131 = 9'h83 == pht_ridx ? pht_131 : _GEN_130; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_132 = 9'h84 == pht_ridx ? pht_132 : _GEN_131; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_133 = 9'h85 == pht_ridx ? pht_133 : _GEN_132; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_134 = 9'h86 == pht_ridx ? pht_134 : _GEN_133; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_135 = 9'h87 == pht_ridx ? pht_135 : _GEN_134; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_136 = 9'h88 == pht_ridx ? pht_136 : _GEN_135; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_137 = 9'h89 == pht_ridx ? pht_137 : _GEN_136; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_138 = 9'h8a == pht_ridx ? pht_138 : _GEN_137; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_139 = 9'h8b == pht_ridx ? pht_139 : _GEN_138; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_140 = 9'h8c == pht_ridx ? pht_140 : _GEN_139; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_141 = 9'h8d == pht_ridx ? pht_141 : _GEN_140; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_142 = 9'h8e == pht_ridx ? pht_142 : _GEN_141; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_143 = 9'h8f == pht_ridx ? pht_143 : _GEN_142; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_144 = 9'h90 == pht_ridx ? pht_144 : _GEN_143; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_145 = 9'h91 == pht_ridx ? pht_145 : _GEN_144; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_146 = 9'h92 == pht_ridx ? pht_146 : _GEN_145; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_147 = 9'h93 == pht_ridx ? pht_147 : _GEN_146; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_148 = 9'h94 == pht_ridx ? pht_148 : _GEN_147; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_149 = 9'h95 == pht_ridx ? pht_149 : _GEN_148; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_150 = 9'h96 == pht_ridx ? pht_150 : _GEN_149; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_151 = 9'h97 == pht_ridx ? pht_151 : _GEN_150; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_152 = 9'h98 == pht_ridx ? pht_152 : _GEN_151; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_153 = 9'h99 == pht_ridx ? pht_153 : _GEN_152; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_154 = 9'h9a == pht_ridx ? pht_154 : _GEN_153; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_155 = 9'h9b == pht_ridx ? pht_155 : _GEN_154; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_156 = 9'h9c == pht_ridx ? pht_156 : _GEN_155; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_157 = 9'h9d == pht_ridx ? pht_157 : _GEN_156; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_158 = 9'h9e == pht_ridx ? pht_158 : _GEN_157; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_159 = 9'h9f == pht_ridx ? pht_159 : _GEN_158; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_160 = 9'ha0 == pht_ridx ? pht_160 : _GEN_159; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_161 = 9'ha1 == pht_ridx ? pht_161 : _GEN_160; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_162 = 9'ha2 == pht_ridx ? pht_162 : _GEN_161; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_163 = 9'ha3 == pht_ridx ? pht_163 : _GEN_162; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_164 = 9'ha4 == pht_ridx ? pht_164 : _GEN_163; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_165 = 9'ha5 == pht_ridx ? pht_165 : _GEN_164; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_166 = 9'ha6 == pht_ridx ? pht_166 : _GEN_165; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_167 = 9'ha7 == pht_ridx ? pht_167 : _GEN_166; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_168 = 9'ha8 == pht_ridx ? pht_168 : _GEN_167; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_169 = 9'ha9 == pht_ridx ? pht_169 : _GEN_168; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_170 = 9'haa == pht_ridx ? pht_170 : _GEN_169; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_171 = 9'hab == pht_ridx ? pht_171 : _GEN_170; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_172 = 9'hac == pht_ridx ? pht_172 : _GEN_171; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_173 = 9'had == pht_ridx ? pht_173 : _GEN_172; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_174 = 9'hae == pht_ridx ? pht_174 : _GEN_173; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_175 = 9'haf == pht_ridx ? pht_175 : _GEN_174; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_176 = 9'hb0 == pht_ridx ? pht_176 : _GEN_175; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_177 = 9'hb1 == pht_ridx ? pht_177 : _GEN_176; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_178 = 9'hb2 == pht_ridx ? pht_178 : _GEN_177; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_179 = 9'hb3 == pht_ridx ? pht_179 : _GEN_178; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_180 = 9'hb4 == pht_ridx ? pht_180 : _GEN_179; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_181 = 9'hb5 == pht_ridx ? pht_181 : _GEN_180; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_182 = 9'hb6 == pht_ridx ? pht_182 : _GEN_181; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_183 = 9'hb7 == pht_ridx ? pht_183 : _GEN_182; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_184 = 9'hb8 == pht_ridx ? pht_184 : _GEN_183; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_185 = 9'hb9 == pht_ridx ? pht_185 : _GEN_184; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_186 = 9'hba == pht_ridx ? pht_186 : _GEN_185; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_187 = 9'hbb == pht_ridx ? pht_187 : _GEN_186; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_188 = 9'hbc == pht_ridx ? pht_188 : _GEN_187; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_189 = 9'hbd == pht_ridx ? pht_189 : _GEN_188; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_190 = 9'hbe == pht_ridx ? pht_190 : _GEN_189; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_191 = 9'hbf == pht_ridx ? pht_191 : _GEN_190; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_192 = 9'hc0 == pht_ridx ? pht_192 : _GEN_191; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_193 = 9'hc1 == pht_ridx ? pht_193 : _GEN_192; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_194 = 9'hc2 == pht_ridx ? pht_194 : _GEN_193; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_195 = 9'hc3 == pht_ridx ? pht_195 : _GEN_194; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_196 = 9'hc4 == pht_ridx ? pht_196 : _GEN_195; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_197 = 9'hc5 == pht_ridx ? pht_197 : _GEN_196; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_198 = 9'hc6 == pht_ridx ? pht_198 : _GEN_197; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_199 = 9'hc7 == pht_ridx ? pht_199 : _GEN_198; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_200 = 9'hc8 == pht_ridx ? pht_200 : _GEN_199; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_201 = 9'hc9 == pht_ridx ? pht_201 : _GEN_200; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_202 = 9'hca == pht_ridx ? pht_202 : _GEN_201; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_203 = 9'hcb == pht_ridx ? pht_203 : _GEN_202; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_204 = 9'hcc == pht_ridx ? pht_204 : _GEN_203; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_205 = 9'hcd == pht_ridx ? pht_205 : _GEN_204; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_206 = 9'hce == pht_ridx ? pht_206 : _GEN_205; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_207 = 9'hcf == pht_ridx ? pht_207 : _GEN_206; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_208 = 9'hd0 == pht_ridx ? pht_208 : _GEN_207; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_209 = 9'hd1 == pht_ridx ? pht_209 : _GEN_208; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_210 = 9'hd2 == pht_ridx ? pht_210 : _GEN_209; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_211 = 9'hd3 == pht_ridx ? pht_211 : _GEN_210; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_212 = 9'hd4 == pht_ridx ? pht_212 : _GEN_211; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_213 = 9'hd5 == pht_ridx ? pht_213 : _GEN_212; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_214 = 9'hd6 == pht_ridx ? pht_214 : _GEN_213; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_215 = 9'hd7 == pht_ridx ? pht_215 : _GEN_214; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_216 = 9'hd8 == pht_ridx ? pht_216 : _GEN_215; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_217 = 9'hd9 == pht_ridx ? pht_217 : _GEN_216; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_218 = 9'hda == pht_ridx ? pht_218 : _GEN_217; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_219 = 9'hdb == pht_ridx ? pht_219 : _GEN_218; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_220 = 9'hdc == pht_ridx ? pht_220 : _GEN_219; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_221 = 9'hdd == pht_ridx ? pht_221 : _GEN_220; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_222 = 9'hde == pht_ridx ? pht_222 : _GEN_221; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_223 = 9'hdf == pht_ridx ? pht_223 : _GEN_222; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_224 = 9'he0 == pht_ridx ? pht_224 : _GEN_223; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_225 = 9'he1 == pht_ridx ? pht_225 : _GEN_224; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_226 = 9'he2 == pht_ridx ? pht_226 : _GEN_225; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_227 = 9'he3 == pht_ridx ? pht_227 : _GEN_226; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_228 = 9'he4 == pht_ridx ? pht_228 : _GEN_227; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_229 = 9'he5 == pht_ridx ? pht_229 : _GEN_228; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_230 = 9'he6 == pht_ridx ? pht_230 : _GEN_229; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_231 = 9'he7 == pht_ridx ? pht_231 : _GEN_230; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_232 = 9'he8 == pht_ridx ? pht_232 : _GEN_231; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_233 = 9'he9 == pht_ridx ? pht_233 : _GEN_232; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_234 = 9'hea == pht_ridx ? pht_234 : _GEN_233; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_235 = 9'heb == pht_ridx ? pht_235 : _GEN_234; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_236 = 9'hec == pht_ridx ? pht_236 : _GEN_235; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_237 = 9'hed == pht_ridx ? pht_237 : _GEN_236; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_238 = 9'hee == pht_ridx ? pht_238 : _GEN_237; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_239 = 9'hef == pht_ridx ? pht_239 : _GEN_238; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_240 = 9'hf0 == pht_ridx ? pht_240 : _GEN_239; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_241 = 9'hf1 == pht_ridx ? pht_241 : _GEN_240; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_242 = 9'hf2 == pht_ridx ? pht_242 : _GEN_241; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_243 = 9'hf3 == pht_ridx ? pht_243 : _GEN_242; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_244 = 9'hf4 == pht_ridx ? pht_244 : _GEN_243; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_245 = 9'hf5 == pht_ridx ? pht_245 : _GEN_244; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_246 = 9'hf6 == pht_ridx ? pht_246 : _GEN_245; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_247 = 9'hf7 == pht_ridx ? pht_247 : _GEN_246; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_248 = 9'hf8 == pht_ridx ? pht_248 : _GEN_247; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_249 = 9'hf9 == pht_ridx ? pht_249 : _GEN_248; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_250 = 9'hfa == pht_ridx ? pht_250 : _GEN_249; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_251 = 9'hfb == pht_ridx ? pht_251 : _GEN_250; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_252 = 9'hfc == pht_ridx ? pht_252 : _GEN_251; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_253 = 9'hfd == pht_ridx ? pht_253 : _GEN_252; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_254 = 9'hfe == pht_ridx ? pht_254 : _GEN_253; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_255 = 9'hff == pht_ridx ? pht_255 : _GEN_254; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_256 = 9'h100 == pht_ridx ? pht_256 : _GEN_255; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_257 = 9'h101 == pht_ridx ? pht_257 : _GEN_256; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_258 = 9'h102 == pht_ridx ? pht_258 : _GEN_257; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_259 = 9'h103 == pht_ridx ? pht_259 : _GEN_258; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_260 = 9'h104 == pht_ridx ? pht_260 : _GEN_259; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_261 = 9'h105 == pht_ridx ? pht_261 : _GEN_260; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_262 = 9'h106 == pht_ridx ? pht_262 : _GEN_261; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_263 = 9'h107 == pht_ridx ? pht_263 : _GEN_262; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_264 = 9'h108 == pht_ridx ? pht_264 : _GEN_263; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_265 = 9'h109 == pht_ridx ? pht_265 : _GEN_264; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_266 = 9'h10a == pht_ridx ? pht_266 : _GEN_265; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_267 = 9'h10b == pht_ridx ? pht_267 : _GEN_266; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_268 = 9'h10c == pht_ridx ? pht_268 : _GEN_267; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_269 = 9'h10d == pht_ridx ? pht_269 : _GEN_268; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_270 = 9'h10e == pht_ridx ? pht_270 : _GEN_269; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_271 = 9'h10f == pht_ridx ? pht_271 : _GEN_270; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_272 = 9'h110 == pht_ridx ? pht_272 : _GEN_271; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_273 = 9'h111 == pht_ridx ? pht_273 : _GEN_272; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_274 = 9'h112 == pht_ridx ? pht_274 : _GEN_273; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_275 = 9'h113 == pht_ridx ? pht_275 : _GEN_274; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_276 = 9'h114 == pht_ridx ? pht_276 : _GEN_275; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_277 = 9'h115 == pht_ridx ? pht_277 : _GEN_276; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_278 = 9'h116 == pht_ridx ? pht_278 : _GEN_277; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_279 = 9'h117 == pht_ridx ? pht_279 : _GEN_278; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_280 = 9'h118 == pht_ridx ? pht_280 : _GEN_279; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_281 = 9'h119 == pht_ridx ? pht_281 : _GEN_280; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_282 = 9'h11a == pht_ridx ? pht_282 : _GEN_281; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_283 = 9'h11b == pht_ridx ? pht_283 : _GEN_282; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_284 = 9'h11c == pht_ridx ? pht_284 : _GEN_283; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_285 = 9'h11d == pht_ridx ? pht_285 : _GEN_284; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_286 = 9'h11e == pht_ridx ? pht_286 : _GEN_285; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_287 = 9'h11f == pht_ridx ? pht_287 : _GEN_286; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_288 = 9'h120 == pht_ridx ? pht_288 : _GEN_287; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_289 = 9'h121 == pht_ridx ? pht_289 : _GEN_288; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_290 = 9'h122 == pht_ridx ? pht_290 : _GEN_289; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_291 = 9'h123 == pht_ridx ? pht_291 : _GEN_290; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_292 = 9'h124 == pht_ridx ? pht_292 : _GEN_291; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_293 = 9'h125 == pht_ridx ? pht_293 : _GEN_292; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_294 = 9'h126 == pht_ridx ? pht_294 : _GEN_293; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_295 = 9'h127 == pht_ridx ? pht_295 : _GEN_294; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_296 = 9'h128 == pht_ridx ? pht_296 : _GEN_295; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_297 = 9'h129 == pht_ridx ? pht_297 : _GEN_296; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_298 = 9'h12a == pht_ridx ? pht_298 : _GEN_297; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_299 = 9'h12b == pht_ridx ? pht_299 : _GEN_298; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_300 = 9'h12c == pht_ridx ? pht_300 : _GEN_299; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_301 = 9'h12d == pht_ridx ? pht_301 : _GEN_300; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_302 = 9'h12e == pht_ridx ? pht_302 : _GEN_301; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_303 = 9'h12f == pht_ridx ? pht_303 : _GEN_302; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_304 = 9'h130 == pht_ridx ? pht_304 : _GEN_303; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_305 = 9'h131 == pht_ridx ? pht_305 : _GEN_304; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_306 = 9'h132 == pht_ridx ? pht_306 : _GEN_305; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_307 = 9'h133 == pht_ridx ? pht_307 : _GEN_306; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_308 = 9'h134 == pht_ridx ? pht_308 : _GEN_307; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_309 = 9'h135 == pht_ridx ? pht_309 : _GEN_308; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_310 = 9'h136 == pht_ridx ? pht_310 : _GEN_309; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_311 = 9'h137 == pht_ridx ? pht_311 : _GEN_310; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_312 = 9'h138 == pht_ridx ? pht_312 : _GEN_311; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_313 = 9'h139 == pht_ridx ? pht_313 : _GEN_312; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_314 = 9'h13a == pht_ridx ? pht_314 : _GEN_313; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_315 = 9'h13b == pht_ridx ? pht_315 : _GEN_314; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_316 = 9'h13c == pht_ridx ? pht_316 : _GEN_315; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_317 = 9'h13d == pht_ridx ? pht_317 : _GEN_316; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_318 = 9'h13e == pht_ridx ? pht_318 : _GEN_317; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_319 = 9'h13f == pht_ridx ? pht_319 : _GEN_318; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_320 = 9'h140 == pht_ridx ? pht_320 : _GEN_319; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_321 = 9'h141 == pht_ridx ? pht_321 : _GEN_320; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_322 = 9'h142 == pht_ridx ? pht_322 : _GEN_321; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_323 = 9'h143 == pht_ridx ? pht_323 : _GEN_322; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_324 = 9'h144 == pht_ridx ? pht_324 : _GEN_323; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_325 = 9'h145 == pht_ridx ? pht_325 : _GEN_324; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_326 = 9'h146 == pht_ridx ? pht_326 : _GEN_325; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_327 = 9'h147 == pht_ridx ? pht_327 : _GEN_326; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_328 = 9'h148 == pht_ridx ? pht_328 : _GEN_327; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_329 = 9'h149 == pht_ridx ? pht_329 : _GEN_328; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_330 = 9'h14a == pht_ridx ? pht_330 : _GEN_329; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_331 = 9'h14b == pht_ridx ? pht_331 : _GEN_330; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_332 = 9'h14c == pht_ridx ? pht_332 : _GEN_331; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_333 = 9'h14d == pht_ridx ? pht_333 : _GEN_332; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_334 = 9'h14e == pht_ridx ? pht_334 : _GEN_333; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_335 = 9'h14f == pht_ridx ? pht_335 : _GEN_334; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_336 = 9'h150 == pht_ridx ? pht_336 : _GEN_335; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_337 = 9'h151 == pht_ridx ? pht_337 : _GEN_336; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_338 = 9'h152 == pht_ridx ? pht_338 : _GEN_337; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_339 = 9'h153 == pht_ridx ? pht_339 : _GEN_338; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_340 = 9'h154 == pht_ridx ? pht_340 : _GEN_339; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_341 = 9'h155 == pht_ridx ? pht_341 : _GEN_340; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_342 = 9'h156 == pht_ridx ? pht_342 : _GEN_341; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_343 = 9'h157 == pht_ridx ? pht_343 : _GEN_342; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_344 = 9'h158 == pht_ridx ? pht_344 : _GEN_343; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_345 = 9'h159 == pht_ridx ? pht_345 : _GEN_344; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_346 = 9'h15a == pht_ridx ? pht_346 : _GEN_345; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_347 = 9'h15b == pht_ridx ? pht_347 : _GEN_346; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_348 = 9'h15c == pht_ridx ? pht_348 : _GEN_347; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_349 = 9'h15d == pht_ridx ? pht_349 : _GEN_348; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_350 = 9'h15e == pht_ridx ? pht_350 : _GEN_349; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_351 = 9'h15f == pht_ridx ? pht_351 : _GEN_350; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_352 = 9'h160 == pht_ridx ? pht_352 : _GEN_351; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_353 = 9'h161 == pht_ridx ? pht_353 : _GEN_352; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_354 = 9'h162 == pht_ridx ? pht_354 : _GEN_353; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_355 = 9'h163 == pht_ridx ? pht_355 : _GEN_354; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_356 = 9'h164 == pht_ridx ? pht_356 : _GEN_355; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_357 = 9'h165 == pht_ridx ? pht_357 : _GEN_356; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_358 = 9'h166 == pht_ridx ? pht_358 : _GEN_357; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_359 = 9'h167 == pht_ridx ? pht_359 : _GEN_358; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_360 = 9'h168 == pht_ridx ? pht_360 : _GEN_359; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_361 = 9'h169 == pht_ridx ? pht_361 : _GEN_360; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_362 = 9'h16a == pht_ridx ? pht_362 : _GEN_361; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_363 = 9'h16b == pht_ridx ? pht_363 : _GEN_362; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_364 = 9'h16c == pht_ridx ? pht_364 : _GEN_363; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_365 = 9'h16d == pht_ridx ? pht_365 : _GEN_364; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_366 = 9'h16e == pht_ridx ? pht_366 : _GEN_365; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_367 = 9'h16f == pht_ridx ? pht_367 : _GEN_366; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_368 = 9'h170 == pht_ridx ? pht_368 : _GEN_367; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_369 = 9'h171 == pht_ridx ? pht_369 : _GEN_368; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_370 = 9'h172 == pht_ridx ? pht_370 : _GEN_369; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_371 = 9'h173 == pht_ridx ? pht_371 : _GEN_370; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_372 = 9'h174 == pht_ridx ? pht_372 : _GEN_371; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_373 = 9'h175 == pht_ridx ? pht_373 : _GEN_372; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_374 = 9'h176 == pht_ridx ? pht_374 : _GEN_373; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_375 = 9'h177 == pht_ridx ? pht_375 : _GEN_374; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_376 = 9'h178 == pht_ridx ? pht_376 : _GEN_375; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_377 = 9'h179 == pht_ridx ? pht_377 : _GEN_376; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_378 = 9'h17a == pht_ridx ? pht_378 : _GEN_377; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_379 = 9'h17b == pht_ridx ? pht_379 : _GEN_378; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_380 = 9'h17c == pht_ridx ? pht_380 : _GEN_379; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_381 = 9'h17d == pht_ridx ? pht_381 : _GEN_380; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_382 = 9'h17e == pht_ridx ? pht_382 : _GEN_381; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_383 = 9'h17f == pht_ridx ? pht_383 : _GEN_382; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_384 = 9'h180 == pht_ridx ? pht_384 : _GEN_383; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_385 = 9'h181 == pht_ridx ? pht_385 : _GEN_384; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_386 = 9'h182 == pht_ridx ? pht_386 : _GEN_385; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_387 = 9'h183 == pht_ridx ? pht_387 : _GEN_386; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_388 = 9'h184 == pht_ridx ? pht_388 : _GEN_387; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_389 = 9'h185 == pht_ridx ? pht_389 : _GEN_388; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_390 = 9'h186 == pht_ridx ? pht_390 : _GEN_389; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_391 = 9'h187 == pht_ridx ? pht_391 : _GEN_390; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_392 = 9'h188 == pht_ridx ? pht_392 : _GEN_391; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_393 = 9'h189 == pht_ridx ? pht_393 : _GEN_392; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_394 = 9'h18a == pht_ridx ? pht_394 : _GEN_393; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_395 = 9'h18b == pht_ridx ? pht_395 : _GEN_394; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_396 = 9'h18c == pht_ridx ? pht_396 : _GEN_395; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_397 = 9'h18d == pht_ridx ? pht_397 : _GEN_396; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_398 = 9'h18e == pht_ridx ? pht_398 : _GEN_397; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_399 = 9'h18f == pht_ridx ? pht_399 : _GEN_398; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_400 = 9'h190 == pht_ridx ? pht_400 : _GEN_399; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_401 = 9'h191 == pht_ridx ? pht_401 : _GEN_400; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_402 = 9'h192 == pht_ridx ? pht_402 : _GEN_401; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_403 = 9'h193 == pht_ridx ? pht_403 : _GEN_402; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_404 = 9'h194 == pht_ridx ? pht_404 : _GEN_403; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_405 = 9'h195 == pht_ridx ? pht_405 : _GEN_404; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_406 = 9'h196 == pht_ridx ? pht_406 : _GEN_405; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_407 = 9'h197 == pht_ridx ? pht_407 : _GEN_406; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_408 = 9'h198 == pht_ridx ? pht_408 : _GEN_407; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_409 = 9'h199 == pht_ridx ? pht_409 : _GEN_408; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_410 = 9'h19a == pht_ridx ? pht_410 : _GEN_409; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_411 = 9'h19b == pht_ridx ? pht_411 : _GEN_410; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_412 = 9'h19c == pht_ridx ? pht_412 : _GEN_411; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_413 = 9'h19d == pht_ridx ? pht_413 : _GEN_412; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_414 = 9'h19e == pht_ridx ? pht_414 : _GEN_413; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_415 = 9'h19f == pht_ridx ? pht_415 : _GEN_414; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_416 = 9'h1a0 == pht_ridx ? pht_416 : _GEN_415; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_417 = 9'h1a1 == pht_ridx ? pht_417 : _GEN_416; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_418 = 9'h1a2 == pht_ridx ? pht_418 : _GEN_417; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_419 = 9'h1a3 == pht_ridx ? pht_419 : _GEN_418; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_420 = 9'h1a4 == pht_ridx ? pht_420 : _GEN_419; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_421 = 9'h1a5 == pht_ridx ? pht_421 : _GEN_420; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_422 = 9'h1a6 == pht_ridx ? pht_422 : _GEN_421; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_423 = 9'h1a7 == pht_ridx ? pht_423 : _GEN_422; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_424 = 9'h1a8 == pht_ridx ? pht_424 : _GEN_423; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_425 = 9'h1a9 == pht_ridx ? pht_425 : _GEN_424; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_426 = 9'h1aa == pht_ridx ? pht_426 : _GEN_425; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_427 = 9'h1ab == pht_ridx ? pht_427 : _GEN_426; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_428 = 9'h1ac == pht_ridx ? pht_428 : _GEN_427; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_429 = 9'h1ad == pht_ridx ? pht_429 : _GEN_428; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_430 = 9'h1ae == pht_ridx ? pht_430 : _GEN_429; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_431 = 9'h1af == pht_ridx ? pht_431 : _GEN_430; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_432 = 9'h1b0 == pht_ridx ? pht_432 : _GEN_431; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_433 = 9'h1b1 == pht_ridx ? pht_433 : _GEN_432; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_434 = 9'h1b2 == pht_ridx ? pht_434 : _GEN_433; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_435 = 9'h1b3 == pht_ridx ? pht_435 : _GEN_434; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_436 = 9'h1b4 == pht_ridx ? pht_436 : _GEN_435; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_437 = 9'h1b5 == pht_ridx ? pht_437 : _GEN_436; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_438 = 9'h1b6 == pht_ridx ? pht_438 : _GEN_437; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_439 = 9'h1b7 == pht_ridx ? pht_439 : _GEN_438; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_440 = 9'h1b8 == pht_ridx ? pht_440 : _GEN_439; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_441 = 9'h1b9 == pht_ridx ? pht_441 : _GEN_440; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_442 = 9'h1ba == pht_ridx ? pht_442 : _GEN_441; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_443 = 9'h1bb == pht_ridx ? pht_443 : _GEN_442; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_444 = 9'h1bc == pht_ridx ? pht_444 : _GEN_443; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_445 = 9'h1bd == pht_ridx ? pht_445 : _GEN_444; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_446 = 9'h1be == pht_ridx ? pht_446 : _GEN_445; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_447 = 9'h1bf == pht_ridx ? pht_447 : _GEN_446; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_448 = 9'h1c0 == pht_ridx ? pht_448 : _GEN_447; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_449 = 9'h1c1 == pht_ridx ? pht_449 : _GEN_448; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_450 = 9'h1c2 == pht_ridx ? pht_450 : _GEN_449; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_451 = 9'h1c3 == pht_ridx ? pht_451 : _GEN_450; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_452 = 9'h1c4 == pht_ridx ? pht_452 : _GEN_451; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_453 = 9'h1c5 == pht_ridx ? pht_453 : _GEN_452; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_454 = 9'h1c6 == pht_ridx ? pht_454 : _GEN_453; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_455 = 9'h1c7 == pht_ridx ? pht_455 : _GEN_454; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_456 = 9'h1c8 == pht_ridx ? pht_456 : _GEN_455; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_457 = 9'h1c9 == pht_ridx ? pht_457 : _GEN_456; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_458 = 9'h1ca == pht_ridx ? pht_458 : _GEN_457; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_459 = 9'h1cb == pht_ridx ? pht_459 : _GEN_458; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_460 = 9'h1cc == pht_ridx ? pht_460 : _GEN_459; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_461 = 9'h1cd == pht_ridx ? pht_461 : _GEN_460; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_462 = 9'h1ce == pht_ridx ? pht_462 : _GEN_461; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_463 = 9'h1cf == pht_ridx ? pht_463 : _GEN_462; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_464 = 9'h1d0 == pht_ridx ? pht_464 : _GEN_463; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_465 = 9'h1d1 == pht_ridx ? pht_465 : _GEN_464; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_466 = 9'h1d2 == pht_ridx ? pht_466 : _GEN_465; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_467 = 9'h1d3 == pht_ridx ? pht_467 : _GEN_466; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_468 = 9'h1d4 == pht_ridx ? pht_468 : _GEN_467; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_469 = 9'h1d5 == pht_ridx ? pht_469 : _GEN_468; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_470 = 9'h1d6 == pht_ridx ? pht_470 : _GEN_469; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_471 = 9'h1d7 == pht_ridx ? pht_471 : _GEN_470; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_472 = 9'h1d8 == pht_ridx ? pht_472 : _GEN_471; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_473 = 9'h1d9 == pht_ridx ? pht_473 : _GEN_472; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_474 = 9'h1da == pht_ridx ? pht_474 : _GEN_473; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_475 = 9'h1db == pht_ridx ? pht_475 : _GEN_474; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_476 = 9'h1dc == pht_ridx ? pht_476 : _GEN_475; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_477 = 9'h1dd == pht_ridx ? pht_477 : _GEN_476; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_478 = 9'h1de == pht_ridx ? pht_478 : _GEN_477; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_479 = 9'h1df == pht_ridx ? pht_479 : _GEN_478; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_480 = 9'h1e0 == pht_ridx ? pht_480 : _GEN_479; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_481 = 9'h1e1 == pht_ridx ? pht_481 : _GEN_480; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_482 = 9'h1e2 == pht_ridx ? pht_482 : _GEN_481; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_483 = 9'h1e3 == pht_ridx ? pht_483 : _GEN_482; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_484 = 9'h1e4 == pht_ridx ? pht_484 : _GEN_483; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_485 = 9'h1e5 == pht_ridx ? pht_485 : _GEN_484; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_486 = 9'h1e6 == pht_ridx ? pht_486 : _GEN_485; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_487 = 9'h1e7 == pht_ridx ? pht_487 : _GEN_486; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_488 = 9'h1e8 == pht_ridx ? pht_488 : _GEN_487; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_489 = 9'h1e9 == pht_ridx ? pht_489 : _GEN_488; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_490 = 9'h1ea == pht_ridx ? pht_490 : _GEN_489; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_491 = 9'h1eb == pht_ridx ? pht_491 : _GEN_490; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_492 = 9'h1ec == pht_ridx ? pht_492 : _GEN_491; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_493 = 9'h1ed == pht_ridx ? pht_493 : _GEN_492; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_494 = 9'h1ee == pht_ridx ? pht_494 : _GEN_493; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_495 = 9'h1ef == pht_ridx ? pht_495 : _GEN_494; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_496 = 9'h1f0 == pht_ridx ? pht_496 : _GEN_495; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_497 = 9'h1f1 == pht_ridx ? pht_497 : _GEN_496; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_498 = 9'h1f2 == pht_ridx ? pht_498 : _GEN_497; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_499 = 9'h1f3 == pht_ridx ? pht_499 : _GEN_498; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_500 = 9'h1f4 == pht_ridx ? pht_500 : _GEN_499; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_501 = 9'h1f5 == pht_ridx ? pht_501 : _GEN_500; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_502 = 9'h1f6 == pht_ridx ? pht_502 : _GEN_501; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_503 = 9'h1f7 == pht_ridx ? pht_503 : _GEN_502; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_504 = 9'h1f8 == pht_ridx ? pht_504 : _GEN_503; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_505 = 9'h1f9 == pht_ridx ? pht_505 : _GEN_504; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_506 = 9'h1fa == pht_ridx ? pht_506 : _GEN_505; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_507 = 9'h1fb == pht_ridx ? pht_507 : _GEN_506; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_508 = 9'h1fc == pht_ridx ? pht_508 : _GEN_507; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_509 = 9'h1fd == pht_ridx ? pht_509 : _GEN_508; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_510 = 9'h1fe == pht_ridx ? pht_510 : _GEN_509; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_511 = 9'h1ff == pht_ridx ? pht_511 : _GEN_510; // @[BPU.scala 33:{30,30}]
  wire  pht_taken = _GEN_511 >= 2'h2; // @[BPU.scala 33:30]
  wire [36:0] _GEN_513 = btb_0_valid & btb_0_tag == io_pc[38:2] ? btb_0_target : 37'h0; // @[BPU.scala 39:67 41:17 37:30]
  wire [36:0] _GEN_515 = btb_1_valid & btb_1_tag == io_pc[38:2] ? btb_1_target : _GEN_513; // @[BPU.scala 39:67 41:17]
  wire [36:0] _GEN_517 = btb_2_valid & btb_2_tag == io_pc[38:2] ? btb_2_target : _GEN_515; // @[BPU.scala 39:67 41:17]
  wire [36:0] _GEN_519 = btb_3_valid & btb_3_tag == io_pc[38:2] ? btb_3_target : _GEN_517; // @[BPU.scala 39:67 41:17]
  wire [36:0] _GEN_521 = btb_4_valid & btb_4_tag == io_pc[38:2] ? btb_4_target : _GEN_519; // @[BPU.scala 39:67 41:17]
  wire [36:0] _GEN_523 = btb_5_valid & btb_5_tag == io_pc[38:2] ? btb_5_target : _GEN_521; // @[BPU.scala 39:67 41:17]
  wire [36:0] _GEN_525 = btb_6_valid & btb_6_tag == io_pc[38:2] ? btb_6_target : _GEN_523; // @[BPU.scala 39:67 41:17]
  wire [36:0] _GEN_527 = btb_7_valid & btb_7_tag == io_pc[38:2] ? btb_7_target : _GEN_525; // @[BPU.scala 39:67 41:17]
  wire [36:0] _GEN_529 = btb_8_valid & btb_8_tag == io_pc[38:2] ? btb_8_target : _GEN_527; // @[BPU.scala 39:67 41:17]
  wire  _GEN_530 = btb_9_valid & btb_9_tag == io_pc[38:2] | (btb_8_valid & btb_8_tag == io_pc[38:2] | (btb_7_valid &
    btb_7_tag == io_pc[38:2] | (btb_6_valid & btb_6_tag == io_pc[38:2] | (btb_5_valid & btb_5_tag == io_pc[38:2] | (
    btb_4_valid & btb_4_tag == io_pc[38:2] | (btb_3_valid & btb_3_tag == io_pc[38:2] | (btb_2_valid & btb_2_tag == io_pc
    [38:2] | (btb_1_valid & btb_1_tag == io_pc[38:2] | btb_0_valid & btb_0_tag == io_pc[38:2])))))))); // @[BPU.scala 39:67 40:17]
  wire [36:0] _GEN_531 = btb_9_valid & btb_9_tag == io_pc[38:2] ? btb_9_target : _GEN_529; // @[BPU.scala 39:67 41:17]
  wire [36:0] _GEN_533 = btb_10_valid & btb_10_tag == io_pc[38:2] ? btb_10_target : _GEN_531; // @[BPU.scala 39:67 41:17]
  wire [36:0] _GEN_535 = btb_11_valid & btb_11_tag == io_pc[38:2] ? btb_11_target : _GEN_533; // @[BPU.scala 39:67 41:17]
  wire [36:0] _GEN_537 = btb_12_valid & btb_12_tag == io_pc[38:2] ? btb_12_target : _GEN_535; // @[BPU.scala 39:67 41:17]
  wire [36:0] _GEN_539 = btb_13_valid & btb_13_tag == io_pc[38:2] ? btb_13_target : _GEN_537; // @[BPU.scala 39:67 41:17]
  wire [36:0] _GEN_541 = btb_14_valid & btb_14_tag == io_pc[38:2] ? btb_14_target : _GEN_539; // @[BPU.scala 39:67 41:17]
  wire  btb_rhit = btb_15_valid & btb_15_tag == io_pc[38:2] | (btb_14_valid & btb_14_tag == io_pc[38:2] | (btb_13_valid
     & btb_13_tag == io_pc[38:2] | (btb_12_valid & btb_12_tag == io_pc[38:2] | (btb_11_valid & btb_11_tag == io_pc[38:2]
     | (btb_10_valid & btb_10_tag == io_pc[38:2] | _GEN_530))))); // @[BPU.scala 39:67 40:17]
  wire [36:0] btb_rdata = btb_15_valid & btb_15_tag == io_pc[38:2] ? btb_15_target : _GEN_541; // @[BPU.scala 39:67 41:17]
  wire [63:0] _io_out_T_1 = io_pc + 64'h4; // @[BPU.scala 46:19]
  wire [38:0] _io_out_T_2 = {btb_rdata,2'h0}; // @[Cat.scala 33:92]
  wire [24:0] _io_out_T_5 = _io_out_T_2[38] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _io_out_T_6 = {_io_out_T_5,btb_rdata,2'h0}; // @[Cat.scala 33:92]
  wire [8:0] pht_widx = io_jmp_packet_bp_pc[10:2] ^ ghr; // @[BPU.scala 52:53]
  wire [7:0] _ghr_T_1 = {ghr[7:1],io_jmp_packet_bp_taken}; // @[Cat.scala 33:92]
  wire [1:0] _pht_T_1 = io_jmp_packet_bp_taken ? 2'h2 : 2'h0; // @[BPU.scala 60:19]
  wire [1:0] _pht_T_2 = io_jmp_packet_bp_taken ? 2'h3 : 2'h1; // @[BPU.scala 61:19]
  wire [1:0] _pht_T_3 = io_jmp_packet_bp_taken ? 2'h3 : 2'h2; // @[BPU.scala 62:19]
  wire [1:0] _GEN_546 = 9'h1 == pht_widx ? pht_1 : pht_0; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_547 = 9'h2 == pht_widx ? pht_2 : _GEN_546; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_548 = 9'h3 == pht_widx ? pht_3 : _GEN_547; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_549 = 9'h4 == pht_widx ? pht_4 : _GEN_548; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_550 = 9'h5 == pht_widx ? pht_5 : _GEN_549; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_551 = 9'h6 == pht_widx ? pht_6 : _GEN_550; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_552 = 9'h7 == pht_widx ? pht_7 : _GEN_551; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_553 = 9'h8 == pht_widx ? pht_8 : _GEN_552; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_554 = 9'h9 == pht_widx ? pht_9 : _GEN_553; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_555 = 9'ha == pht_widx ? pht_10 : _GEN_554; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_556 = 9'hb == pht_widx ? pht_11 : _GEN_555; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_557 = 9'hc == pht_widx ? pht_12 : _GEN_556; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_558 = 9'hd == pht_widx ? pht_13 : _GEN_557; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_559 = 9'he == pht_widx ? pht_14 : _GEN_558; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_560 = 9'hf == pht_widx ? pht_15 : _GEN_559; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_561 = 9'h10 == pht_widx ? pht_16 : _GEN_560; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_562 = 9'h11 == pht_widx ? pht_17 : _GEN_561; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_563 = 9'h12 == pht_widx ? pht_18 : _GEN_562; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_564 = 9'h13 == pht_widx ? pht_19 : _GEN_563; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_565 = 9'h14 == pht_widx ? pht_20 : _GEN_564; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_566 = 9'h15 == pht_widx ? pht_21 : _GEN_565; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_567 = 9'h16 == pht_widx ? pht_22 : _GEN_566; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_568 = 9'h17 == pht_widx ? pht_23 : _GEN_567; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_569 = 9'h18 == pht_widx ? pht_24 : _GEN_568; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_570 = 9'h19 == pht_widx ? pht_25 : _GEN_569; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_571 = 9'h1a == pht_widx ? pht_26 : _GEN_570; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_572 = 9'h1b == pht_widx ? pht_27 : _GEN_571; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_573 = 9'h1c == pht_widx ? pht_28 : _GEN_572; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_574 = 9'h1d == pht_widx ? pht_29 : _GEN_573; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_575 = 9'h1e == pht_widx ? pht_30 : _GEN_574; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_576 = 9'h1f == pht_widx ? pht_31 : _GEN_575; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_577 = 9'h20 == pht_widx ? pht_32 : _GEN_576; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_578 = 9'h21 == pht_widx ? pht_33 : _GEN_577; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_579 = 9'h22 == pht_widx ? pht_34 : _GEN_578; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_580 = 9'h23 == pht_widx ? pht_35 : _GEN_579; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_581 = 9'h24 == pht_widx ? pht_36 : _GEN_580; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_582 = 9'h25 == pht_widx ? pht_37 : _GEN_581; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_583 = 9'h26 == pht_widx ? pht_38 : _GEN_582; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_584 = 9'h27 == pht_widx ? pht_39 : _GEN_583; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_585 = 9'h28 == pht_widx ? pht_40 : _GEN_584; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_586 = 9'h29 == pht_widx ? pht_41 : _GEN_585; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_587 = 9'h2a == pht_widx ? pht_42 : _GEN_586; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_588 = 9'h2b == pht_widx ? pht_43 : _GEN_587; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_589 = 9'h2c == pht_widx ? pht_44 : _GEN_588; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_590 = 9'h2d == pht_widx ? pht_45 : _GEN_589; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_591 = 9'h2e == pht_widx ? pht_46 : _GEN_590; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_592 = 9'h2f == pht_widx ? pht_47 : _GEN_591; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_593 = 9'h30 == pht_widx ? pht_48 : _GEN_592; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_594 = 9'h31 == pht_widx ? pht_49 : _GEN_593; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_595 = 9'h32 == pht_widx ? pht_50 : _GEN_594; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_596 = 9'h33 == pht_widx ? pht_51 : _GEN_595; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_597 = 9'h34 == pht_widx ? pht_52 : _GEN_596; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_598 = 9'h35 == pht_widx ? pht_53 : _GEN_597; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_599 = 9'h36 == pht_widx ? pht_54 : _GEN_598; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_600 = 9'h37 == pht_widx ? pht_55 : _GEN_599; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_601 = 9'h38 == pht_widx ? pht_56 : _GEN_600; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_602 = 9'h39 == pht_widx ? pht_57 : _GEN_601; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_603 = 9'h3a == pht_widx ? pht_58 : _GEN_602; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_604 = 9'h3b == pht_widx ? pht_59 : _GEN_603; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_605 = 9'h3c == pht_widx ? pht_60 : _GEN_604; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_606 = 9'h3d == pht_widx ? pht_61 : _GEN_605; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_607 = 9'h3e == pht_widx ? pht_62 : _GEN_606; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_608 = 9'h3f == pht_widx ? pht_63 : _GEN_607; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_609 = 9'h40 == pht_widx ? pht_64 : _GEN_608; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_610 = 9'h41 == pht_widx ? pht_65 : _GEN_609; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_611 = 9'h42 == pht_widx ? pht_66 : _GEN_610; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_612 = 9'h43 == pht_widx ? pht_67 : _GEN_611; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_613 = 9'h44 == pht_widx ? pht_68 : _GEN_612; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_614 = 9'h45 == pht_widx ? pht_69 : _GEN_613; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_615 = 9'h46 == pht_widx ? pht_70 : _GEN_614; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_616 = 9'h47 == pht_widx ? pht_71 : _GEN_615; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_617 = 9'h48 == pht_widx ? pht_72 : _GEN_616; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_618 = 9'h49 == pht_widx ? pht_73 : _GEN_617; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_619 = 9'h4a == pht_widx ? pht_74 : _GEN_618; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_620 = 9'h4b == pht_widx ? pht_75 : _GEN_619; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_621 = 9'h4c == pht_widx ? pht_76 : _GEN_620; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_622 = 9'h4d == pht_widx ? pht_77 : _GEN_621; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_623 = 9'h4e == pht_widx ? pht_78 : _GEN_622; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_624 = 9'h4f == pht_widx ? pht_79 : _GEN_623; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_625 = 9'h50 == pht_widx ? pht_80 : _GEN_624; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_626 = 9'h51 == pht_widx ? pht_81 : _GEN_625; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_627 = 9'h52 == pht_widx ? pht_82 : _GEN_626; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_628 = 9'h53 == pht_widx ? pht_83 : _GEN_627; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_629 = 9'h54 == pht_widx ? pht_84 : _GEN_628; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_630 = 9'h55 == pht_widx ? pht_85 : _GEN_629; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_631 = 9'h56 == pht_widx ? pht_86 : _GEN_630; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_632 = 9'h57 == pht_widx ? pht_87 : _GEN_631; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_633 = 9'h58 == pht_widx ? pht_88 : _GEN_632; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_634 = 9'h59 == pht_widx ? pht_89 : _GEN_633; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_635 = 9'h5a == pht_widx ? pht_90 : _GEN_634; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_636 = 9'h5b == pht_widx ? pht_91 : _GEN_635; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_637 = 9'h5c == pht_widx ? pht_92 : _GEN_636; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_638 = 9'h5d == pht_widx ? pht_93 : _GEN_637; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_639 = 9'h5e == pht_widx ? pht_94 : _GEN_638; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_640 = 9'h5f == pht_widx ? pht_95 : _GEN_639; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_641 = 9'h60 == pht_widx ? pht_96 : _GEN_640; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_642 = 9'h61 == pht_widx ? pht_97 : _GEN_641; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_643 = 9'h62 == pht_widx ? pht_98 : _GEN_642; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_644 = 9'h63 == pht_widx ? pht_99 : _GEN_643; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_645 = 9'h64 == pht_widx ? pht_100 : _GEN_644; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_646 = 9'h65 == pht_widx ? pht_101 : _GEN_645; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_647 = 9'h66 == pht_widx ? pht_102 : _GEN_646; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_648 = 9'h67 == pht_widx ? pht_103 : _GEN_647; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_649 = 9'h68 == pht_widx ? pht_104 : _GEN_648; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_650 = 9'h69 == pht_widx ? pht_105 : _GEN_649; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_651 = 9'h6a == pht_widx ? pht_106 : _GEN_650; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_652 = 9'h6b == pht_widx ? pht_107 : _GEN_651; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_653 = 9'h6c == pht_widx ? pht_108 : _GEN_652; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_654 = 9'h6d == pht_widx ? pht_109 : _GEN_653; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_655 = 9'h6e == pht_widx ? pht_110 : _GEN_654; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_656 = 9'h6f == pht_widx ? pht_111 : _GEN_655; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_657 = 9'h70 == pht_widx ? pht_112 : _GEN_656; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_658 = 9'h71 == pht_widx ? pht_113 : _GEN_657; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_659 = 9'h72 == pht_widx ? pht_114 : _GEN_658; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_660 = 9'h73 == pht_widx ? pht_115 : _GEN_659; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_661 = 9'h74 == pht_widx ? pht_116 : _GEN_660; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_662 = 9'h75 == pht_widx ? pht_117 : _GEN_661; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_663 = 9'h76 == pht_widx ? pht_118 : _GEN_662; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_664 = 9'h77 == pht_widx ? pht_119 : _GEN_663; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_665 = 9'h78 == pht_widx ? pht_120 : _GEN_664; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_666 = 9'h79 == pht_widx ? pht_121 : _GEN_665; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_667 = 9'h7a == pht_widx ? pht_122 : _GEN_666; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_668 = 9'h7b == pht_widx ? pht_123 : _GEN_667; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_669 = 9'h7c == pht_widx ? pht_124 : _GEN_668; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_670 = 9'h7d == pht_widx ? pht_125 : _GEN_669; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_671 = 9'h7e == pht_widx ? pht_126 : _GEN_670; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_672 = 9'h7f == pht_widx ? pht_127 : _GEN_671; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_673 = 9'h80 == pht_widx ? pht_128 : _GEN_672; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_674 = 9'h81 == pht_widx ? pht_129 : _GEN_673; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_675 = 9'h82 == pht_widx ? pht_130 : _GEN_674; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_676 = 9'h83 == pht_widx ? pht_131 : _GEN_675; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_677 = 9'h84 == pht_widx ? pht_132 : _GEN_676; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_678 = 9'h85 == pht_widx ? pht_133 : _GEN_677; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_679 = 9'h86 == pht_widx ? pht_134 : _GEN_678; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_680 = 9'h87 == pht_widx ? pht_135 : _GEN_679; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_681 = 9'h88 == pht_widx ? pht_136 : _GEN_680; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_682 = 9'h89 == pht_widx ? pht_137 : _GEN_681; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_683 = 9'h8a == pht_widx ? pht_138 : _GEN_682; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_684 = 9'h8b == pht_widx ? pht_139 : _GEN_683; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_685 = 9'h8c == pht_widx ? pht_140 : _GEN_684; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_686 = 9'h8d == pht_widx ? pht_141 : _GEN_685; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_687 = 9'h8e == pht_widx ? pht_142 : _GEN_686; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_688 = 9'h8f == pht_widx ? pht_143 : _GEN_687; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_689 = 9'h90 == pht_widx ? pht_144 : _GEN_688; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_690 = 9'h91 == pht_widx ? pht_145 : _GEN_689; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_691 = 9'h92 == pht_widx ? pht_146 : _GEN_690; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_692 = 9'h93 == pht_widx ? pht_147 : _GEN_691; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_693 = 9'h94 == pht_widx ? pht_148 : _GEN_692; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_694 = 9'h95 == pht_widx ? pht_149 : _GEN_693; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_695 = 9'h96 == pht_widx ? pht_150 : _GEN_694; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_696 = 9'h97 == pht_widx ? pht_151 : _GEN_695; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_697 = 9'h98 == pht_widx ? pht_152 : _GEN_696; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_698 = 9'h99 == pht_widx ? pht_153 : _GEN_697; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_699 = 9'h9a == pht_widx ? pht_154 : _GEN_698; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_700 = 9'h9b == pht_widx ? pht_155 : _GEN_699; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_701 = 9'h9c == pht_widx ? pht_156 : _GEN_700; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_702 = 9'h9d == pht_widx ? pht_157 : _GEN_701; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_703 = 9'h9e == pht_widx ? pht_158 : _GEN_702; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_704 = 9'h9f == pht_widx ? pht_159 : _GEN_703; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_705 = 9'ha0 == pht_widx ? pht_160 : _GEN_704; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_706 = 9'ha1 == pht_widx ? pht_161 : _GEN_705; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_707 = 9'ha2 == pht_widx ? pht_162 : _GEN_706; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_708 = 9'ha3 == pht_widx ? pht_163 : _GEN_707; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_709 = 9'ha4 == pht_widx ? pht_164 : _GEN_708; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_710 = 9'ha5 == pht_widx ? pht_165 : _GEN_709; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_711 = 9'ha6 == pht_widx ? pht_166 : _GEN_710; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_712 = 9'ha7 == pht_widx ? pht_167 : _GEN_711; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_713 = 9'ha8 == pht_widx ? pht_168 : _GEN_712; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_714 = 9'ha9 == pht_widx ? pht_169 : _GEN_713; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_715 = 9'haa == pht_widx ? pht_170 : _GEN_714; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_716 = 9'hab == pht_widx ? pht_171 : _GEN_715; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_717 = 9'hac == pht_widx ? pht_172 : _GEN_716; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_718 = 9'had == pht_widx ? pht_173 : _GEN_717; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_719 = 9'hae == pht_widx ? pht_174 : _GEN_718; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_720 = 9'haf == pht_widx ? pht_175 : _GEN_719; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_721 = 9'hb0 == pht_widx ? pht_176 : _GEN_720; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_722 = 9'hb1 == pht_widx ? pht_177 : _GEN_721; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_723 = 9'hb2 == pht_widx ? pht_178 : _GEN_722; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_724 = 9'hb3 == pht_widx ? pht_179 : _GEN_723; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_725 = 9'hb4 == pht_widx ? pht_180 : _GEN_724; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_726 = 9'hb5 == pht_widx ? pht_181 : _GEN_725; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_727 = 9'hb6 == pht_widx ? pht_182 : _GEN_726; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_728 = 9'hb7 == pht_widx ? pht_183 : _GEN_727; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_729 = 9'hb8 == pht_widx ? pht_184 : _GEN_728; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_730 = 9'hb9 == pht_widx ? pht_185 : _GEN_729; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_731 = 9'hba == pht_widx ? pht_186 : _GEN_730; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_732 = 9'hbb == pht_widx ? pht_187 : _GEN_731; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_733 = 9'hbc == pht_widx ? pht_188 : _GEN_732; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_734 = 9'hbd == pht_widx ? pht_189 : _GEN_733; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_735 = 9'hbe == pht_widx ? pht_190 : _GEN_734; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_736 = 9'hbf == pht_widx ? pht_191 : _GEN_735; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_737 = 9'hc0 == pht_widx ? pht_192 : _GEN_736; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_738 = 9'hc1 == pht_widx ? pht_193 : _GEN_737; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_739 = 9'hc2 == pht_widx ? pht_194 : _GEN_738; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_740 = 9'hc3 == pht_widx ? pht_195 : _GEN_739; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_741 = 9'hc4 == pht_widx ? pht_196 : _GEN_740; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_742 = 9'hc5 == pht_widx ? pht_197 : _GEN_741; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_743 = 9'hc6 == pht_widx ? pht_198 : _GEN_742; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_744 = 9'hc7 == pht_widx ? pht_199 : _GEN_743; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_745 = 9'hc8 == pht_widx ? pht_200 : _GEN_744; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_746 = 9'hc9 == pht_widx ? pht_201 : _GEN_745; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_747 = 9'hca == pht_widx ? pht_202 : _GEN_746; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_748 = 9'hcb == pht_widx ? pht_203 : _GEN_747; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_749 = 9'hcc == pht_widx ? pht_204 : _GEN_748; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_750 = 9'hcd == pht_widx ? pht_205 : _GEN_749; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_751 = 9'hce == pht_widx ? pht_206 : _GEN_750; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_752 = 9'hcf == pht_widx ? pht_207 : _GEN_751; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_753 = 9'hd0 == pht_widx ? pht_208 : _GEN_752; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_754 = 9'hd1 == pht_widx ? pht_209 : _GEN_753; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_755 = 9'hd2 == pht_widx ? pht_210 : _GEN_754; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_756 = 9'hd3 == pht_widx ? pht_211 : _GEN_755; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_757 = 9'hd4 == pht_widx ? pht_212 : _GEN_756; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_758 = 9'hd5 == pht_widx ? pht_213 : _GEN_757; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_759 = 9'hd6 == pht_widx ? pht_214 : _GEN_758; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_760 = 9'hd7 == pht_widx ? pht_215 : _GEN_759; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_761 = 9'hd8 == pht_widx ? pht_216 : _GEN_760; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_762 = 9'hd9 == pht_widx ? pht_217 : _GEN_761; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_763 = 9'hda == pht_widx ? pht_218 : _GEN_762; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_764 = 9'hdb == pht_widx ? pht_219 : _GEN_763; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_765 = 9'hdc == pht_widx ? pht_220 : _GEN_764; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_766 = 9'hdd == pht_widx ? pht_221 : _GEN_765; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_767 = 9'hde == pht_widx ? pht_222 : _GEN_766; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_768 = 9'hdf == pht_widx ? pht_223 : _GEN_767; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_769 = 9'he0 == pht_widx ? pht_224 : _GEN_768; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_770 = 9'he1 == pht_widx ? pht_225 : _GEN_769; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_771 = 9'he2 == pht_widx ? pht_226 : _GEN_770; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_772 = 9'he3 == pht_widx ? pht_227 : _GEN_771; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_773 = 9'he4 == pht_widx ? pht_228 : _GEN_772; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_774 = 9'he5 == pht_widx ? pht_229 : _GEN_773; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_775 = 9'he6 == pht_widx ? pht_230 : _GEN_774; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_776 = 9'he7 == pht_widx ? pht_231 : _GEN_775; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_777 = 9'he8 == pht_widx ? pht_232 : _GEN_776; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_778 = 9'he9 == pht_widx ? pht_233 : _GEN_777; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_779 = 9'hea == pht_widx ? pht_234 : _GEN_778; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_780 = 9'heb == pht_widx ? pht_235 : _GEN_779; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_781 = 9'hec == pht_widx ? pht_236 : _GEN_780; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_782 = 9'hed == pht_widx ? pht_237 : _GEN_781; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_783 = 9'hee == pht_widx ? pht_238 : _GEN_782; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_784 = 9'hef == pht_widx ? pht_239 : _GEN_783; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_785 = 9'hf0 == pht_widx ? pht_240 : _GEN_784; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_786 = 9'hf1 == pht_widx ? pht_241 : _GEN_785; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_787 = 9'hf2 == pht_widx ? pht_242 : _GEN_786; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_788 = 9'hf3 == pht_widx ? pht_243 : _GEN_787; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_789 = 9'hf4 == pht_widx ? pht_244 : _GEN_788; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_790 = 9'hf5 == pht_widx ? pht_245 : _GEN_789; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_791 = 9'hf6 == pht_widx ? pht_246 : _GEN_790; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_792 = 9'hf7 == pht_widx ? pht_247 : _GEN_791; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_793 = 9'hf8 == pht_widx ? pht_248 : _GEN_792; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_794 = 9'hf9 == pht_widx ? pht_249 : _GEN_793; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_795 = 9'hfa == pht_widx ? pht_250 : _GEN_794; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_796 = 9'hfb == pht_widx ? pht_251 : _GEN_795; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_797 = 9'hfc == pht_widx ? pht_252 : _GEN_796; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_798 = 9'hfd == pht_widx ? pht_253 : _GEN_797; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_799 = 9'hfe == pht_widx ? pht_254 : _GEN_798; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_800 = 9'hff == pht_widx ? pht_255 : _GEN_799; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_801 = 9'h100 == pht_widx ? pht_256 : _GEN_800; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_802 = 9'h101 == pht_widx ? pht_257 : _GEN_801; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_803 = 9'h102 == pht_widx ? pht_258 : _GEN_802; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_804 = 9'h103 == pht_widx ? pht_259 : _GEN_803; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_805 = 9'h104 == pht_widx ? pht_260 : _GEN_804; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_806 = 9'h105 == pht_widx ? pht_261 : _GEN_805; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_807 = 9'h106 == pht_widx ? pht_262 : _GEN_806; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_808 = 9'h107 == pht_widx ? pht_263 : _GEN_807; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_809 = 9'h108 == pht_widx ? pht_264 : _GEN_808; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_810 = 9'h109 == pht_widx ? pht_265 : _GEN_809; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_811 = 9'h10a == pht_widx ? pht_266 : _GEN_810; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_812 = 9'h10b == pht_widx ? pht_267 : _GEN_811; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_813 = 9'h10c == pht_widx ? pht_268 : _GEN_812; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_814 = 9'h10d == pht_widx ? pht_269 : _GEN_813; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_815 = 9'h10e == pht_widx ? pht_270 : _GEN_814; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_816 = 9'h10f == pht_widx ? pht_271 : _GEN_815; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_817 = 9'h110 == pht_widx ? pht_272 : _GEN_816; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_818 = 9'h111 == pht_widx ? pht_273 : _GEN_817; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_819 = 9'h112 == pht_widx ? pht_274 : _GEN_818; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_820 = 9'h113 == pht_widx ? pht_275 : _GEN_819; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_821 = 9'h114 == pht_widx ? pht_276 : _GEN_820; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_822 = 9'h115 == pht_widx ? pht_277 : _GEN_821; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_823 = 9'h116 == pht_widx ? pht_278 : _GEN_822; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_824 = 9'h117 == pht_widx ? pht_279 : _GEN_823; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_825 = 9'h118 == pht_widx ? pht_280 : _GEN_824; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_826 = 9'h119 == pht_widx ? pht_281 : _GEN_825; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_827 = 9'h11a == pht_widx ? pht_282 : _GEN_826; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_828 = 9'h11b == pht_widx ? pht_283 : _GEN_827; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_829 = 9'h11c == pht_widx ? pht_284 : _GEN_828; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_830 = 9'h11d == pht_widx ? pht_285 : _GEN_829; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_831 = 9'h11e == pht_widx ? pht_286 : _GEN_830; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_832 = 9'h11f == pht_widx ? pht_287 : _GEN_831; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_833 = 9'h120 == pht_widx ? pht_288 : _GEN_832; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_834 = 9'h121 == pht_widx ? pht_289 : _GEN_833; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_835 = 9'h122 == pht_widx ? pht_290 : _GEN_834; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_836 = 9'h123 == pht_widx ? pht_291 : _GEN_835; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_837 = 9'h124 == pht_widx ? pht_292 : _GEN_836; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_838 = 9'h125 == pht_widx ? pht_293 : _GEN_837; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_839 = 9'h126 == pht_widx ? pht_294 : _GEN_838; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_840 = 9'h127 == pht_widx ? pht_295 : _GEN_839; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_841 = 9'h128 == pht_widx ? pht_296 : _GEN_840; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_842 = 9'h129 == pht_widx ? pht_297 : _GEN_841; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_843 = 9'h12a == pht_widx ? pht_298 : _GEN_842; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_844 = 9'h12b == pht_widx ? pht_299 : _GEN_843; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_845 = 9'h12c == pht_widx ? pht_300 : _GEN_844; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_846 = 9'h12d == pht_widx ? pht_301 : _GEN_845; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_847 = 9'h12e == pht_widx ? pht_302 : _GEN_846; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_848 = 9'h12f == pht_widx ? pht_303 : _GEN_847; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_849 = 9'h130 == pht_widx ? pht_304 : _GEN_848; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_850 = 9'h131 == pht_widx ? pht_305 : _GEN_849; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_851 = 9'h132 == pht_widx ? pht_306 : _GEN_850; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_852 = 9'h133 == pht_widx ? pht_307 : _GEN_851; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_853 = 9'h134 == pht_widx ? pht_308 : _GEN_852; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_854 = 9'h135 == pht_widx ? pht_309 : _GEN_853; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_855 = 9'h136 == pht_widx ? pht_310 : _GEN_854; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_856 = 9'h137 == pht_widx ? pht_311 : _GEN_855; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_857 = 9'h138 == pht_widx ? pht_312 : _GEN_856; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_858 = 9'h139 == pht_widx ? pht_313 : _GEN_857; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_859 = 9'h13a == pht_widx ? pht_314 : _GEN_858; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_860 = 9'h13b == pht_widx ? pht_315 : _GEN_859; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_861 = 9'h13c == pht_widx ? pht_316 : _GEN_860; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_862 = 9'h13d == pht_widx ? pht_317 : _GEN_861; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_863 = 9'h13e == pht_widx ? pht_318 : _GEN_862; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_864 = 9'h13f == pht_widx ? pht_319 : _GEN_863; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_865 = 9'h140 == pht_widx ? pht_320 : _GEN_864; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_866 = 9'h141 == pht_widx ? pht_321 : _GEN_865; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_867 = 9'h142 == pht_widx ? pht_322 : _GEN_866; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_868 = 9'h143 == pht_widx ? pht_323 : _GEN_867; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_869 = 9'h144 == pht_widx ? pht_324 : _GEN_868; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_870 = 9'h145 == pht_widx ? pht_325 : _GEN_869; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_871 = 9'h146 == pht_widx ? pht_326 : _GEN_870; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_872 = 9'h147 == pht_widx ? pht_327 : _GEN_871; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_873 = 9'h148 == pht_widx ? pht_328 : _GEN_872; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_874 = 9'h149 == pht_widx ? pht_329 : _GEN_873; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_875 = 9'h14a == pht_widx ? pht_330 : _GEN_874; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_876 = 9'h14b == pht_widx ? pht_331 : _GEN_875; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_877 = 9'h14c == pht_widx ? pht_332 : _GEN_876; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_878 = 9'h14d == pht_widx ? pht_333 : _GEN_877; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_879 = 9'h14e == pht_widx ? pht_334 : _GEN_878; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_880 = 9'h14f == pht_widx ? pht_335 : _GEN_879; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_881 = 9'h150 == pht_widx ? pht_336 : _GEN_880; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_882 = 9'h151 == pht_widx ? pht_337 : _GEN_881; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_883 = 9'h152 == pht_widx ? pht_338 : _GEN_882; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_884 = 9'h153 == pht_widx ? pht_339 : _GEN_883; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_885 = 9'h154 == pht_widx ? pht_340 : _GEN_884; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_886 = 9'h155 == pht_widx ? pht_341 : _GEN_885; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_887 = 9'h156 == pht_widx ? pht_342 : _GEN_886; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_888 = 9'h157 == pht_widx ? pht_343 : _GEN_887; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_889 = 9'h158 == pht_widx ? pht_344 : _GEN_888; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_890 = 9'h159 == pht_widx ? pht_345 : _GEN_889; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_891 = 9'h15a == pht_widx ? pht_346 : _GEN_890; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_892 = 9'h15b == pht_widx ? pht_347 : _GEN_891; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_893 = 9'h15c == pht_widx ? pht_348 : _GEN_892; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_894 = 9'h15d == pht_widx ? pht_349 : _GEN_893; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_895 = 9'h15e == pht_widx ? pht_350 : _GEN_894; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_896 = 9'h15f == pht_widx ? pht_351 : _GEN_895; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_897 = 9'h160 == pht_widx ? pht_352 : _GEN_896; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_898 = 9'h161 == pht_widx ? pht_353 : _GEN_897; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_899 = 9'h162 == pht_widx ? pht_354 : _GEN_898; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_900 = 9'h163 == pht_widx ? pht_355 : _GEN_899; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_901 = 9'h164 == pht_widx ? pht_356 : _GEN_900; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_902 = 9'h165 == pht_widx ? pht_357 : _GEN_901; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_903 = 9'h166 == pht_widx ? pht_358 : _GEN_902; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_904 = 9'h167 == pht_widx ? pht_359 : _GEN_903; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_905 = 9'h168 == pht_widx ? pht_360 : _GEN_904; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_906 = 9'h169 == pht_widx ? pht_361 : _GEN_905; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_907 = 9'h16a == pht_widx ? pht_362 : _GEN_906; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_908 = 9'h16b == pht_widx ? pht_363 : _GEN_907; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_909 = 9'h16c == pht_widx ? pht_364 : _GEN_908; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_910 = 9'h16d == pht_widx ? pht_365 : _GEN_909; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_911 = 9'h16e == pht_widx ? pht_366 : _GEN_910; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_912 = 9'h16f == pht_widx ? pht_367 : _GEN_911; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_913 = 9'h170 == pht_widx ? pht_368 : _GEN_912; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_914 = 9'h171 == pht_widx ? pht_369 : _GEN_913; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_915 = 9'h172 == pht_widx ? pht_370 : _GEN_914; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_916 = 9'h173 == pht_widx ? pht_371 : _GEN_915; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_917 = 9'h174 == pht_widx ? pht_372 : _GEN_916; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_918 = 9'h175 == pht_widx ? pht_373 : _GEN_917; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_919 = 9'h176 == pht_widx ? pht_374 : _GEN_918; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_920 = 9'h177 == pht_widx ? pht_375 : _GEN_919; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_921 = 9'h178 == pht_widx ? pht_376 : _GEN_920; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_922 = 9'h179 == pht_widx ? pht_377 : _GEN_921; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_923 = 9'h17a == pht_widx ? pht_378 : _GEN_922; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_924 = 9'h17b == pht_widx ? pht_379 : _GEN_923; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_925 = 9'h17c == pht_widx ? pht_380 : _GEN_924; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_926 = 9'h17d == pht_widx ? pht_381 : _GEN_925; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_927 = 9'h17e == pht_widx ? pht_382 : _GEN_926; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_928 = 9'h17f == pht_widx ? pht_383 : _GEN_927; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_929 = 9'h180 == pht_widx ? pht_384 : _GEN_928; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_930 = 9'h181 == pht_widx ? pht_385 : _GEN_929; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_931 = 9'h182 == pht_widx ? pht_386 : _GEN_930; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_932 = 9'h183 == pht_widx ? pht_387 : _GEN_931; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_933 = 9'h184 == pht_widx ? pht_388 : _GEN_932; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_934 = 9'h185 == pht_widx ? pht_389 : _GEN_933; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_935 = 9'h186 == pht_widx ? pht_390 : _GEN_934; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_936 = 9'h187 == pht_widx ? pht_391 : _GEN_935; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_937 = 9'h188 == pht_widx ? pht_392 : _GEN_936; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_938 = 9'h189 == pht_widx ? pht_393 : _GEN_937; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_939 = 9'h18a == pht_widx ? pht_394 : _GEN_938; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_940 = 9'h18b == pht_widx ? pht_395 : _GEN_939; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_941 = 9'h18c == pht_widx ? pht_396 : _GEN_940; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_942 = 9'h18d == pht_widx ? pht_397 : _GEN_941; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_943 = 9'h18e == pht_widx ? pht_398 : _GEN_942; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_944 = 9'h18f == pht_widx ? pht_399 : _GEN_943; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_945 = 9'h190 == pht_widx ? pht_400 : _GEN_944; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_946 = 9'h191 == pht_widx ? pht_401 : _GEN_945; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_947 = 9'h192 == pht_widx ? pht_402 : _GEN_946; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_948 = 9'h193 == pht_widx ? pht_403 : _GEN_947; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_949 = 9'h194 == pht_widx ? pht_404 : _GEN_948; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_950 = 9'h195 == pht_widx ? pht_405 : _GEN_949; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_951 = 9'h196 == pht_widx ? pht_406 : _GEN_950; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_952 = 9'h197 == pht_widx ? pht_407 : _GEN_951; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_953 = 9'h198 == pht_widx ? pht_408 : _GEN_952; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_954 = 9'h199 == pht_widx ? pht_409 : _GEN_953; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_955 = 9'h19a == pht_widx ? pht_410 : _GEN_954; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_956 = 9'h19b == pht_widx ? pht_411 : _GEN_955; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_957 = 9'h19c == pht_widx ? pht_412 : _GEN_956; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_958 = 9'h19d == pht_widx ? pht_413 : _GEN_957; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_959 = 9'h19e == pht_widx ? pht_414 : _GEN_958; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_960 = 9'h19f == pht_widx ? pht_415 : _GEN_959; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_961 = 9'h1a0 == pht_widx ? pht_416 : _GEN_960; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_962 = 9'h1a1 == pht_widx ? pht_417 : _GEN_961; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_963 = 9'h1a2 == pht_widx ? pht_418 : _GEN_962; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_964 = 9'h1a3 == pht_widx ? pht_419 : _GEN_963; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_965 = 9'h1a4 == pht_widx ? pht_420 : _GEN_964; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_966 = 9'h1a5 == pht_widx ? pht_421 : _GEN_965; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_967 = 9'h1a6 == pht_widx ? pht_422 : _GEN_966; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_968 = 9'h1a7 == pht_widx ? pht_423 : _GEN_967; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_969 = 9'h1a8 == pht_widx ? pht_424 : _GEN_968; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_970 = 9'h1a9 == pht_widx ? pht_425 : _GEN_969; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_971 = 9'h1aa == pht_widx ? pht_426 : _GEN_970; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_972 = 9'h1ab == pht_widx ? pht_427 : _GEN_971; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_973 = 9'h1ac == pht_widx ? pht_428 : _GEN_972; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_974 = 9'h1ad == pht_widx ? pht_429 : _GEN_973; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_975 = 9'h1ae == pht_widx ? pht_430 : _GEN_974; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_976 = 9'h1af == pht_widx ? pht_431 : _GEN_975; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_977 = 9'h1b0 == pht_widx ? pht_432 : _GEN_976; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_978 = 9'h1b1 == pht_widx ? pht_433 : _GEN_977; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_979 = 9'h1b2 == pht_widx ? pht_434 : _GEN_978; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_980 = 9'h1b3 == pht_widx ? pht_435 : _GEN_979; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_981 = 9'h1b4 == pht_widx ? pht_436 : _GEN_980; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_982 = 9'h1b5 == pht_widx ? pht_437 : _GEN_981; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_983 = 9'h1b6 == pht_widx ? pht_438 : _GEN_982; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_984 = 9'h1b7 == pht_widx ? pht_439 : _GEN_983; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_985 = 9'h1b8 == pht_widx ? pht_440 : _GEN_984; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_986 = 9'h1b9 == pht_widx ? pht_441 : _GEN_985; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_987 = 9'h1ba == pht_widx ? pht_442 : _GEN_986; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_988 = 9'h1bb == pht_widx ? pht_443 : _GEN_987; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_989 = 9'h1bc == pht_widx ? pht_444 : _GEN_988; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_990 = 9'h1bd == pht_widx ? pht_445 : _GEN_989; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_991 = 9'h1be == pht_widx ? pht_446 : _GEN_990; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_992 = 9'h1bf == pht_widx ? pht_447 : _GEN_991; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_993 = 9'h1c0 == pht_widx ? pht_448 : _GEN_992; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_994 = 9'h1c1 == pht_widx ? pht_449 : _GEN_993; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_995 = 9'h1c2 == pht_widx ? pht_450 : _GEN_994; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_996 = 9'h1c3 == pht_widx ? pht_451 : _GEN_995; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_997 = 9'h1c4 == pht_widx ? pht_452 : _GEN_996; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_998 = 9'h1c5 == pht_widx ? pht_453 : _GEN_997; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_999 = 9'h1c6 == pht_widx ? pht_454 : _GEN_998; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1000 = 9'h1c7 == pht_widx ? pht_455 : _GEN_999; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1001 = 9'h1c8 == pht_widx ? pht_456 : _GEN_1000; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1002 = 9'h1c9 == pht_widx ? pht_457 : _GEN_1001; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1003 = 9'h1ca == pht_widx ? pht_458 : _GEN_1002; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1004 = 9'h1cb == pht_widx ? pht_459 : _GEN_1003; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1005 = 9'h1cc == pht_widx ? pht_460 : _GEN_1004; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1006 = 9'h1cd == pht_widx ? pht_461 : _GEN_1005; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1007 = 9'h1ce == pht_widx ? pht_462 : _GEN_1006; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1008 = 9'h1cf == pht_widx ? pht_463 : _GEN_1007; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1009 = 9'h1d0 == pht_widx ? pht_464 : _GEN_1008; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1010 = 9'h1d1 == pht_widx ? pht_465 : _GEN_1009; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1011 = 9'h1d2 == pht_widx ? pht_466 : _GEN_1010; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1012 = 9'h1d3 == pht_widx ? pht_467 : _GEN_1011; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1013 = 9'h1d4 == pht_widx ? pht_468 : _GEN_1012; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1014 = 9'h1d5 == pht_widx ? pht_469 : _GEN_1013; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1015 = 9'h1d6 == pht_widx ? pht_470 : _GEN_1014; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1016 = 9'h1d7 == pht_widx ? pht_471 : _GEN_1015; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1017 = 9'h1d8 == pht_widx ? pht_472 : _GEN_1016; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1018 = 9'h1d9 == pht_widx ? pht_473 : _GEN_1017; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1019 = 9'h1da == pht_widx ? pht_474 : _GEN_1018; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1020 = 9'h1db == pht_widx ? pht_475 : _GEN_1019; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1021 = 9'h1dc == pht_widx ? pht_476 : _GEN_1020; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1022 = 9'h1dd == pht_widx ? pht_477 : _GEN_1021; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1023 = 9'h1de == pht_widx ? pht_478 : _GEN_1022; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1024 = 9'h1df == pht_widx ? pht_479 : _GEN_1023; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1025 = 9'h1e0 == pht_widx ? pht_480 : _GEN_1024; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1026 = 9'h1e1 == pht_widx ? pht_481 : _GEN_1025; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1027 = 9'h1e2 == pht_widx ? pht_482 : _GEN_1026; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1028 = 9'h1e3 == pht_widx ? pht_483 : _GEN_1027; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1029 = 9'h1e4 == pht_widx ? pht_484 : _GEN_1028; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1030 = 9'h1e5 == pht_widx ? pht_485 : _GEN_1029; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1031 = 9'h1e6 == pht_widx ? pht_486 : _GEN_1030; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1032 = 9'h1e7 == pht_widx ? pht_487 : _GEN_1031; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1033 = 9'h1e8 == pht_widx ? pht_488 : _GEN_1032; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1034 = 9'h1e9 == pht_widx ? pht_489 : _GEN_1033; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1035 = 9'h1ea == pht_widx ? pht_490 : _GEN_1034; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1036 = 9'h1eb == pht_widx ? pht_491 : _GEN_1035; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1037 = 9'h1ec == pht_widx ? pht_492 : _GEN_1036; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1038 = 9'h1ed == pht_widx ? pht_493 : _GEN_1037; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1039 = 9'h1ee == pht_widx ? pht_494 : _GEN_1038; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1040 = 9'h1ef == pht_widx ? pht_495 : _GEN_1039; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1041 = 9'h1f0 == pht_widx ? pht_496 : _GEN_1040; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1042 = 9'h1f1 == pht_widx ? pht_497 : _GEN_1041; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1043 = 9'h1f2 == pht_widx ? pht_498 : _GEN_1042; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1044 = 9'h1f3 == pht_widx ? pht_499 : _GEN_1043; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1045 = 9'h1f4 == pht_widx ? pht_500 : _GEN_1044; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1046 = 9'h1f5 == pht_widx ? pht_501 : _GEN_1045; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1047 = 9'h1f6 == pht_widx ? pht_502 : _GEN_1046; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1048 = 9'h1f7 == pht_widx ? pht_503 : _GEN_1047; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1049 = 9'h1f8 == pht_widx ? pht_504 : _GEN_1048; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1050 = 9'h1f9 == pht_widx ? pht_505 : _GEN_1049; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1051 = 9'h1fa == pht_widx ? pht_506 : _GEN_1050; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1052 = 9'h1fb == pht_widx ? pht_507 : _GEN_1051; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1053 = 9'h1fc == pht_widx ? pht_508 : _GEN_1052; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1054 = 9'h1fd == pht_widx ? pht_509 : _GEN_1053; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1055 = 9'h1fe == pht_widx ? pht_510 : _GEN_1054; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1056 = 9'h1ff == pht_widx ? pht_511 : _GEN_1055; // @[Mux.scala 81:{61,61}]
  wire [1:0] _pht_T_5 = 2'h1 == _GEN_1056 ? _pht_T_1 : {{1'd0}, io_jmp_packet_bp_taken}; // @[Mux.scala 81:58]
  wire [1:0] _pht_T_7 = 2'h2 == _GEN_1056 ? _pht_T_2 : _pht_T_5; // @[Mux.scala 81:58]
  wire [3:0] _GEN_2085 = btb_1_valid & btb_1_tag == io_jmp_packet_bp_pc[38:2] ? 4'h1 : 4'h0; // @[BPU.scala 71:81 73:20]
  wire [3:0] _GEN_2087 = btb_2_valid & btb_2_tag == io_jmp_packet_bp_pc[38:2] ? 4'h2 : _GEN_2085; // @[BPU.scala 71:81 73:20]
  wire [3:0] _GEN_2089 = btb_3_valid & btb_3_tag == io_jmp_packet_bp_pc[38:2] ? 4'h3 : _GEN_2087; // @[BPU.scala 71:81 73:20]
  wire [3:0] _GEN_2091 = btb_4_valid & btb_4_tag == io_jmp_packet_bp_pc[38:2] ? 4'h4 : _GEN_2089; // @[BPU.scala 71:81 73:20]
  wire [3:0] _GEN_2093 = btb_5_valid & btb_5_tag == io_jmp_packet_bp_pc[38:2] ? 4'h5 : _GEN_2091; // @[BPU.scala 71:81 73:20]
  wire [3:0] _GEN_2095 = btb_6_valid & btb_6_tag == io_jmp_packet_bp_pc[38:2] ? 4'h6 : _GEN_2093; // @[BPU.scala 71:81 73:20]
  wire [3:0] _GEN_2097 = btb_7_valid & btb_7_tag == io_jmp_packet_bp_pc[38:2] ? 4'h7 : _GEN_2095; // @[BPU.scala 71:81 73:20]
  wire [3:0] _GEN_2099 = btb_8_valid & btb_8_tag == io_jmp_packet_bp_pc[38:2] ? 4'h8 : _GEN_2097; // @[BPU.scala 71:81 73:20]
  wire  _GEN_2100 = btb_9_valid & btb_9_tag == io_jmp_packet_bp_pc[38:2] | (btb_8_valid & btb_8_tag ==
    io_jmp_packet_bp_pc[38:2] | (btb_7_valid & btb_7_tag == io_jmp_packet_bp_pc[38:2] | (btb_6_valid & btb_6_tag ==
    io_jmp_packet_bp_pc[38:2] | (btb_5_valid & btb_5_tag == io_jmp_packet_bp_pc[38:2] | (btb_4_valid & btb_4_tag ==
    io_jmp_packet_bp_pc[38:2] | (btb_3_valid & btb_3_tag == io_jmp_packet_bp_pc[38:2] | (btb_2_valid & btb_2_tag ==
    io_jmp_packet_bp_pc[38:2] | (btb_1_valid & btb_1_tag == io_jmp_packet_bp_pc[38:2] | btb_0_valid & btb_0_tag ==
    io_jmp_packet_bp_pc[38:2])))))))); // @[BPU.scala 71:81 72:20]
  wire [3:0] _GEN_2101 = btb_9_valid & btb_9_tag == io_jmp_packet_bp_pc[38:2] ? 4'h9 : _GEN_2099; // @[BPU.scala 71:81 73:20]
  wire [3:0] _GEN_2103 = btb_10_valid & btb_10_tag == io_jmp_packet_bp_pc[38:2] ? 4'ha : _GEN_2101; // @[BPU.scala 71:81 73:20]
  wire [3:0] _GEN_2105 = btb_11_valid & btb_11_tag == io_jmp_packet_bp_pc[38:2] ? 4'hb : _GEN_2103; // @[BPU.scala 71:81 73:20]
  wire [3:0] _GEN_2107 = btb_12_valid & btb_12_tag == io_jmp_packet_bp_pc[38:2] ? 4'hc : _GEN_2105; // @[BPU.scala 71:81 73:20]
  wire [3:0] _GEN_2109 = btb_13_valid & btb_13_tag == io_jmp_packet_bp_pc[38:2] ? 4'hd : _GEN_2107; // @[BPU.scala 71:81 73:20]
  wire [3:0] _GEN_2111 = btb_14_valid & btb_14_tag == io_jmp_packet_bp_pc[38:2] ? 4'he : _GEN_2109; // @[BPU.scala 71:81 73:20]
  wire  btb_whit = btb_15_valid & btb_15_tag == io_jmp_packet_bp_pc[38:2] | (btb_14_valid & btb_14_tag ==
    io_jmp_packet_bp_pc[38:2] | (btb_13_valid & btb_13_tag == io_jmp_packet_bp_pc[38:2] | (btb_12_valid & btb_12_tag ==
    io_jmp_packet_bp_pc[38:2] | (btb_11_valid & btb_11_tag == io_jmp_packet_bp_pc[38:2] | (btb_10_valid & btb_10_tag ==
    io_jmp_packet_bp_pc[38:2] | _GEN_2100))))); // @[BPU.scala 71:81 72:20]
  wire [3:0] btb_whit_way = btb_15_valid & btb_15_tag == io_jmp_packet_bp_pc[38:2] ? 4'hf : _GEN_2111; // @[BPU.scala 71:81 73:20]
  wire [3:0] _btb_replace_idx_T = {btb_replace_idx_prng_io_out_3,btb_replace_idx_prng_io_out_2,
    btb_replace_idx_prng_io_out_1,btb_replace_idx_prng_io_out_0}; // @[PRNG.scala 95:17]
  wire [3:0] btb_replace_idx = btb_whit ? btb_whit_way : _btb_replace_idx_T; // @[BPU.scala 77:25]
  wire  _GEN_2114 = 4'h0 == btb_replace_idx | btb_0_valid; // @[BPU.scala 28:20 79:{33,33}]
  wire  _GEN_2115 = 4'h1 == btb_replace_idx | btb_1_valid; // @[BPU.scala 28:20 79:{33,33}]
  wire  _GEN_2116 = 4'h2 == btb_replace_idx | btb_2_valid; // @[BPU.scala 28:20 79:{33,33}]
  wire  _GEN_2117 = 4'h3 == btb_replace_idx | btb_3_valid; // @[BPU.scala 28:20 79:{33,33}]
  wire  _GEN_2118 = 4'h4 == btb_replace_idx | btb_4_valid; // @[BPU.scala 28:20 79:{33,33}]
  wire  _GEN_2119 = 4'h5 == btb_replace_idx | btb_5_valid; // @[BPU.scala 28:20 79:{33,33}]
  wire  _GEN_2120 = 4'h6 == btb_replace_idx | btb_6_valid; // @[BPU.scala 28:20 79:{33,33}]
  wire  _GEN_2121 = 4'h7 == btb_replace_idx | btb_7_valid; // @[BPU.scala 28:20 79:{33,33}]
  wire  _GEN_2122 = 4'h8 == btb_replace_idx | btb_8_valid; // @[BPU.scala 28:20 79:{33,33}]
  wire  _GEN_2123 = 4'h9 == btb_replace_idx | btb_9_valid; // @[BPU.scala 28:20 79:{33,33}]
  wire  _GEN_2124 = 4'ha == btb_replace_idx | btb_10_valid; // @[BPU.scala 28:20 79:{33,33}]
  wire  _GEN_2125 = 4'hb == btb_replace_idx | btb_11_valid; // @[BPU.scala 28:20 79:{33,33}]
  wire  _GEN_2126 = 4'hc == btb_replace_idx | btb_12_valid; // @[BPU.scala 28:20 79:{33,33}]
  wire  _GEN_2127 = 4'hd == btb_replace_idx | btb_13_valid; // @[BPU.scala 28:20 79:{33,33}]
  wire  _GEN_2128 = 4'he == btb_replace_idx | btb_14_valid; // @[BPU.scala 28:20 79:{33,33}]
  wire  _GEN_2129 = 4'hf == btb_replace_idx | btb_15_valid; // @[BPU.scala 28:20 79:{33,33}]
  MaxPeriodFibonacciLFSR btb_replace_idx_prng ( // @[PRNG.scala 91:22]
    .clock(btb_replace_idx_prng_clock),
    .reset(btb_replace_idx_prng_reset),
    .io_out_0(btb_replace_idx_prng_io_out_0),
    .io_out_1(btb_replace_idx_prng_io_out_1),
    .io_out_2(btb_replace_idx_prng_io_out_2),
    .io_out_3(btb_replace_idx_prng_io_out_3)
  );
  assign io_out = pht_taken & btb_rhit ? _io_out_T_6 : _io_out_T_1; // @[BPU.scala 46:10 47:31 48:12]
  assign btb_replace_idx_prng_clock = clock;
  assign btb_replace_idx_prng_reset = reset;
  always @(posedge clock) begin
    if (reset) begin // @[BPU.scala 26:20]
      ghr <= 9'h0; // @[BPU.scala 26:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      ghr <= {{1'd0}, _ghr_T_1}; // @[BPU.scala 54:9]
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_0 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h0 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_0 <= _pht_T_3;
        end else begin
          pht_0 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_1 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_1 <= _pht_T_3;
        end else begin
          pht_1 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_2 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h2 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_2 <= _pht_T_3;
        end else begin
          pht_2 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_3 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h3 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_3 <= _pht_T_3;
        end else begin
          pht_3 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_4 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h4 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_4 <= _pht_T_3;
        end else begin
          pht_4 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_5 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h5 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_5 <= _pht_T_3;
        end else begin
          pht_5 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_6 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h6 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_6 <= _pht_T_3;
        end else begin
          pht_6 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_7 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h7 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_7 <= _pht_T_3;
        end else begin
          pht_7 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_8 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h8 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_8 <= _pht_T_3;
        end else begin
          pht_8 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_9 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h9 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_9 <= _pht_T_3;
        end else begin
          pht_9 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_10 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'ha == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_10 <= _pht_T_3;
        end else begin
          pht_10 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_11 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hb == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_11 <= _pht_T_3;
        end else begin
          pht_11 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_12 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hc == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_12 <= _pht_T_3;
        end else begin
          pht_12 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_13 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hd == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_13 <= _pht_T_3;
        end else begin
          pht_13 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_14 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'he == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_14 <= _pht_T_3;
        end else begin
          pht_14 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_15 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hf == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_15 <= _pht_T_3;
        end else begin
          pht_15 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_16 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h10 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_16 <= _pht_T_3;
        end else begin
          pht_16 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_17 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h11 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_17 <= _pht_T_3;
        end else begin
          pht_17 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_18 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h12 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_18 <= _pht_T_3;
        end else begin
          pht_18 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_19 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h13 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_19 <= _pht_T_3;
        end else begin
          pht_19 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_20 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h14 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_20 <= _pht_T_3;
        end else begin
          pht_20 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_21 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h15 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_21 <= _pht_T_3;
        end else begin
          pht_21 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_22 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h16 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_22 <= _pht_T_3;
        end else begin
          pht_22 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_23 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h17 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_23 <= _pht_T_3;
        end else begin
          pht_23 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_24 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h18 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_24 <= _pht_T_3;
        end else begin
          pht_24 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_25 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h19 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_25 <= _pht_T_3;
        end else begin
          pht_25 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_26 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1a == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_26 <= _pht_T_3;
        end else begin
          pht_26 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_27 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1b == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_27 <= _pht_T_3;
        end else begin
          pht_27 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_28 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1c == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_28 <= _pht_T_3;
        end else begin
          pht_28 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_29 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1d == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_29 <= _pht_T_3;
        end else begin
          pht_29 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_30 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1e == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_30 <= _pht_T_3;
        end else begin
          pht_30 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_31 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1f == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_31 <= _pht_T_3;
        end else begin
          pht_31 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_32 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h20 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_32 <= _pht_T_3;
        end else begin
          pht_32 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_33 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h21 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_33 <= _pht_T_3;
        end else begin
          pht_33 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_34 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h22 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_34 <= _pht_T_3;
        end else begin
          pht_34 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_35 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h23 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_35 <= _pht_T_3;
        end else begin
          pht_35 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_36 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h24 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_36 <= _pht_T_3;
        end else begin
          pht_36 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_37 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h25 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_37 <= _pht_T_3;
        end else begin
          pht_37 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_38 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h26 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_38 <= _pht_T_3;
        end else begin
          pht_38 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_39 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h27 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_39 <= _pht_T_3;
        end else begin
          pht_39 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_40 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h28 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_40 <= _pht_T_3;
        end else begin
          pht_40 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_41 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h29 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_41 <= _pht_T_3;
        end else begin
          pht_41 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_42 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h2a == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_42 <= _pht_T_3;
        end else begin
          pht_42 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_43 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h2b == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_43 <= _pht_T_3;
        end else begin
          pht_43 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_44 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h2c == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_44 <= _pht_T_3;
        end else begin
          pht_44 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_45 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h2d == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_45 <= _pht_T_3;
        end else begin
          pht_45 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_46 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h2e == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_46 <= _pht_T_3;
        end else begin
          pht_46 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_47 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h2f == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_47 <= _pht_T_3;
        end else begin
          pht_47 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_48 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h30 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_48 <= _pht_T_3;
        end else begin
          pht_48 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_49 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h31 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_49 <= _pht_T_3;
        end else begin
          pht_49 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_50 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h32 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_50 <= _pht_T_3;
        end else begin
          pht_50 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_51 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h33 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_51 <= _pht_T_3;
        end else begin
          pht_51 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_52 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h34 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_52 <= _pht_T_3;
        end else begin
          pht_52 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_53 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h35 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_53 <= _pht_T_3;
        end else begin
          pht_53 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_54 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h36 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_54 <= _pht_T_3;
        end else begin
          pht_54 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_55 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h37 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_55 <= _pht_T_3;
        end else begin
          pht_55 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_56 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h38 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_56 <= _pht_T_3;
        end else begin
          pht_56 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_57 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h39 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_57 <= _pht_T_3;
        end else begin
          pht_57 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_58 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h3a == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_58 <= _pht_T_3;
        end else begin
          pht_58 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_59 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h3b == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_59 <= _pht_T_3;
        end else begin
          pht_59 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_60 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h3c == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_60 <= _pht_T_3;
        end else begin
          pht_60 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_61 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h3d == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_61 <= _pht_T_3;
        end else begin
          pht_61 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_62 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h3e == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_62 <= _pht_T_3;
        end else begin
          pht_62 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_63 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h3f == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_63 <= _pht_T_3;
        end else begin
          pht_63 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_64 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h40 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_64 <= _pht_T_3;
        end else begin
          pht_64 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_65 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h41 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_65 <= _pht_T_3;
        end else begin
          pht_65 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_66 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h42 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_66 <= _pht_T_3;
        end else begin
          pht_66 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_67 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h43 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_67 <= _pht_T_3;
        end else begin
          pht_67 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_68 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h44 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_68 <= _pht_T_3;
        end else begin
          pht_68 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_69 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h45 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_69 <= _pht_T_3;
        end else begin
          pht_69 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_70 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h46 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_70 <= _pht_T_3;
        end else begin
          pht_70 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_71 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h47 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_71 <= _pht_T_3;
        end else begin
          pht_71 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_72 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h48 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_72 <= _pht_T_3;
        end else begin
          pht_72 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_73 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h49 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_73 <= _pht_T_3;
        end else begin
          pht_73 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_74 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h4a == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_74 <= _pht_T_3;
        end else begin
          pht_74 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_75 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h4b == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_75 <= _pht_T_3;
        end else begin
          pht_75 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_76 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h4c == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_76 <= _pht_T_3;
        end else begin
          pht_76 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_77 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h4d == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_77 <= _pht_T_3;
        end else begin
          pht_77 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_78 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h4e == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_78 <= _pht_T_3;
        end else begin
          pht_78 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_79 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h4f == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_79 <= _pht_T_3;
        end else begin
          pht_79 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_80 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h50 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_80 <= _pht_T_3;
        end else begin
          pht_80 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_81 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h51 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_81 <= _pht_T_3;
        end else begin
          pht_81 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_82 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h52 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_82 <= _pht_T_3;
        end else begin
          pht_82 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_83 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h53 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_83 <= _pht_T_3;
        end else begin
          pht_83 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_84 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h54 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_84 <= _pht_T_3;
        end else begin
          pht_84 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_85 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h55 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_85 <= _pht_T_3;
        end else begin
          pht_85 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_86 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h56 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_86 <= _pht_T_3;
        end else begin
          pht_86 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_87 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h57 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_87 <= _pht_T_3;
        end else begin
          pht_87 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_88 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h58 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_88 <= _pht_T_3;
        end else begin
          pht_88 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_89 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h59 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_89 <= _pht_T_3;
        end else begin
          pht_89 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_90 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h5a == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_90 <= _pht_T_3;
        end else begin
          pht_90 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_91 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h5b == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_91 <= _pht_T_3;
        end else begin
          pht_91 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_92 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h5c == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_92 <= _pht_T_3;
        end else begin
          pht_92 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_93 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h5d == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_93 <= _pht_T_3;
        end else begin
          pht_93 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_94 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h5e == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_94 <= _pht_T_3;
        end else begin
          pht_94 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_95 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h5f == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_95 <= _pht_T_3;
        end else begin
          pht_95 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_96 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h60 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_96 <= _pht_T_3;
        end else begin
          pht_96 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_97 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h61 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_97 <= _pht_T_3;
        end else begin
          pht_97 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_98 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h62 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_98 <= _pht_T_3;
        end else begin
          pht_98 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_99 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h63 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_99 <= _pht_T_3;
        end else begin
          pht_99 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_100 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h64 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_100 <= _pht_T_3;
        end else begin
          pht_100 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_101 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h65 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_101 <= _pht_T_3;
        end else begin
          pht_101 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_102 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h66 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_102 <= _pht_T_3;
        end else begin
          pht_102 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_103 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h67 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_103 <= _pht_T_3;
        end else begin
          pht_103 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_104 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h68 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_104 <= _pht_T_3;
        end else begin
          pht_104 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_105 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h69 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_105 <= _pht_T_3;
        end else begin
          pht_105 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_106 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h6a == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_106 <= _pht_T_3;
        end else begin
          pht_106 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_107 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h6b == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_107 <= _pht_T_3;
        end else begin
          pht_107 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_108 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h6c == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_108 <= _pht_T_3;
        end else begin
          pht_108 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_109 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h6d == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_109 <= _pht_T_3;
        end else begin
          pht_109 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_110 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h6e == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_110 <= _pht_T_3;
        end else begin
          pht_110 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_111 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h6f == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_111 <= _pht_T_3;
        end else begin
          pht_111 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_112 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h70 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_112 <= _pht_T_3;
        end else begin
          pht_112 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_113 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h71 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_113 <= _pht_T_3;
        end else begin
          pht_113 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_114 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h72 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_114 <= _pht_T_3;
        end else begin
          pht_114 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_115 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h73 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_115 <= _pht_T_3;
        end else begin
          pht_115 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_116 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h74 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_116 <= _pht_T_3;
        end else begin
          pht_116 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_117 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h75 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_117 <= _pht_T_3;
        end else begin
          pht_117 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_118 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h76 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_118 <= _pht_T_3;
        end else begin
          pht_118 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_119 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h77 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_119 <= _pht_T_3;
        end else begin
          pht_119 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_120 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h78 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_120 <= _pht_T_3;
        end else begin
          pht_120 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_121 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h79 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_121 <= _pht_T_3;
        end else begin
          pht_121 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_122 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h7a == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_122 <= _pht_T_3;
        end else begin
          pht_122 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_123 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h7b == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_123 <= _pht_T_3;
        end else begin
          pht_123 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_124 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h7c == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_124 <= _pht_T_3;
        end else begin
          pht_124 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_125 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h7d == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_125 <= _pht_T_3;
        end else begin
          pht_125 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_126 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h7e == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_126 <= _pht_T_3;
        end else begin
          pht_126 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_127 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h7f == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_127 <= _pht_T_3;
        end else begin
          pht_127 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_128 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h80 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_128 <= _pht_T_3;
        end else begin
          pht_128 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_129 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h81 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_129 <= _pht_T_3;
        end else begin
          pht_129 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_130 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h82 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_130 <= _pht_T_3;
        end else begin
          pht_130 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_131 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h83 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_131 <= _pht_T_3;
        end else begin
          pht_131 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_132 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h84 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_132 <= _pht_T_3;
        end else begin
          pht_132 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_133 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h85 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_133 <= _pht_T_3;
        end else begin
          pht_133 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_134 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h86 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_134 <= _pht_T_3;
        end else begin
          pht_134 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_135 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h87 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_135 <= _pht_T_3;
        end else begin
          pht_135 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_136 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h88 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_136 <= _pht_T_3;
        end else begin
          pht_136 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_137 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h89 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_137 <= _pht_T_3;
        end else begin
          pht_137 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_138 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h8a == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_138 <= _pht_T_3;
        end else begin
          pht_138 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_139 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h8b == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_139 <= _pht_T_3;
        end else begin
          pht_139 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_140 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h8c == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_140 <= _pht_T_3;
        end else begin
          pht_140 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_141 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h8d == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_141 <= _pht_T_3;
        end else begin
          pht_141 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_142 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h8e == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_142 <= _pht_T_3;
        end else begin
          pht_142 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_143 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h8f == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_143 <= _pht_T_3;
        end else begin
          pht_143 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_144 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h90 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_144 <= _pht_T_3;
        end else begin
          pht_144 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_145 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h91 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_145 <= _pht_T_3;
        end else begin
          pht_145 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_146 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h92 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_146 <= _pht_T_3;
        end else begin
          pht_146 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_147 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h93 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_147 <= _pht_T_3;
        end else begin
          pht_147 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_148 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h94 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_148 <= _pht_T_3;
        end else begin
          pht_148 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_149 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h95 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_149 <= _pht_T_3;
        end else begin
          pht_149 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_150 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h96 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_150 <= _pht_T_3;
        end else begin
          pht_150 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_151 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h97 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_151 <= _pht_T_3;
        end else begin
          pht_151 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_152 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h98 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_152 <= _pht_T_3;
        end else begin
          pht_152 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_153 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h99 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_153 <= _pht_T_3;
        end else begin
          pht_153 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_154 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h9a == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_154 <= _pht_T_3;
        end else begin
          pht_154 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_155 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h9b == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_155 <= _pht_T_3;
        end else begin
          pht_155 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_156 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h9c == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_156 <= _pht_T_3;
        end else begin
          pht_156 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_157 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h9d == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_157 <= _pht_T_3;
        end else begin
          pht_157 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_158 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h9e == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_158 <= _pht_T_3;
        end else begin
          pht_158 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_159 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h9f == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_159 <= _pht_T_3;
        end else begin
          pht_159 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_160 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'ha0 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_160 <= _pht_T_3;
        end else begin
          pht_160 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_161 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'ha1 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_161 <= _pht_T_3;
        end else begin
          pht_161 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_162 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'ha2 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_162 <= _pht_T_3;
        end else begin
          pht_162 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_163 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'ha3 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_163 <= _pht_T_3;
        end else begin
          pht_163 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_164 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'ha4 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_164 <= _pht_T_3;
        end else begin
          pht_164 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_165 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'ha5 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_165 <= _pht_T_3;
        end else begin
          pht_165 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_166 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'ha6 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_166 <= _pht_T_3;
        end else begin
          pht_166 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_167 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'ha7 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_167 <= _pht_T_3;
        end else begin
          pht_167 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_168 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'ha8 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_168 <= _pht_T_3;
        end else begin
          pht_168 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_169 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'ha9 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_169 <= _pht_T_3;
        end else begin
          pht_169 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_170 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'haa == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_170 <= _pht_T_3;
        end else begin
          pht_170 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_171 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hab == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_171 <= _pht_T_3;
        end else begin
          pht_171 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_172 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hac == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_172 <= _pht_T_3;
        end else begin
          pht_172 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_173 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'had == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_173 <= _pht_T_3;
        end else begin
          pht_173 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_174 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hae == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_174 <= _pht_T_3;
        end else begin
          pht_174 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_175 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'haf == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_175 <= _pht_T_3;
        end else begin
          pht_175 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_176 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hb0 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_176 <= _pht_T_3;
        end else begin
          pht_176 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_177 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hb1 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_177 <= _pht_T_3;
        end else begin
          pht_177 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_178 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hb2 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_178 <= _pht_T_3;
        end else begin
          pht_178 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_179 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hb3 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_179 <= _pht_T_3;
        end else begin
          pht_179 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_180 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hb4 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_180 <= _pht_T_3;
        end else begin
          pht_180 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_181 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hb5 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_181 <= _pht_T_3;
        end else begin
          pht_181 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_182 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hb6 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_182 <= _pht_T_3;
        end else begin
          pht_182 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_183 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hb7 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_183 <= _pht_T_3;
        end else begin
          pht_183 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_184 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hb8 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_184 <= _pht_T_3;
        end else begin
          pht_184 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_185 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hb9 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_185 <= _pht_T_3;
        end else begin
          pht_185 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_186 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hba == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_186 <= _pht_T_3;
        end else begin
          pht_186 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_187 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hbb == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_187 <= _pht_T_3;
        end else begin
          pht_187 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_188 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hbc == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_188 <= _pht_T_3;
        end else begin
          pht_188 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_189 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hbd == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_189 <= _pht_T_3;
        end else begin
          pht_189 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_190 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hbe == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_190 <= _pht_T_3;
        end else begin
          pht_190 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_191 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hbf == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_191 <= _pht_T_3;
        end else begin
          pht_191 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_192 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hc0 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_192 <= _pht_T_3;
        end else begin
          pht_192 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_193 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hc1 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_193 <= _pht_T_3;
        end else begin
          pht_193 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_194 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hc2 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_194 <= _pht_T_3;
        end else begin
          pht_194 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_195 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hc3 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_195 <= _pht_T_3;
        end else begin
          pht_195 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_196 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hc4 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_196 <= _pht_T_3;
        end else begin
          pht_196 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_197 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hc5 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_197 <= _pht_T_3;
        end else begin
          pht_197 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_198 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hc6 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_198 <= _pht_T_3;
        end else begin
          pht_198 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_199 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hc7 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_199 <= _pht_T_3;
        end else begin
          pht_199 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_200 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hc8 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_200 <= _pht_T_3;
        end else begin
          pht_200 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_201 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hc9 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_201 <= _pht_T_3;
        end else begin
          pht_201 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_202 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hca == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_202 <= _pht_T_3;
        end else begin
          pht_202 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_203 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hcb == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_203 <= _pht_T_3;
        end else begin
          pht_203 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_204 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hcc == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_204 <= _pht_T_3;
        end else begin
          pht_204 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_205 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hcd == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_205 <= _pht_T_3;
        end else begin
          pht_205 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_206 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hce == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_206 <= _pht_T_3;
        end else begin
          pht_206 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_207 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hcf == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_207 <= _pht_T_3;
        end else begin
          pht_207 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_208 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hd0 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_208 <= _pht_T_3;
        end else begin
          pht_208 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_209 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hd1 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_209 <= _pht_T_3;
        end else begin
          pht_209 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_210 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hd2 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_210 <= _pht_T_3;
        end else begin
          pht_210 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_211 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hd3 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_211 <= _pht_T_3;
        end else begin
          pht_211 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_212 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hd4 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_212 <= _pht_T_3;
        end else begin
          pht_212 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_213 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hd5 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_213 <= _pht_T_3;
        end else begin
          pht_213 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_214 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hd6 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_214 <= _pht_T_3;
        end else begin
          pht_214 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_215 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hd7 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_215 <= _pht_T_3;
        end else begin
          pht_215 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_216 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hd8 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_216 <= _pht_T_3;
        end else begin
          pht_216 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_217 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hd9 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_217 <= _pht_T_3;
        end else begin
          pht_217 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_218 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hda == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_218 <= _pht_T_3;
        end else begin
          pht_218 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_219 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hdb == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_219 <= _pht_T_3;
        end else begin
          pht_219 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_220 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hdc == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_220 <= _pht_T_3;
        end else begin
          pht_220 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_221 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hdd == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_221 <= _pht_T_3;
        end else begin
          pht_221 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_222 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hde == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_222 <= _pht_T_3;
        end else begin
          pht_222 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_223 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hdf == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_223 <= _pht_T_3;
        end else begin
          pht_223 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_224 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'he0 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_224 <= _pht_T_3;
        end else begin
          pht_224 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_225 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'he1 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_225 <= _pht_T_3;
        end else begin
          pht_225 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_226 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'he2 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_226 <= _pht_T_3;
        end else begin
          pht_226 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_227 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'he3 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_227 <= _pht_T_3;
        end else begin
          pht_227 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_228 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'he4 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_228 <= _pht_T_3;
        end else begin
          pht_228 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_229 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'he5 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_229 <= _pht_T_3;
        end else begin
          pht_229 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_230 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'he6 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_230 <= _pht_T_3;
        end else begin
          pht_230 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_231 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'he7 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_231 <= _pht_T_3;
        end else begin
          pht_231 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_232 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'he8 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_232 <= _pht_T_3;
        end else begin
          pht_232 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_233 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'he9 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_233 <= _pht_T_3;
        end else begin
          pht_233 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_234 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hea == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_234 <= _pht_T_3;
        end else begin
          pht_234 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_235 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'heb == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_235 <= _pht_T_3;
        end else begin
          pht_235 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_236 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hec == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_236 <= _pht_T_3;
        end else begin
          pht_236 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_237 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hed == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_237 <= _pht_T_3;
        end else begin
          pht_237 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_238 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hee == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_238 <= _pht_T_3;
        end else begin
          pht_238 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_239 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hef == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_239 <= _pht_T_3;
        end else begin
          pht_239 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_240 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hf0 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_240 <= _pht_T_3;
        end else begin
          pht_240 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_241 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hf1 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_241 <= _pht_T_3;
        end else begin
          pht_241 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_242 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hf2 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_242 <= _pht_T_3;
        end else begin
          pht_242 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_243 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hf3 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_243 <= _pht_T_3;
        end else begin
          pht_243 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_244 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hf4 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_244 <= _pht_T_3;
        end else begin
          pht_244 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_245 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hf5 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_245 <= _pht_T_3;
        end else begin
          pht_245 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_246 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hf6 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_246 <= _pht_T_3;
        end else begin
          pht_246 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_247 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hf7 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_247 <= _pht_T_3;
        end else begin
          pht_247 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_248 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hf8 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_248 <= _pht_T_3;
        end else begin
          pht_248 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_249 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hf9 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_249 <= _pht_T_3;
        end else begin
          pht_249 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_250 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hfa == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_250 <= _pht_T_3;
        end else begin
          pht_250 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_251 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hfb == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_251 <= _pht_T_3;
        end else begin
          pht_251 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_252 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hfc == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_252 <= _pht_T_3;
        end else begin
          pht_252 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_253 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hfd == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_253 <= _pht_T_3;
        end else begin
          pht_253 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_254 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hfe == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_254 <= _pht_T_3;
        end else begin
          pht_254 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_255 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hff == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_255 <= _pht_T_3;
        end else begin
          pht_255 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_256 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h100 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_256 <= _pht_T_3;
        end else begin
          pht_256 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_257 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h101 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_257 <= _pht_T_3;
        end else begin
          pht_257 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_258 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h102 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_258 <= _pht_T_3;
        end else begin
          pht_258 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_259 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h103 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_259 <= _pht_T_3;
        end else begin
          pht_259 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_260 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h104 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_260 <= _pht_T_3;
        end else begin
          pht_260 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_261 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h105 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_261 <= _pht_T_3;
        end else begin
          pht_261 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_262 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h106 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_262 <= _pht_T_3;
        end else begin
          pht_262 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_263 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h107 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_263 <= _pht_T_3;
        end else begin
          pht_263 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_264 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h108 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_264 <= _pht_T_3;
        end else begin
          pht_264 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_265 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h109 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_265 <= _pht_T_3;
        end else begin
          pht_265 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_266 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h10a == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_266 <= _pht_T_3;
        end else begin
          pht_266 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_267 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h10b == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_267 <= _pht_T_3;
        end else begin
          pht_267 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_268 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h10c == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_268 <= _pht_T_3;
        end else begin
          pht_268 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_269 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h10d == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_269 <= _pht_T_3;
        end else begin
          pht_269 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_270 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h10e == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_270 <= _pht_T_3;
        end else begin
          pht_270 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_271 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h10f == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_271 <= _pht_T_3;
        end else begin
          pht_271 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_272 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h110 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_272 <= _pht_T_3;
        end else begin
          pht_272 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_273 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h111 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_273 <= _pht_T_3;
        end else begin
          pht_273 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_274 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h112 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_274 <= _pht_T_3;
        end else begin
          pht_274 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_275 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h113 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_275 <= _pht_T_3;
        end else begin
          pht_275 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_276 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h114 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_276 <= _pht_T_3;
        end else begin
          pht_276 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_277 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h115 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_277 <= _pht_T_3;
        end else begin
          pht_277 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_278 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h116 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_278 <= _pht_T_3;
        end else begin
          pht_278 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_279 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h117 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_279 <= _pht_T_3;
        end else begin
          pht_279 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_280 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h118 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_280 <= _pht_T_3;
        end else begin
          pht_280 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_281 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h119 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_281 <= _pht_T_3;
        end else begin
          pht_281 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_282 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h11a == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_282 <= _pht_T_3;
        end else begin
          pht_282 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_283 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h11b == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_283 <= _pht_T_3;
        end else begin
          pht_283 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_284 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h11c == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_284 <= _pht_T_3;
        end else begin
          pht_284 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_285 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h11d == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_285 <= _pht_T_3;
        end else begin
          pht_285 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_286 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h11e == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_286 <= _pht_T_3;
        end else begin
          pht_286 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_287 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h11f == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_287 <= _pht_T_3;
        end else begin
          pht_287 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_288 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h120 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_288 <= _pht_T_3;
        end else begin
          pht_288 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_289 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h121 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_289 <= _pht_T_3;
        end else begin
          pht_289 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_290 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h122 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_290 <= _pht_T_3;
        end else begin
          pht_290 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_291 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h123 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_291 <= _pht_T_3;
        end else begin
          pht_291 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_292 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h124 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_292 <= _pht_T_3;
        end else begin
          pht_292 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_293 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h125 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_293 <= _pht_T_3;
        end else begin
          pht_293 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_294 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h126 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_294 <= _pht_T_3;
        end else begin
          pht_294 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_295 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h127 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_295 <= _pht_T_3;
        end else begin
          pht_295 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_296 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h128 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_296 <= _pht_T_3;
        end else begin
          pht_296 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_297 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h129 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_297 <= _pht_T_3;
        end else begin
          pht_297 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_298 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h12a == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_298 <= _pht_T_3;
        end else begin
          pht_298 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_299 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h12b == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_299 <= _pht_T_3;
        end else begin
          pht_299 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_300 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h12c == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_300 <= _pht_T_3;
        end else begin
          pht_300 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_301 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h12d == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_301 <= _pht_T_3;
        end else begin
          pht_301 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_302 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h12e == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_302 <= _pht_T_3;
        end else begin
          pht_302 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_303 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h12f == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_303 <= _pht_T_3;
        end else begin
          pht_303 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_304 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h130 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_304 <= _pht_T_3;
        end else begin
          pht_304 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_305 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h131 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_305 <= _pht_T_3;
        end else begin
          pht_305 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_306 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h132 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_306 <= _pht_T_3;
        end else begin
          pht_306 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_307 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h133 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_307 <= _pht_T_3;
        end else begin
          pht_307 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_308 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h134 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_308 <= _pht_T_3;
        end else begin
          pht_308 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_309 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h135 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_309 <= _pht_T_3;
        end else begin
          pht_309 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_310 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h136 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_310 <= _pht_T_3;
        end else begin
          pht_310 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_311 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h137 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_311 <= _pht_T_3;
        end else begin
          pht_311 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_312 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h138 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_312 <= _pht_T_3;
        end else begin
          pht_312 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_313 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h139 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_313 <= _pht_T_3;
        end else begin
          pht_313 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_314 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h13a == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_314 <= _pht_T_3;
        end else begin
          pht_314 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_315 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h13b == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_315 <= _pht_T_3;
        end else begin
          pht_315 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_316 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h13c == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_316 <= _pht_T_3;
        end else begin
          pht_316 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_317 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h13d == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_317 <= _pht_T_3;
        end else begin
          pht_317 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_318 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h13e == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_318 <= _pht_T_3;
        end else begin
          pht_318 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_319 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h13f == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_319 <= _pht_T_3;
        end else begin
          pht_319 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_320 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h140 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_320 <= _pht_T_3;
        end else begin
          pht_320 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_321 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h141 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_321 <= _pht_T_3;
        end else begin
          pht_321 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_322 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h142 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_322 <= _pht_T_3;
        end else begin
          pht_322 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_323 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h143 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_323 <= _pht_T_3;
        end else begin
          pht_323 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_324 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h144 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_324 <= _pht_T_3;
        end else begin
          pht_324 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_325 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h145 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_325 <= _pht_T_3;
        end else begin
          pht_325 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_326 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h146 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_326 <= _pht_T_3;
        end else begin
          pht_326 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_327 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h147 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_327 <= _pht_T_3;
        end else begin
          pht_327 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_328 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h148 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_328 <= _pht_T_3;
        end else begin
          pht_328 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_329 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h149 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_329 <= _pht_T_3;
        end else begin
          pht_329 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_330 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h14a == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_330 <= _pht_T_3;
        end else begin
          pht_330 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_331 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h14b == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_331 <= _pht_T_3;
        end else begin
          pht_331 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_332 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h14c == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_332 <= _pht_T_3;
        end else begin
          pht_332 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_333 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h14d == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_333 <= _pht_T_3;
        end else begin
          pht_333 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_334 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h14e == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_334 <= _pht_T_3;
        end else begin
          pht_334 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_335 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h14f == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_335 <= _pht_T_3;
        end else begin
          pht_335 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_336 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h150 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_336 <= _pht_T_3;
        end else begin
          pht_336 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_337 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h151 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_337 <= _pht_T_3;
        end else begin
          pht_337 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_338 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h152 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_338 <= _pht_T_3;
        end else begin
          pht_338 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_339 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h153 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_339 <= _pht_T_3;
        end else begin
          pht_339 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_340 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h154 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_340 <= _pht_T_3;
        end else begin
          pht_340 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_341 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h155 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_341 <= _pht_T_3;
        end else begin
          pht_341 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_342 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h156 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_342 <= _pht_T_3;
        end else begin
          pht_342 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_343 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h157 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_343 <= _pht_T_3;
        end else begin
          pht_343 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_344 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h158 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_344 <= _pht_T_3;
        end else begin
          pht_344 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_345 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h159 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_345 <= _pht_T_3;
        end else begin
          pht_345 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_346 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h15a == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_346 <= _pht_T_3;
        end else begin
          pht_346 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_347 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h15b == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_347 <= _pht_T_3;
        end else begin
          pht_347 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_348 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h15c == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_348 <= _pht_T_3;
        end else begin
          pht_348 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_349 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h15d == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_349 <= _pht_T_3;
        end else begin
          pht_349 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_350 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h15e == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_350 <= _pht_T_3;
        end else begin
          pht_350 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_351 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h15f == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_351 <= _pht_T_3;
        end else begin
          pht_351 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_352 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h160 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_352 <= _pht_T_3;
        end else begin
          pht_352 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_353 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h161 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_353 <= _pht_T_3;
        end else begin
          pht_353 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_354 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h162 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_354 <= _pht_T_3;
        end else begin
          pht_354 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_355 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h163 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_355 <= _pht_T_3;
        end else begin
          pht_355 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_356 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h164 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_356 <= _pht_T_3;
        end else begin
          pht_356 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_357 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h165 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_357 <= _pht_T_3;
        end else begin
          pht_357 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_358 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h166 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_358 <= _pht_T_3;
        end else begin
          pht_358 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_359 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h167 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_359 <= _pht_T_3;
        end else begin
          pht_359 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_360 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h168 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_360 <= _pht_T_3;
        end else begin
          pht_360 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_361 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h169 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_361 <= _pht_T_3;
        end else begin
          pht_361 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_362 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h16a == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_362 <= _pht_T_3;
        end else begin
          pht_362 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_363 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h16b == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_363 <= _pht_T_3;
        end else begin
          pht_363 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_364 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h16c == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_364 <= _pht_T_3;
        end else begin
          pht_364 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_365 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h16d == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_365 <= _pht_T_3;
        end else begin
          pht_365 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_366 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h16e == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_366 <= _pht_T_3;
        end else begin
          pht_366 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_367 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h16f == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_367 <= _pht_T_3;
        end else begin
          pht_367 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_368 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h170 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_368 <= _pht_T_3;
        end else begin
          pht_368 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_369 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h171 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_369 <= _pht_T_3;
        end else begin
          pht_369 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_370 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h172 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_370 <= _pht_T_3;
        end else begin
          pht_370 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_371 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h173 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_371 <= _pht_T_3;
        end else begin
          pht_371 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_372 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h174 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_372 <= _pht_T_3;
        end else begin
          pht_372 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_373 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h175 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_373 <= _pht_T_3;
        end else begin
          pht_373 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_374 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h176 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_374 <= _pht_T_3;
        end else begin
          pht_374 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_375 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h177 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_375 <= _pht_T_3;
        end else begin
          pht_375 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_376 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h178 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_376 <= _pht_T_3;
        end else begin
          pht_376 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_377 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h179 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_377 <= _pht_T_3;
        end else begin
          pht_377 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_378 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h17a == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_378 <= _pht_T_3;
        end else begin
          pht_378 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_379 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h17b == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_379 <= _pht_T_3;
        end else begin
          pht_379 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_380 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h17c == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_380 <= _pht_T_3;
        end else begin
          pht_380 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_381 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h17d == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_381 <= _pht_T_3;
        end else begin
          pht_381 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_382 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h17e == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_382 <= _pht_T_3;
        end else begin
          pht_382 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_383 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h17f == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_383 <= _pht_T_3;
        end else begin
          pht_383 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_384 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h180 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_384 <= _pht_T_3;
        end else begin
          pht_384 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_385 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h181 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_385 <= _pht_T_3;
        end else begin
          pht_385 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_386 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h182 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_386 <= _pht_T_3;
        end else begin
          pht_386 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_387 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h183 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_387 <= _pht_T_3;
        end else begin
          pht_387 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_388 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h184 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_388 <= _pht_T_3;
        end else begin
          pht_388 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_389 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h185 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_389 <= _pht_T_3;
        end else begin
          pht_389 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_390 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h186 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_390 <= _pht_T_3;
        end else begin
          pht_390 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_391 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h187 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_391 <= _pht_T_3;
        end else begin
          pht_391 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_392 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h188 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_392 <= _pht_T_3;
        end else begin
          pht_392 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_393 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h189 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_393 <= _pht_T_3;
        end else begin
          pht_393 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_394 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h18a == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_394 <= _pht_T_3;
        end else begin
          pht_394 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_395 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h18b == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_395 <= _pht_T_3;
        end else begin
          pht_395 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_396 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h18c == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_396 <= _pht_T_3;
        end else begin
          pht_396 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_397 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h18d == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_397 <= _pht_T_3;
        end else begin
          pht_397 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_398 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h18e == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_398 <= _pht_T_3;
        end else begin
          pht_398 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_399 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h18f == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_399 <= _pht_T_3;
        end else begin
          pht_399 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_400 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h190 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_400 <= _pht_T_3;
        end else begin
          pht_400 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_401 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h191 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_401 <= _pht_T_3;
        end else begin
          pht_401 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_402 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h192 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_402 <= _pht_T_3;
        end else begin
          pht_402 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_403 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h193 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_403 <= _pht_T_3;
        end else begin
          pht_403 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_404 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h194 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_404 <= _pht_T_3;
        end else begin
          pht_404 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_405 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h195 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_405 <= _pht_T_3;
        end else begin
          pht_405 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_406 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h196 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_406 <= _pht_T_3;
        end else begin
          pht_406 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_407 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h197 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_407 <= _pht_T_3;
        end else begin
          pht_407 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_408 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h198 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_408 <= _pht_T_3;
        end else begin
          pht_408 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_409 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h199 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_409 <= _pht_T_3;
        end else begin
          pht_409 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_410 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h19a == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_410 <= _pht_T_3;
        end else begin
          pht_410 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_411 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h19b == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_411 <= _pht_T_3;
        end else begin
          pht_411 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_412 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h19c == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_412 <= _pht_T_3;
        end else begin
          pht_412 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_413 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h19d == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_413 <= _pht_T_3;
        end else begin
          pht_413 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_414 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h19e == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_414 <= _pht_T_3;
        end else begin
          pht_414 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_415 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h19f == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_415 <= _pht_T_3;
        end else begin
          pht_415 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_416 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1a0 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_416 <= _pht_T_3;
        end else begin
          pht_416 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_417 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1a1 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_417 <= _pht_T_3;
        end else begin
          pht_417 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_418 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1a2 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_418 <= _pht_T_3;
        end else begin
          pht_418 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_419 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1a3 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_419 <= _pht_T_3;
        end else begin
          pht_419 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_420 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1a4 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_420 <= _pht_T_3;
        end else begin
          pht_420 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_421 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1a5 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_421 <= _pht_T_3;
        end else begin
          pht_421 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_422 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1a6 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_422 <= _pht_T_3;
        end else begin
          pht_422 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_423 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1a7 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_423 <= _pht_T_3;
        end else begin
          pht_423 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_424 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1a8 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_424 <= _pht_T_3;
        end else begin
          pht_424 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_425 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1a9 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_425 <= _pht_T_3;
        end else begin
          pht_425 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_426 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1aa == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_426 <= _pht_T_3;
        end else begin
          pht_426 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_427 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1ab == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_427 <= _pht_T_3;
        end else begin
          pht_427 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_428 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1ac == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_428 <= _pht_T_3;
        end else begin
          pht_428 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_429 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1ad == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_429 <= _pht_T_3;
        end else begin
          pht_429 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_430 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1ae == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_430 <= _pht_T_3;
        end else begin
          pht_430 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_431 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1af == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_431 <= _pht_T_3;
        end else begin
          pht_431 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_432 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1b0 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_432 <= _pht_T_3;
        end else begin
          pht_432 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_433 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1b1 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_433 <= _pht_T_3;
        end else begin
          pht_433 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_434 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1b2 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_434 <= _pht_T_3;
        end else begin
          pht_434 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_435 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1b3 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_435 <= _pht_T_3;
        end else begin
          pht_435 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_436 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1b4 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_436 <= _pht_T_3;
        end else begin
          pht_436 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_437 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1b5 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_437 <= _pht_T_3;
        end else begin
          pht_437 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_438 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1b6 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_438 <= _pht_T_3;
        end else begin
          pht_438 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_439 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1b7 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_439 <= _pht_T_3;
        end else begin
          pht_439 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_440 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1b8 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_440 <= _pht_T_3;
        end else begin
          pht_440 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_441 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1b9 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_441 <= _pht_T_3;
        end else begin
          pht_441 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_442 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1ba == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_442 <= _pht_T_3;
        end else begin
          pht_442 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_443 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1bb == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_443 <= _pht_T_3;
        end else begin
          pht_443 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_444 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1bc == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_444 <= _pht_T_3;
        end else begin
          pht_444 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_445 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1bd == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_445 <= _pht_T_3;
        end else begin
          pht_445 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_446 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1be == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_446 <= _pht_T_3;
        end else begin
          pht_446 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_447 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1bf == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_447 <= _pht_T_3;
        end else begin
          pht_447 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_448 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1c0 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_448 <= _pht_T_3;
        end else begin
          pht_448 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_449 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1c1 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_449 <= _pht_T_3;
        end else begin
          pht_449 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_450 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1c2 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_450 <= _pht_T_3;
        end else begin
          pht_450 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_451 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1c3 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_451 <= _pht_T_3;
        end else begin
          pht_451 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_452 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1c4 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_452 <= _pht_T_3;
        end else begin
          pht_452 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_453 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1c5 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_453 <= _pht_T_3;
        end else begin
          pht_453 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_454 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1c6 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_454 <= _pht_T_3;
        end else begin
          pht_454 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_455 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1c7 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_455 <= _pht_T_3;
        end else begin
          pht_455 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_456 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1c8 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_456 <= _pht_T_3;
        end else begin
          pht_456 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_457 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1c9 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_457 <= _pht_T_3;
        end else begin
          pht_457 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_458 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1ca == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_458 <= _pht_T_3;
        end else begin
          pht_458 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_459 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1cb == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_459 <= _pht_T_3;
        end else begin
          pht_459 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_460 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1cc == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_460 <= _pht_T_3;
        end else begin
          pht_460 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_461 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1cd == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_461 <= _pht_T_3;
        end else begin
          pht_461 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_462 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1ce == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_462 <= _pht_T_3;
        end else begin
          pht_462 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_463 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1cf == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_463 <= _pht_T_3;
        end else begin
          pht_463 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_464 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1d0 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_464 <= _pht_T_3;
        end else begin
          pht_464 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_465 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1d1 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_465 <= _pht_T_3;
        end else begin
          pht_465 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_466 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1d2 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_466 <= _pht_T_3;
        end else begin
          pht_466 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_467 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1d3 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_467 <= _pht_T_3;
        end else begin
          pht_467 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_468 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1d4 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_468 <= _pht_T_3;
        end else begin
          pht_468 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_469 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1d5 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_469 <= _pht_T_3;
        end else begin
          pht_469 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_470 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1d6 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_470 <= _pht_T_3;
        end else begin
          pht_470 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_471 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1d7 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_471 <= _pht_T_3;
        end else begin
          pht_471 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_472 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1d8 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_472 <= _pht_T_3;
        end else begin
          pht_472 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_473 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1d9 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_473 <= _pht_T_3;
        end else begin
          pht_473 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_474 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1da == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_474 <= _pht_T_3;
        end else begin
          pht_474 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_475 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1db == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_475 <= _pht_T_3;
        end else begin
          pht_475 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_476 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1dc == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_476 <= _pht_T_3;
        end else begin
          pht_476 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_477 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1dd == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_477 <= _pht_T_3;
        end else begin
          pht_477 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_478 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1de == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_478 <= _pht_T_3;
        end else begin
          pht_478 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_479 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1df == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_479 <= _pht_T_3;
        end else begin
          pht_479 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_480 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1e0 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_480 <= _pht_T_3;
        end else begin
          pht_480 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_481 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1e1 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_481 <= _pht_T_3;
        end else begin
          pht_481 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_482 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1e2 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_482 <= _pht_T_3;
        end else begin
          pht_482 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_483 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1e3 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_483 <= _pht_T_3;
        end else begin
          pht_483 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_484 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1e4 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_484 <= _pht_T_3;
        end else begin
          pht_484 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_485 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1e5 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_485 <= _pht_T_3;
        end else begin
          pht_485 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_486 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1e6 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_486 <= _pht_T_3;
        end else begin
          pht_486 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_487 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1e7 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_487 <= _pht_T_3;
        end else begin
          pht_487 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_488 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1e8 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_488 <= _pht_T_3;
        end else begin
          pht_488 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_489 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1e9 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_489 <= _pht_T_3;
        end else begin
          pht_489 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_490 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1ea == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_490 <= _pht_T_3;
        end else begin
          pht_490 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_491 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1eb == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_491 <= _pht_T_3;
        end else begin
          pht_491 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_492 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1ec == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_492 <= _pht_T_3;
        end else begin
          pht_492 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_493 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1ed == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_493 <= _pht_T_3;
        end else begin
          pht_493 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_494 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1ee == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_494 <= _pht_T_3;
        end else begin
          pht_494 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_495 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1ef == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_495 <= _pht_T_3;
        end else begin
          pht_495 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_496 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1f0 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_496 <= _pht_T_3;
        end else begin
          pht_496 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_497 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1f1 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_497 <= _pht_T_3;
        end else begin
          pht_497 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_498 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1f2 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_498 <= _pht_T_3;
        end else begin
          pht_498 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_499 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1f3 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_499 <= _pht_T_3;
        end else begin
          pht_499 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_500 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1f4 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_500 <= _pht_T_3;
        end else begin
          pht_500 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_501 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1f5 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_501 <= _pht_T_3;
        end else begin
          pht_501 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_502 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1f6 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_502 <= _pht_T_3;
        end else begin
          pht_502 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_503 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1f7 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_503 <= _pht_T_3;
        end else begin
          pht_503 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_504 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1f8 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_504 <= _pht_T_3;
        end else begin
          pht_504 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_505 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1f9 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_505 <= _pht_T_3;
        end else begin
          pht_505 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_506 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1fa == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_506 <= _pht_T_3;
        end else begin
          pht_506 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_507 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1fb == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_507 <= _pht_T_3;
        end else begin
          pht_507 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_508 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1fc == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_508 <= _pht_T_3;
        end else begin
          pht_508 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_509 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1fd == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_509 <= _pht_T_3;
        end else begin
          pht_509 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_510 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1fe == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_510 <= _pht_T_3;
        end else begin
          pht_510 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_511 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1ff == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_511 <= _pht_T_3;
        end else begin
          pht_511 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_0_tag <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'h0 == btb_replace_idx) begin // @[BPU.scala 80:33]
        btb_0_tag <= io_jmp_packet_bp_pc[38:2]; // @[BPU.scala 80:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_0_target <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'h0 == btb_replace_idx) begin // @[BPU.scala 81:33]
        btb_0_target <= io_jmp_packet_target[38:2]; // @[BPU.scala 81:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_0_valid <= 1'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      btb_0_valid <= _GEN_2114;
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_1_tag <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'h1 == btb_replace_idx) begin // @[BPU.scala 80:33]
        btb_1_tag <= io_jmp_packet_bp_pc[38:2]; // @[BPU.scala 80:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_1_target <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'h1 == btb_replace_idx) begin // @[BPU.scala 81:33]
        btb_1_target <= io_jmp_packet_target[38:2]; // @[BPU.scala 81:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_1_valid <= 1'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      btb_1_valid <= _GEN_2115;
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_2_tag <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'h2 == btb_replace_idx) begin // @[BPU.scala 80:33]
        btb_2_tag <= io_jmp_packet_bp_pc[38:2]; // @[BPU.scala 80:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_2_target <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'h2 == btb_replace_idx) begin // @[BPU.scala 81:33]
        btb_2_target <= io_jmp_packet_target[38:2]; // @[BPU.scala 81:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_2_valid <= 1'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      btb_2_valid <= _GEN_2116;
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_3_tag <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'h3 == btb_replace_idx) begin // @[BPU.scala 80:33]
        btb_3_tag <= io_jmp_packet_bp_pc[38:2]; // @[BPU.scala 80:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_3_target <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'h3 == btb_replace_idx) begin // @[BPU.scala 81:33]
        btb_3_target <= io_jmp_packet_target[38:2]; // @[BPU.scala 81:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_3_valid <= 1'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      btb_3_valid <= _GEN_2117;
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_4_tag <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'h4 == btb_replace_idx) begin // @[BPU.scala 80:33]
        btb_4_tag <= io_jmp_packet_bp_pc[38:2]; // @[BPU.scala 80:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_4_target <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'h4 == btb_replace_idx) begin // @[BPU.scala 81:33]
        btb_4_target <= io_jmp_packet_target[38:2]; // @[BPU.scala 81:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_4_valid <= 1'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      btb_4_valid <= _GEN_2118;
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_5_tag <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'h5 == btb_replace_idx) begin // @[BPU.scala 80:33]
        btb_5_tag <= io_jmp_packet_bp_pc[38:2]; // @[BPU.scala 80:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_5_target <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'h5 == btb_replace_idx) begin // @[BPU.scala 81:33]
        btb_5_target <= io_jmp_packet_target[38:2]; // @[BPU.scala 81:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_5_valid <= 1'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      btb_5_valid <= _GEN_2119;
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_6_tag <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'h6 == btb_replace_idx) begin // @[BPU.scala 80:33]
        btb_6_tag <= io_jmp_packet_bp_pc[38:2]; // @[BPU.scala 80:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_6_target <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'h6 == btb_replace_idx) begin // @[BPU.scala 81:33]
        btb_6_target <= io_jmp_packet_target[38:2]; // @[BPU.scala 81:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_6_valid <= 1'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      btb_6_valid <= _GEN_2120;
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_7_tag <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'h7 == btb_replace_idx) begin // @[BPU.scala 80:33]
        btb_7_tag <= io_jmp_packet_bp_pc[38:2]; // @[BPU.scala 80:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_7_target <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'h7 == btb_replace_idx) begin // @[BPU.scala 81:33]
        btb_7_target <= io_jmp_packet_target[38:2]; // @[BPU.scala 81:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_7_valid <= 1'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      btb_7_valid <= _GEN_2121;
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_8_tag <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'h8 == btb_replace_idx) begin // @[BPU.scala 80:33]
        btb_8_tag <= io_jmp_packet_bp_pc[38:2]; // @[BPU.scala 80:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_8_target <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'h8 == btb_replace_idx) begin // @[BPU.scala 81:33]
        btb_8_target <= io_jmp_packet_target[38:2]; // @[BPU.scala 81:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_8_valid <= 1'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      btb_8_valid <= _GEN_2122;
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_9_tag <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'h9 == btb_replace_idx) begin // @[BPU.scala 80:33]
        btb_9_tag <= io_jmp_packet_bp_pc[38:2]; // @[BPU.scala 80:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_9_target <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'h9 == btb_replace_idx) begin // @[BPU.scala 81:33]
        btb_9_target <= io_jmp_packet_target[38:2]; // @[BPU.scala 81:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_9_valid <= 1'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      btb_9_valid <= _GEN_2123;
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_10_tag <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'ha == btb_replace_idx) begin // @[BPU.scala 80:33]
        btb_10_tag <= io_jmp_packet_bp_pc[38:2]; // @[BPU.scala 80:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_10_target <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'ha == btb_replace_idx) begin // @[BPU.scala 81:33]
        btb_10_target <= io_jmp_packet_target[38:2]; // @[BPU.scala 81:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_10_valid <= 1'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      btb_10_valid <= _GEN_2124;
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_11_tag <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'hb == btb_replace_idx) begin // @[BPU.scala 80:33]
        btb_11_tag <= io_jmp_packet_bp_pc[38:2]; // @[BPU.scala 80:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_11_target <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'hb == btb_replace_idx) begin // @[BPU.scala 81:33]
        btb_11_target <= io_jmp_packet_target[38:2]; // @[BPU.scala 81:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_11_valid <= 1'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      btb_11_valid <= _GEN_2125;
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_12_tag <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'hc == btb_replace_idx) begin // @[BPU.scala 80:33]
        btb_12_tag <= io_jmp_packet_bp_pc[38:2]; // @[BPU.scala 80:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_12_target <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'hc == btb_replace_idx) begin // @[BPU.scala 81:33]
        btb_12_target <= io_jmp_packet_target[38:2]; // @[BPU.scala 81:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_12_valid <= 1'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      btb_12_valid <= _GEN_2126;
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_13_tag <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'hd == btb_replace_idx) begin // @[BPU.scala 80:33]
        btb_13_tag <= io_jmp_packet_bp_pc[38:2]; // @[BPU.scala 80:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_13_target <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'hd == btb_replace_idx) begin // @[BPU.scala 81:33]
        btb_13_target <= io_jmp_packet_target[38:2]; // @[BPU.scala 81:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_13_valid <= 1'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      btb_13_valid <= _GEN_2127;
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_14_tag <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'he == btb_replace_idx) begin // @[BPU.scala 80:33]
        btb_14_tag <= io_jmp_packet_bp_pc[38:2]; // @[BPU.scala 80:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_14_target <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'he == btb_replace_idx) begin // @[BPU.scala 81:33]
        btb_14_target <= io_jmp_packet_target[38:2]; // @[BPU.scala 81:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_14_valid <= 1'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      btb_14_valid <= _GEN_2128;
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_15_tag <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'hf == btb_replace_idx) begin // @[BPU.scala 80:33]
        btb_15_tag <= io_jmp_packet_bp_pc[38:2]; // @[BPU.scala 80:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_15_target <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'hf == btb_replace_idx) begin // @[BPU.scala 81:33]
        btb_15_target <= io_jmp_packet_target[38:2]; // @[BPU.scala 81:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_15_valid <= 1'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      btb_15_valid <= _GEN_2129;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ghr = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  pht_0 = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  pht_1 = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  pht_2 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  pht_3 = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  pht_4 = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  pht_5 = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  pht_6 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  pht_7 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  pht_8 = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  pht_9 = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  pht_10 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  pht_11 = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  pht_12 = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  pht_13 = _RAND_14[1:0];
  _RAND_15 = {1{`RANDOM}};
  pht_14 = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  pht_15 = _RAND_16[1:0];
  _RAND_17 = {1{`RANDOM}};
  pht_16 = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  pht_17 = _RAND_18[1:0];
  _RAND_19 = {1{`RANDOM}};
  pht_18 = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  pht_19 = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  pht_20 = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  pht_21 = _RAND_22[1:0];
  _RAND_23 = {1{`RANDOM}};
  pht_22 = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  pht_23 = _RAND_24[1:0];
  _RAND_25 = {1{`RANDOM}};
  pht_24 = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  pht_25 = _RAND_26[1:0];
  _RAND_27 = {1{`RANDOM}};
  pht_26 = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  pht_27 = _RAND_28[1:0];
  _RAND_29 = {1{`RANDOM}};
  pht_28 = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  pht_29 = _RAND_30[1:0];
  _RAND_31 = {1{`RANDOM}};
  pht_30 = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  pht_31 = _RAND_32[1:0];
  _RAND_33 = {1{`RANDOM}};
  pht_32 = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  pht_33 = _RAND_34[1:0];
  _RAND_35 = {1{`RANDOM}};
  pht_34 = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  pht_35 = _RAND_36[1:0];
  _RAND_37 = {1{`RANDOM}};
  pht_36 = _RAND_37[1:0];
  _RAND_38 = {1{`RANDOM}};
  pht_37 = _RAND_38[1:0];
  _RAND_39 = {1{`RANDOM}};
  pht_38 = _RAND_39[1:0];
  _RAND_40 = {1{`RANDOM}};
  pht_39 = _RAND_40[1:0];
  _RAND_41 = {1{`RANDOM}};
  pht_40 = _RAND_41[1:0];
  _RAND_42 = {1{`RANDOM}};
  pht_41 = _RAND_42[1:0];
  _RAND_43 = {1{`RANDOM}};
  pht_42 = _RAND_43[1:0];
  _RAND_44 = {1{`RANDOM}};
  pht_43 = _RAND_44[1:0];
  _RAND_45 = {1{`RANDOM}};
  pht_44 = _RAND_45[1:0];
  _RAND_46 = {1{`RANDOM}};
  pht_45 = _RAND_46[1:0];
  _RAND_47 = {1{`RANDOM}};
  pht_46 = _RAND_47[1:0];
  _RAND_48 = {1{`RANDOM}};
  pht_47 = _RAND_48[1:0];
  _RAND_49 = {1{`RANDOM}};
  pht_48 = _RAND_49[1:0];
  _RAND_50 = {1{`RANDOM}};
  pht_49 = _RAND_50[1:0];
  _RAND_51 = {1{`RANDOM}};
  pht_50 = _RAND_51[1:0];
  _RAND_52 = {1{`RANDOM}};
  pht_51 = _RAND_52[1:0];
  _RAND_53 = {1{`RANDOM}};
  pht_52 = _RAND_53[1:0];
  _RAND_54 = {1{`RANDOM}};
  pht_53 = _RAND_54[1:0];
  _RAND_55 = {1{`RANDOM}};
  pht_54 = _RAND_55[1:0];
  _RAND_56 = {1{`RANDOM}};
  pht_55 = _RAND_56[1:0];
  _RAND_57 = {1{`RANDOM}};
  pht_56 = _RAND_57[1:0];
  _RAND_58 = {1{`RANDOM}};
  pht_57 = _RAND_58[1:0];
  _RAND_59 = {1{`RANDOM}};
  pht_58 = _RAND_59[1:0];
  _RAND_60 = {1{`RANDOM}};
  pht_59 = _RAND_60[1:0];
  _RAND_61 = {1{`RANDOM}};
  pht_60 = _RAND_61[1:0];
  _RAND_62 = {1{`RANDOM}};
  pht_61 = _RAND_62[1:0];
  _RAND_63 = {1{`RANDOM}};
  pht_62 = _RAND_63[1:0];
  _RAND_64 = {1{`RANDOM}};
  pht_63 = _RAND_64[1:0];
  _RAND_65 = {1{`RANDOM}};
  pht_64 = _RAND_65[1:0];
  _RAND_66 = {1{`RANDOM}};
  pht_65 = _RAND_66[1:0];
  _RAND_67 = {1{`RANDOM}};
  pht_66 = _RAND_67[1:0];
  _RAND_68 = {1{`RANDOM}};
  pht_67 = _RAND_68[1:0];
  _RAND_69 = {1{`RANDOM}};
  pht_68 = _RAND_69[1:0];
  _RAND_70 = {1{`RANDOM}};
  pht_69 = _RAND_70[1:0];
  _RAND_71 = {1{`RANDOM}};
  pht_70 = _RAND_71[1:0];
  _RAND_72 = {1{`RANDOM}};
  pht_71 = _RAND_72[1:0];
  _RAND_73 = {1{`RANDOM}};
  pht_72 = _RAND_73[1:0];
  _RAND_74 = {1{`RANDOM}};
  pht_73 = _RAND_74[1:0];
  _RAND_75 = {1{`RANDOM}};
  pht_74 = _RAND_75[1:0];
  _RAND_76 = {1{`RANDOM}};
  pht_75 = _RAND_76[1:0];
  _RAND_77 = {1{`RANDOM}};
  pht_76 = _RAND_77[1:0];
  _RAND_78 = {1{`RANDOM}};
  pht_77 = _RAND_78[1:0];
  _RAND_79 = {1{`RANDOM}};
  pht_78 = _RAND_79[1:0];
  _RAND_80 = {1{`RANDOM}};
  pht_79 = _RAND_80[1:0];
  _RAND_81 = {1{`RANDOM}};
  pht_80 = _RAND_81[1:0];
  _RAND_82 = {1{`RANDOM}};
  pht_81 = _RAND_82[1:0];
  _RAND_83 = {1{`RANDOM}};
  pht_82 = _RAND_83[1:0];
  _RAND_84 = {1{`RANDOM}};
  pht_83 = _RAND_84[1:0];
  _RAND_85 = {1{`RANDOM}};
  pht_84 = _RAND_85[1:0];
  _RAND_86 = {1{`RANDOM}};
  pht_85 = _RAND_86[1:0];
  _RAND_87 = {1{`RANDOM}};
  pht_86 = _RAND_87[1:0];
  _RAND_88 = {1{`RANDOM}};
  pht_87 = _RAND_88[1:0];
  _RAND_89 = {1{`RANDOM}};
  pht_88 = _RAND_89[1:0];
  _RAND_90 = {1{`RANDOM}};
  pht_89 = _RAND_90[1:0];
  _RAND_91 = {1{`RANDOM}};
  pht_90 = _RAND_91[1:0];
  _RAND_92 = {1{`RANDOM}};
  pht_91 = _RAND_92[1:0];
  _RAND_93 = {1{`RANDOM}};
  pht_92 = _RAND_93[1:0];
  _RAND_94 = {1{`RANDOM}};
  pht_93 = _RAND_94[1:0];
  _RAND_95 = {1{`RANDOM}};
  pht_94 = _RAND_95[1:0];
  _RAND_96 = {1{`RANDOM}};
  pht_95 = _RAND_96[1:0];
  _RAND_97 = {1{`RANDOM}};
  pht_96 = _RAND_97[1:0];
  _RAND_98 = {1{`RANDOM}};
  pht_97 = _RAND_98[1:0];
  _RAND_99 = {1{`RANDOM}};
  pht_98 = _RAND_99[1:0];
  _RAND_100 = {1{`RANDOM}};
  pht_99 = _RAND_100[1:0];
  _RAND_101 = {1{`RANDOM}};
  pht_100 = _RAND_101[1:0];
  _RAND_102 = {1{`RANDOM}};
  pht_101 = _RAND_102[1:0];
  _RAND_103 = {1{`RANDOM}};
  pht_102 = _RAND_103[1:0];
  _RAND_104 = {1{`RANDOM}};
  pht_103 = _RAND_104[1:0];
  _RAND_105 = {1{`RANDOM}};
  pht_104 = _RAND_105[1:0];
  _RAND_106 = {1{`RANDOM}};
  pht_105 = _RAND_106[1:0];
  _RAND_107 = {1{`RANDOM}};
  pht_106 = _RAND_107[1:0];
  _RAND_108 = {1{`RANDOM}};
  pht_107 = _RAND_108[1:0];
  _RAND_109 = {1{`RANDOM}};
  pht_108 = _RAND_109[1:0];
  _RAND_110 = {1{`RANDOM}};
  pht_109 = _RAND_110[1:0];
  _RAND_111 = {1{`RANDOM}};
  pht_110 = _RAND_111[1:0];
  _RAND_112 = {1{`RANDOM}};
  pht_111 = _RAND_112[1:0];
  _RAND_113 = {1{`RANDOM}};
  pht_112 = _RAND_113[1:0];
  _RAND_114 = {1{`RANDOM}};
  pht_113 = _RAND_114[1:0];
  _RAND_115 = {1{`RANDOM}};
  pht_114 = _RAND_115[1:0];
  _RAND_116 = {1{`RANDOM}};
  pht_115 = _RAND_116[1:0];
  _RAND_117 = {1{`RANDOM}};
  pht_116 = _RAND_117[1:0];
  _RAND_118 = {1{`RANDOM}};
  pht_117 = _RAND_118[1:0];
  _RAND_119 = {1{`RANDOM}};
  pht_118 = _RAND_119[1:0];
  _RAND_120 = {1{`RANDOM}};
  pht_119 = _RAND_120[1:0];
  _RAND_121 = {1{`RANDOM}};
  pht_120 = _RAND_121[1:0];
  _RAND_122 = {1{`RANDOM}};
  pht_121 = _RAND_122[1:0];
  _RAND_123 = {1{`RANDOM}};
  pht_122 = _RAND_123[1:0];
  _RAND_124 = {1{`RANDOM}};
  pht_123 = _RAND_124[1:0];
  _RAND_125 = {1{`RANDOM}};
  pht_124 = _RAND_125[1:0];
  _RAND_126 = {1{`RANDOM}};
  pht_125 = _RAND_126[1:0];
  _RAND_127 = {1{`RANDOM}};
  pht_126 = _RAND_127[1:0];
  _RAND_128 = {1{`RANDOM}};
  pht_127 = _RAND_128[1:0];
  _RAND_129 = {1{`RANDOM}};
  pht_128 = _RAND_129[1:0];
  _RAND_130 = {1{`RANDOM}};
  pht_129 = _RAND_130[1:0];
  _RAND_131 = {1{`RANDOM}};
  pht_130 = _RAND_131[1:0];
  _RAND_132 = {1{`RANDOM}};
  pht_131 = _RAND_132[1:0];
  _RAND_133 = {1{`RANDOM}};
  pht_132 = _RAND_133[1:0];
  _RAND_134 = {1{`RANDOM}};
  pht_133 = _RAND_134[1:0];
  _RAND_135 = {1{`RANDOM}};
  pht_134 = _RAND_135[1:0];
  _RAND_136 = {1{`RANDOM}};
  pht_135 = _RAND_136[1:0];
  _RAND_137 = {1{`RANDOM}};
  pht_136 = _RAND_137[1:0];
  _RAND_138 = {1{`RANDOM}};
  pht_137 = _RAND_138[1:0];
  _RAND_139 = {1{`RANDOM}};
  pht_138 = _RAND_139[1:0];
  _RAND_140 = {1{`RANDOM}};
  pht_139 = _RAND_140[1:0];
  _RAND_141 = {1{`RANDOM}};
  pht_140 = _RAND_141[1:0];
  _RAND_142 = {1{`RANDOM}};
  pht_141 = _RAND_142[1:0];
  _RAND_143 = {1{`RANDOM}};
  pht_142 = _RAND_143[1:0];
  _RAND_144 = {1{`RANDOM}};
  pht_143 = _RAND_144[1:0];
  _RAND_145 = {1{`RANDOM}};
  pht_144 = _RAND_145[1:0];
  _RAND_146 = {1{`RANDOM}};
  pht_145 = _RAND_146[1:0];
  _RAND_147 = {1{`RANDOM}};
  pht_146 = _RAND_147[1:0];
  _RAND_148 = {1{`RANDOM}};
  pht_147 = _RAND_148[1:0];
  _RAND_149 = {1{`RANDOM}};
  pht_148 = _RAND_149[1:0];
  _RAND_150 = {1{`RANDOM}};
  pht_149 = _RAND_150[1:0];
  _RAND_151 = {1{`RANDOM}};
  pht_150 = _RAND_151[1:0];
  _RAND_152 = {1{`RANDOM}};
  pht_151 = _RAND_152[1:0];
  _RAND_153 = {1{`RANDOM}};
  pht_152 = _RAND_153[1:0];
  _RAND_154 = {1{`RANDOM}};
  pht_153 = _RAND_154[1:0];
  _RAND_155 = {1{`RANDOM}};
  pht_154 = _RAND_155[1:0];
  _RAND_156 = {1{`RANDOM}};
  pht_155 = _RAND_156[1:0];
  _RAND_157 = {1{`RANDOM}};
  pht_156 = _RAND_157[1:0];
  _RAND_158 = {1{`RANDOM}};
  pht_157 = _RAND_158[1:0];
  _RAND_159 = {1{`RANDOM}};
  pht_158 = _RAND_159[1:0];
  _RAND_160 = {1{`RANDOM}};
  pht_159 = _RAND_160[1:0];
  _RAND_161 = {1{`RANDOM}};
  pht_160 = _RAND_161[1:0];
  _RAND_162 = {1{`RANDOM}};
  pht_161 = _RAND_162[1:0];
  _RAND_163 = {1{`RANDOM}};
  pht_162 = _RAND_163[1:0];
  _RAND_164 = {1{`RANDOM}};
  pht_163 = _RAND_164[1:0];
  _RAND_165 = {1{`RANDOM}};
  pht_164 = _RAND_165[1:0];
  _RAND_166 = {1{`RANDOM}};
  pht_165 = _RAND_166[1:0];
  _RAND_167 = {1{`RANDOM}};
  pht_166 = _RAND_167[1:0];
  _RAND_168 = {1{`RANDOM}};
  pht_167 = _RAND_168[1:0];
  _RAND_169 = {1{`RANDOM}};
  pht_168 = _RAND_169[1:0];
  _RAND_170 = {1{`RANDOM}};
  pht_169 = _RAND_170[1:0];
  _RAND_171 = {1{`RANDOM}};
  pht_170 = _RAND_171[1:0];
  _RAND_172 = {1{`RANDOM}};
  pht_171 = _RAND_172[1:0];
  _RAND_173 = {1{`RANDOM}};
  pht_172 = _RAND_173[1:0];
  _RAND_174 = {1{`RANDOM}};
  pht_173 = _RAND_174[1:0];
  _RAND_175 = {1{`RANDOM}};
  pht_174 = _RAND_175[1:0];
  _RAND_176 = {1{`RANDOM}};
  pht_175 = _RAND_176[1:0];
  _RAND_177 = {1{`RANDOM}};
  pht_176 = _RAND_177[1:0];
  _RAND_178 = {1{`RANDOM}};
  pht_177 = _RAND_178[1:0];
  _RAND_179 = {1{`RANDOM}};
  pht_178 = _RAND_179[1:0];
  _RAND_180 = {1{`RANDOM}};
  pht_179 = _RAND_180[1:0];
  _RAND_181 = {1{`RANDOM}};
  pht_180 = _RAND_181[1:0];
  _RAND_182 = {1{`RANDOM}};
  pht_181 = _RAND_182[1:0];
  _RAND_183 = {1{`RANDOM}};
  pht_182 = _RAND_183[1:0];
  _RAND_184 = {1{`RANDOM}};
  pht_183 = _RAND_184[1:0];
  _RAND_185 = {1{`RANDOM}};
  pht_184 = _RAND_185[1:0];
  _RAND_186 = {1{`RANDOM}};
  pht_185 = _RAND_186[1:0];
  _RAND_187 = {1{`RANDOM}};
  pht_186 = _RAND_187[1:0];
  _RAND_188 = {1{`RANDOM}};
  pht_187 = _RAND_188[1:0];
  _RAND_189 = {1{`RANDOM}};
  pht_188 = _RAND_189[1:0];
  _RAND_190 = {1{`RANDOM}};
  pht_189 = _RAND_190[1:0];
  _RAND_191 = {1{`RANDOM}};
  pht_190 = _RAND_191[1:0];
  _RAND_192 = {1{`RANDOM}};
  pht_191 = _RAND_192[1:0];
  _RAND_193 = {1{`RANDOM}};
  pht_192 = _RAND_193[1:0];
  _RAND_194 = {1{`RANDOM}};
  pht_193 = _RAND_194[1:0];
  _RAND_195 = {1{`RANDOM}};
  pht_194 = _RAND_195[1:0];
  _RAND_196 = {1{`RANDOM}};
  pht_195 = _RAND_196[1:0];
  _RAND_197 = {1{`RANDOM}};
  pht_196 = _RAND_197[1:0];
  _RAND_198 = {1{`RANDOM}};
  pht_197 = _RAND_198[1:0];
  _RAND_199 = {1{`RANDOM}};
  pht_198 = _RAND_199[1:0];
  _RAND_200 = {1{`RANDOM}};
  pht_199 = _RAND_200[1:0];
  _RAND_201 = {1{`RANDOM}};
  pht_200 = _RAND_201[1:0];
  _RAND_202 = {1{`RANDOM}};
  pht_201 = _RAND_202[1:0];
  _RAND_203 = {1{`RANDOM}};
  pht_202 = _RAND_203[1:0];
  _RAND_204 = {1{`RANDOM}};
  pht_203 = _RAND_204[1:0];
  _RAND_205 = {1{`RANDOM}};
  pht_204 = _RAND_205[1:0];
  _RAND_206 = {1{`RANDOM}};
  pht_205 = _RAND_206[1:0];
  _RAND_207 = {1{`RANDOM}};
  pht_206 = _RAND_207[1:0];
  _RAND_208 = {1{`RANDOM}};
  pht_207 = _RAND_208[1:0];
  _RAND_209 = {1{`RANDOM}};
  pht_208 = _RAND_209[1:0];
  _RAND_210 = {1{`RANDOM}};
  pht_209 = _RAND_210[1:0];
  _RAND_211 = {1{`RANDOM}};
  pht_210 = _RAND_211[1:0];
  _RAND_212 = {1{`RANDOM}};
  pht_211 = _RAND_212[1:0];
  _RAND_213 = {1{`RANDOM}};
  pht_212 = _RAND_213[1:0];
  _RAND_214 = {1{`RANDOM}};
  pht_213 = _RAND_214[1:0];
  _RAND_215 = {1{`RANDOM}};
  pht_214 = _RAND_215[1:0];
  _RAND_216 = {1{`RANDOM}};
  pht_215 = _RAND_216[1:0];
  _RAND_217 = {1{`RANDOM}};
  pht_216 = _RAND_217[1:0];
  _RAND_218 = {1{`RANDOM}};
  pht_217 = _RAND_218[1:0];
  _RAND_219 = {1{`RANDOM}};
  pht_218 = _RAND_219[1:0];
  _RAND_220 = {1{`RANDOM}};
  pht_219 = _RAND_220[1:0];
  _RAND_221 = {1{`RANDOM}};
  pht_220 = _RAND_221[1:0];
  _RAND_222 = {1{`RANDOM}};
  pht_221 = _RAND_222[1:0];
  _RAND_223 = {1{`RANDOM}};
  pht_222 = _RAND_223[1:0];
  _RAND_224 = {1{`RANDOM}};
  pht_223 = _RAND_224[1:0];
  _RAND_225 = {1{`RANDOM}};
  pht_224 = _RAND_225[1:0];
  _RAND_226 = {1{`RANDOM}};
  pht_225 = _RAND_226[1:0];
  _RAND_227 = {1{`RANDOM}};
  pht_226 = _RAND_227[1:0];
  _RAND_228 = {1{`RANDOM}};
  pht_227 = _RAND_228[1:0];
  _RAND_229 = {1{`RANDOM}};
  pht_228 = _RAND_229[1:0];
  _RAND_230 = {1{`RANDOM}};
  pht_229 = _RAND_230[1:0];
  _RAND_231 = {1{`RANDOM}};
  pht_230 = _RAND_231[1:0];
  _RAND_232 = {1{`RANDOM}};
  pht_231 = _RAND_232[1:0];
  _RAND_233 = {1{`RANDOM}};
  pht_232 = _RAND_233[1:0];
  _RAND_234 = {1{`RANDOM}};
  pht_233 = _RAND_234[1:0];
  _RAND_235 = {1{`RANDOM}};
  pht_234 = _RAND_235[1:0];
  _RAND_236 = {1{`RANDOM}};
  pht_235 = _RAND_236[1:0];
  _RAND_237 = {1{`RANDOM}};
  pht_236 = _RAND_237[1:0];
  _RAND_238 = {1{`RANDOM}};
  pht_237 = _RAND_238[1:0];
  _RAND_239 = {1{`RANDOM}};
  pht_238 = _RAND_239[1:0];
  _RAND_240 = {1{`RANDOM}};
  pht_239 = _RAND_240[1:0];
  _RAND_241 = {1{`RANDOM}};
  pht_240 = _RAND_241[1:0];
  _RAND_242 = {1{`RANDOM}};
  pht_241 = _RAND_242[1:0];
  _RAND_243 = {1{`RANDOM}};
  pht_242 = _RAND_243[1:0];
  _RAND_244 = {1{`RANDOM}};
  pht_243 = _RAND_244[1:0];
  _RAND_245 = {1{`RANDOM}};
  pht_244 = _RAND_245[1:0];
  _RAND_246 = {1{`RANDOM}};
  pht_245 = _RAND_246[1:0];
  _RAND_247 = {1{`RANDOM}};
  pht_246 = _RAND_247[1:0];
  _RAND_248 = {1{`RANDOM}};
  pht_247 = _RAND_248[1:0];
  _RAND_249 = {1{`RANDOM}};
  pht_248 = _RAND_249[1:0];
  _RAND_250 = {1{`RANDOM}};
  pht_249 = _RAND_250[1:0];
  _RAND_251 = {1{`RANDOM}};
  pht_250 = _RAND_251[1:0];
  _RAND_252 = {1{`RANDOM}};
  pht_251 = _RAND_252[1:0];
  _RAND_253 = {1{`RANDOM}};
  pht_252 = _RAND_253[1:0];
  _RAND_254 = {1{`RANDOM}};
  pht_253 = _RAND_254[1:0];
  _RAND_255 = {1{`RANDOM}};
  pht_254 = _RAND_255[1:0];
  _RAND_256 = {1{`RANDOM}};
  pht_255 = _RAND_256[1:0];
  _RAND_257 = {1{`RANDOM}};
  pht_256 = _RAND_257[1:0];
  _RAND_258 = {1{`RANDOM}};
  pht_257 = _RAND_258[1:0];
  _RAND_259 = {1{`RANDOM}};
  pht_258 = _RAND_259[1:0];
  _RAND_260 = {1{`RANDOM}};
  pht_259 = _RAND_260[1:0];
  _RAND_261 = {1{`RANDOM}};
  pht_260 = _RAND_261[1:0];
  _RAND_262 = {1{`RANDOM}};
  pht_261 = _RAND_262[1:0];
  _RAND_263 = {1{`RANDOM}};
  pht_262 = _RAND_263[1:0];
  _RAND_264 = {1{`RANDOM}};
  pht_263 = _RAND_264[1:0];
  _RAND_265 = {1{`RANDOM}};
  pht_264 = _RAND_265[1:0];
  _RAND_266 = {1{`RANDOM}};
  pht_265 = _RAND_266[1:0];
  _RAND_267 = {1{`RANDOM}};
  pht_266 = _RAND_267[1:0];
  _RAND_268 = {1{`RANDOM}};
  pht_267 = _RAND_268[1:0];
  _RAND_269 = {1{`RANDOM}};
  pht_268 = _RAND_269[1:0];
  _RAND_270 = {1{`RANDOM}};
  pht_269 = _RAND_270[1:0];
  _RAND_271 = {1{`RANDOM}};
  pht_270 = _RAND_271[1:0];
  _RAND_272 = {1{`RANDOM}};
  pht_271 = _RAND_272[1:0];
  _RAND_273 = {1{`RANDOM}};
  pht_272 = _RAND_273[1:0];
  _RAND_274 = {1{`RANDOM}};
  pht_273 = _RAND_274[1:0];
  _RAND_275 = {1{`RANDOM}};
  pht_274 = _RAND_275[1:0];
  _RAND_276 = {1{`RANDOM}};
  pht_275 = _RAND_276[1:0];
  _RAND_277 = {1{`RANDOM}};
  pht_276 = _RAND_277[1:0];
  _RAND_278 = {1{`RANDOM}};
  pht_277 = _RAND_278[1:0];
  _RAND_279 = {1{`RANDOM}};
  pht_278 = _RAND_279[1:0];
  _RAND_280 = {1{`RANDOM}};
  pht_279 = _RAND_280[1:0];
  _RAND_281 = {1{`RANDOM}};
  pht_280 = _RAND_281[1:0];
  _RAND_282 = {1{`RANDOM}};
  pht_281 = _RAND_282[1:0];
  _RAND_283 = {1{`RANDOM}};
  pht_282 = _RAND_283[1:0];
  _RAND_284 = {1{`RANDOM}};
  pht_283 = _RAND_284[1:0];
  _RAND_285 = {1{`RANDOM}};
  pht_284 = _RAND_285[1:0];
  _RAND_286 = {1{`RANDOM}};
  pht_285 = _RAND_286[1:0];
  _RAND_287 = {1{`RANDOM}};
  pht_286 = _RAND_287[1:0];
  _RAND_288 = {1{`RANDOM}};
  pht_287 = _RAND_288[1:0];
  _RAND_289 = {1{`RANDOM}};
  pht_288 = _RAND_289[1:0];
  _RAND_290 = {1{`RANDOM}};
  pht_289 = _RAND_290[1:0];
  _RAND_291 = {1{`RANDOM}};
  pht_290 = _RAND_291[1:0];
  _RAND_292 = {1{`RANDOM}};
  pht_291 = _RAND_292[1:0];
  _RAND_293 = {1{`RANDOM}};
  pht_292 = _RAND_293[1:0];
  _RAND_294 = {1{`RANDOM}};
  pht_293 = _RAND_294[1:0];
  _RAND_295 = {1{`RANDOM}};
  pht_294 = _RAND_295[1:0];
  _RAND_296 = {1{`RANDOM}};
  pht_295 = _RAND_296[1:0];
  _RAND_297 = {1{`RANDOM}};
  pht_296 = _RAND_297[1:0];
  _RAND_298 = {1{`RANDOM}};
  pht_297 = _RAND_298[1:0];
  _RAND_299 = {1{`RANDOM}};
  pht_298 = _RAND_299[1:0];
  _RAND_300 = {1{`RANDOM}};
  pht_299 = _RAND_300[1:0];
  _RAND_301 = {1{`RANDOM}};
  pht_300 = _RAND_301[1:0];
  _RAND_302 = {1{`RANDOM}};
  pht_301 = _RAND_302[1:0];
  _RAND_303 = {1{`RANDOM}};
  pht_302 = _RAND_303[1:0];
  _RAND_304 = {1{`RANDOM}};
  pht_303 = _RAND_304[1:0];
  _RAND_305 = {1{`RANDOM}};
  pht_304 = _RAND_305[1:0];
  _RAND_306 = {1{`RANDOM}};
  pht_305 = _RAND_306[1:0];
  _RAND_307 = {1{`RANDOM}};
  pht_306 = _RAND_307[1:0];
  _RAND_308 = {1{`RANDOM}};
  pht_307 = _RAND_308[1:0];
  _RAND_309 = {1{`RANDOM}};
  pht_308 = _RAND_309[1:0];
  _RAND_310 = {1{`RANDOM}};
  pht_309 = _RAND_310[1:0];
  _RAND_311 = {1{`RANDOM}};
  pht_310 = _RAND_311[1:0];
  _RAND_312 = {1{`RANDOM}};
  pht_311 = _RAND_312[1:0];
  _RAND_313 = {1{`RANDOM}};
  pht_312 = _RAND_313[1:0];
  _RAND_314 = {1{`RANDOM}};
  pht_313 = _RAND_314[1:0];
  _RAND_315 = {1{`RANDOM}};
  pht_314 = _RAND_315[1:0];
  _RAND_316 = {1{`RANDOM}};
  pht_315 = _RAND_316[1:0];
  _RAND_317 = {1{`RANDOM}};
  pht_316 = _RAND_317[1:0];
  _RAND_318 = {1{`RANDOM}};
  pht_317 = _RAND_318[1:0];
  _RAND_319 = {1{`RANDOM}};
  pht_318 = _RAND_319[1:0];
  _RAND_320 = {1{`RANDOM}};
  pht_319 = _RAND_320[1:0];
  _RAND_321 = {1{`RANDOM}};
  pht_320 = _RAND_321[1:0];
  _RAND_322 = {1{`RANDOM}};
  pht_321 = _RAND_322[1:0];
  _RAND_323 = {1{`RANDOM}};
  pht_322 = _RAND_323[1:0];
  _RAND_324 = {1{`RANDOM}};
  pht_323 = _RAND_324[1:0];
  _RAND_325 = {1{`RANDOM}};
  pht_324 = _RAND_325[1:0];
  _RAND_326 = {1{`RANDOM}};
  pht_325 = _RAND_326[1:0];
  _RAND_327 = {1{`RANDOM}};
  pht_326 = _RAND_327[1:0];
  _RAND_328 = {1{`RANDOM}};
  pht_327 = _RAND_328[1:0];
  _RAND_329 = {1{`RANDOM}};
  pht_328 = _RAND_329[1:0];
  _RAND_330 = {1{`RANDOM}};
  pht_329 = _RAND_330[1:0];
  _RAND_331 = {1{`RANDOM}};
  pht_330 = _RAND_331[1:0];
  _RAND_332 = {1{`RANDOM}};
  pht_331 = _RAND_332[1:0];
  _RAND_333 = {1{`RANDOM}};
  pht_332 = _RAND_333[1:0];
  _RAND_334 = {1{`RANDOM}};
  pht_333 = _RAND_334[1:0];
  _RAND_335 = {1{`RANDOM}};
  pht_334 = _RAND_335[1:0];
  _RAND_336 = {1{`RANDOM}};
  pht_335 = _RAND_336[1:0];
  _RAND_337 = {1{`RANDOM}};
  pht_336 = _RAND_337[1:0];
  _RAND_338 = {1{`RANDOM}};
  pht_337 = _RAND_338[1:0];
  _RAND_339 = {1{`RANDOM}};
  pht_338 = _RAND_339[1:0];
  _RAND_340 = {1{`RANDOM}};
  pht_339 = _RAND_340[1:0];
  _RAND_341 = {1{`RANDOM}};
  pht_340 = _RAND_341[1:0];
  _RAND_342 = {1{`RANDOM}};
  pht_341 = _RAND_342[1:0];
  _RAND_343 = {1{`RANDOM}};
  pht_342 = _RAND_343[1:0];
  _RAND_344 = {1{`RANDOM}};
  pht_343 = _RAND_344[1:0];
  _RAND_345 = {1{`RANDOM}};
  pht_344 = _RAND_345[1:0];
  _RAND_346 = {1{`RANDOM}};
  pht_345 = _RAND_346[1:0];
  _RAND_347 = {1{`RANDOM}};
  pht_346 = _RAND_347[1:0];
  _RAND_348 = {1{`RANDOM}};
  pht_347 = _RAND_348[1:0];
  _RAND_349 = {1{`RANDOM}};
  pht_348 = _RAND_349[1:0];
  _RAND_350 = {1{`RANDOM}};
  pht_349 = _RAND_350[1:0];
  _RAND_351 = {1{`RANDOM}};
  pht_350 = _RAND_351[1:0];
  _RAND_352 = {1{`RANDOM}};
  pht_351 = _RAND_352[1:0];
  _RAND_353 = {1{`RANDOM}};
  pht_352 = _RAND_353[1:0];
  _RAND_354 = {1{`RANDOM}};
  pht_353 = _RAND_354[1:0];
  _RAND_355 = {1{`RANDOM}};
  pht_354 = _RAND_355[1:0];
  _RAND_356 = {1{`RANDOM}};
  pht_355 = _RAND_356[1:0];
  _RAND_357 = {1{`RANDOM}};
  pht_356 = _RAND_357[1:0];
  _RAND_358 = {1{`RANDOM}};
  pht_357 = _RAND_358[1:0];
  _RAND_359 = {1{`RANDOM}};
  pht_358 = _RAND_359[1:0];
  _RAND_360 = {1{`RANDOM}};
  pht_359 = _RAND_360[1:0];
  _RAND_361 = {1{`RANDOM}};
  pht_360 = _RAND_361[1:0];
  _RAND_362 = {1{`RANDOM}};
  pht_361 = _RAND_362[1:0];
  _RAND_363 = {1{`RANDOM}};
  pht_362 = _RAND_363[1:0];
  _RAND_364 = {1{`RANDOM}};
  pht_363 = _RAND_364[1:0];
  _RAND_365 = {1{`RANDOM}};
  pht_364 = _RAND_365[1:0];
  _RAND_366 = {1{`RANDOM}};
  pht_365 = _RAND_366[1:0];
  _RAND_367 = {1{`RANDOM}};
  pht_366 = _RAND_367[1:0];
  _RAND_368 = {1{`RANDOM}};
  pht_367 = _RAND_368[1:0];
  _RAND_369 = {1{`RANDOM}};
  pht_368 = _RAND_369[1:0];
  _RAND_370 = {1{`RANDOM}};
  pht_369 = _RAND_370[1:0];
  _RAND_371 = {1{`RANDOM}};
  pht_370 = _RAND_371[1:0];
  _RAND_372 = {1{`RANDOM}};
  pht_371 = _RAND_372[1:0];
  _RAND_373 = {1{`RANDOM}};
  pht_372 = _RAND_373[1:0];
  _RAND_374 = {1{`RANDOM}};
  pht_373 = _RAND_374[1:0];
  _RAND_375 = {1{`RANDOM}};
  pht_374 = _RAND_375[1:0];
  _RAND_376 = {1{`RANDOM}};
  pht_375 = _RAND_376[1:0];
  _RAND_377 = {1{`RANDOM}};
  pht_376 = _RAND_377[1:0];
  _RAND_378 = {1{`RANDOM}};
  pht_377 = _RAND_378[1:0];
  _RAND_379 = {1{`RANDOM}};
  pht_378 = _RAND_379[1:0];
  _RAND_380 = {1{`RANDOM}};
  pht_379 = _RAND_380[1:0];
  _RAND_381 = {1{`RANDOM}};
  pht_380 = _RAND_381[1:0];
  _RAND_382 = {1{`RANDOM}};
  pht_381 = _RAND_382[1:0];
  _RAND_383 = {1{`RANDOM}};
  pht_382 = _RAND_383[1:0];
  _RAND_384 = {1{`RANDOM}};
  pht_383 = _RAND_384[1:0];
  _RAND_385 = {1{`RANDOM}};
  pht_384 = _RAND_385[1:0];
  _RAND_386 = {1{`RANDOM}};
  pht_385 = _RAND_386[1:0];
  _RAND_387 = {1{`RANDOM}};
  pht_386 = _RAND_387[1:0];
  _RAND_388 = {1{`RANDOM}};
  pht_387 = _RAND_388[1:0];
  _RAND_389 = {1{`RANDOM}};
  pht_388 = _RAND_389[1:0];
  _RAND_390 = {1{`RANDOM}};
  pht_389 = _RAND_390[1:0];
  _RAND_391 = {1{`RANDOM}};
  pht_390 = _RAND_391[1:0];
  _RAND_392 = {1{`RANDOM}};
  pht_391 = _RAND_392[1:0];
  _RAND_393 = {1{`RANDOM}};
  pht_392 = _RAND_393[1:0];
  _RAND_394 = {1{`RANDOM}};
  pht_393 = _RAND_394[1:0];
  _RAND_395 = {1{`RANDOM}};
  pht_394 = _RAND_395[1:0];
  _RAND_396 = {1{`RANDOM}};
  pht_395 = _RAND_396[1:0];
  _RAND_397 = {1{`RANDOM}};
  pht_396 = _RAND_397[1:0];
  _RAND_398 = {1{`RANDOM}};
  pht_397 = _RAND_398[1:0];
  _RAND_399 = {1{`RANDOM}};
  pht_398 = _RAND_399[1:0];
  _RAND_400 = {1{`RANDOM}};
  pht_399 = _RAND_400[1:0];
  _RAND_401 = {1{`RANDOM}};
  pht_400 = _RAND_401[1:0];
  _RAND_402 = {1{`RANDOM}};
  pht_401 = _RAND_402[1:0];
  _RAND_403 = {1{`RANDOM}};
  pht_402 = _RAND_403[1:0];
  _RAND_404 = {1{`RANDOM}};
  pht_403 = _RAND_404[1:0];
  _RAND_405 = {1{`RANDOM}};
  pht_404 = _RAND_405[1:0];
  _RAND_406 = {1{`RANDOM}};
  pht_405 = _RAND_406[1:0];
  _RAND_407 = {1{`RANDOM}};
  pht_406 = _RAND_407[1:0];
  _RAND_408 = {1{`RANDOM}};
  pht_407 = _RAND_408[1:0];
  _RAND_409 = {1{`RANDOM}};
  pht_408 = _RAND_409[1:0];
  _RAND_410 = {1{`RANDOM}};
  pht_409 = _RAND_410[1:0];
  _RAND_411 = {1{`RANDOM}};
  pht_410 = _RAND_411[1:0];
  _RAND_412 = {1{`RANDOM}};
  pht_411 = _RAND_412[1:0];
  _RAND_413 = {1{`RANDOM}};
  pht_412 = _RAND_413[1:0];
  _RAND_414 = {1{`RANDOM}};
  pht_413 = _RAND_414[1:0];
  _RAND_415 = {1{`RANDOM}};
  pht_414 = _RAND_415[1:0];
  _RAND_416 = {1{`RANDOM}};
  pht_415 = _RAND_416[1:0];
  _RAND_417 = {1{`RANDOM}};
  pht_416 = _RAND_417[1:0];
  _RAND_418 = {1{`RANDOM}};
  pht_417 = _RAND_418[1:0];
  _RAND_419 = {1{`RANDOM}};
  pht_418 = _RAND_419[1:0];
  _RAND_420 = {1{`RANDOM}};
  pht_419 = _RAND_420[1:0];
  _RAND_421 = {1{`RANDOM}};
  pht_420 = _RAND_421[1:0];
  _RAND_422 = {1{`RANDOM}};
  pht_421 = _RAND_422[1:0];
  _RAND_423 = {1{`RANDOM}};
  pht_422 = _RAND_423[1:0];
  _RAND_424 = {1{`RANDOM}};
  pht_423 = _RAND_424[1:0];
  _RAND_425 = {1{`RANDOM}};
  pht_424 = _RAND_425[1:0];
  _RAND_426 = {1{`RANDOM}};
  pht_425 = _RAND_426[1:0];
  _RAND_427 = {1{`RANDOM}};
  pht_426 = _RAND_427[1:0];
  _RAND_428 = {1{`RANDOM}};
  pht_427 = _RAND_428[1:0];
  _RAND_429 = {1{`RANDOM}};
  pht_428 = _RAND_429[1:0];
  _RAND_430 = {1{`RANDOM}};
  pht_429 = _RAND_430[1:0];
  _RAND_431 = {1{`RANDOM}};
  pht_430 = _RAND_431[1:0];
  _RAND_432 = {1{`RANDOM}};
  pht_431 = _RAND_432[1:0];
  _RAND_433 = {1{`RANDOM}};
  pht_432 = _RAND_433[1:0];
  _RAND_434 = {1{`RANDOM}};
  pht_433 = _RAND_434[1:0];
  _RAND_435 = {1{`RANDOM}};
  pht_434 = _RAND_435[1:0];
  _RAND_436 = {1{`RANDOM}};
  pht_435 = _RAND_436[1:0];
  _RAND_437 = {1{`RANDOM}};
  pht_436 = _RAND_437[1:0];
  _RAND_438 = {1{`RANDOM}};
  pht_437 = _RAND_438[1:0];
  _RAND_439 = {1{`RANDOM}};
  pht_438 = _RAND_439[1:0];
  _RAND_440 = {1{`RANDOM}};
  pht_439 = _RAND_440[1:0];
  _RAND_441 = {1{`RANDOM}};
  pht_440 = _RAND_441[1:0];
  _RAND_442 = {1{`RANDOM}};
  pht_441 = _RAND_442[1:0];
  _RAND_443 = {1{`RANDOM}};
  pht_442 = _RAND_443[1:0];
  _RAND_444 = {1{`RANDOM}};
  pht_443 = _RAND_444[1:0];
  _RAND_445 = {1{`RANDOM}};
  pht_444 = _RAND_445[1:0];
  _RAND_446 = {1{`RANDOM}};
  pht_445 = _RAND_446[1:0];
  _RAND_447 = {1{`RANDOM}};
  pht_446 = _RAND_447[1:0];
  _RAND_448 = {1{`RANDOM}};
  pht_447 = _RAND_448[1:0];
  _RAND_449 = {1{`RANDOM}};
  pht_448 = _RAND_449[1:0];
  _RAND_450 = {1{`RANDOM}};
  pht_449 = _RAND_450[1:0];
  _RAND_451 = {1{`RANDOM}};
  pht_450 = _RAND_451[1:0];
  _RAND_452 = {1{`RANDOM}};
  pht_451 = _RAND_452[1:0];
  _RAND_453 = {1{`RANDOM}};
  pht_452 = _RAND_453[1:0];
  _RAND_454 = {1{`RANDOM}};
  pht_453 = _RAND_454[1:0];
  _RAND_455 = {1{`RANDOM}};
  pht_454 = _RAND_455[1:0];
  _RAND_456 = {1{`RANDOM}};
  pht_455 = _RAND_456[1:0];
  _RAND_457 = {1{`RANDOM}};
  pht_456 = _RAND_457[1:0];
  _RAND_458 = {1{`RANDOM}};
  pht_457 = _RAND_458[1:0];
  _RAND_459 = {1{`RANDOM}};
  pht_458 = _RAND_459[1:0];
  _RAND_460 = {1{`RANDOM}};
  pht_459 = _RAND_460[1:0];
  _RAND_461 = {1{`RANDOM}};
  pht_460 = _RAND_461[1:0];
  _RAND_462 = {1{`RANDOM}};
  pht_461 = _RAND_462[1:0];
  _RAND_463 = {1{`RANDOM}};
  pht_462 = _RAND_463[1:0];
  _RAND_464 = {1{`RANDOM}};
  pht_463 = _RAND_464[1:0];
  _RAND_465 = {1{`RANDOM}};
  pht_464 = _RAND_465[1:0];
  _RAND_466 = {1{`RANDOM}};
  pht_465 = _RAND_466[1:0];
  _RAND_467 = {1{`RANDOM}};
  pht_466 = _RAND_467[1:0];
  _RAND_468 = {1{`RANDOM}};
  pht_467 = _RAND_468[1:0];
  _RAND_469 = {1{`RANDOM}};
  pht_468 = _RAND_469[1:0];
  _RAND_470 = {1{`RANDOM}};
  pht_469 = _RAND_470[1:0];
  _RAND_471 = {1{`RANDOM}};
  pht_470 = _RAND_471[1:0];
  _RAND_472 = {1{`RANDOM}};
  pht_471 = _RAND_472[1:0];
  _RAND_473 = {1{`RANDOM}};
  pht_472 = _RAND_473[1:0];
  _RAND_474 = {1{`RANDOM}};
  pht_473 = _RAND_474[1:0];
  _RAND_475 = {1{`RANDOM}};
  pht_474 = _RAND_475[1:0];
  _RAND_476 = {1{`RANDOM}};
  pht_475 = _RAND_476[1:0];
  _RAND_477 = {1{`RANDOM}};
  pht_476 = _RAND_477[1:0];
  _RAND_478 = {1{`RANDOM}};
  pht_477 = _RAND_478[1:0];
  _RAND_479 = {1{`RANDOM}};
  pht_478 = _RAND_479[1:0];
  _RAND_480 = {1{`RANDOM}};
  pht_479 = _RAND_480[1:0];
  _RAND_481 = {1{`RANDOM}};
  pht_480 = _RAND_481[1:0];
  _RAND_482 = {1{`RANDOM}};
  pht_481 = _RAND_482[1:0];
  _RAND_483 = {1{`RANDOM}};
  pht_482 = _RAND_483[1:0];
  _RAND_484 = {1{`RANDOM}};
  pht_483 = _RAND_484[1:0];
  _RAND_485 = {1{`RANDOM}};
  pht_484 = _RAND_485[1:0];
  _RAND_486 = {1{`RANDOM}};
  pht_485 = _RAND_486[1:0];
  _RAND_487 = {1{`RANDOM}};
  pht_486 = _RAND_487[1:0];
  _RAND_488 = {1{`RANDOM}};
  pht_487 = _RAND_488[1:0];
  _RAND_489 = {1{`RANDOM}};
  pht_488 = _RAND_489[1:0];
  _RAND_490 = {1{`RANDOM}};
  pht_489 = _RAND_490[1:0];
  _RAND_491 = {1{`RANDOM}};
  pht_490 = _RAND_491[1:0];
  _RAND_492 = {1{`RANDOM}};
  pht_491 = _RAND_492[1:0];
  _RAND_493 = {1{`RANDOM}};
  pht_492 = _RAND_493[1:0];
  _RAND_494 = {1{`RANDOM}};
  pht_493 = _RAND_494[1:0];
  _RAND_495 = {1{`RANDOM}};
  pht_494 = _RAND_495[1:0];
  _RAND_496 = {1{`RANDOM}};
  pht_495 = _RAND_496[1:0];
  _RAND_497 = {1{`RANDOM}};
  pht_496 = _RAND_497[1:0];
  _RAND_498 = {1{`RANDOM}};
  pht_497 = _RAND_498[1:0];
  _RAND_499 = {1{`RANDOM}};
  pht_498 = _RAND_499[1:0];
  _RAND_500 = {1{`RANDOM}};
  pht_499 = _RAND_500[1:0];
  _RAND_501 = {1{`RANDOM}};
  pht_500 = _RAND_501[1:0];
  _RAND_502 = {1{`RANDOM}};
  pht_501 = _RAND_502[1:0];
  _RAND_503 = {1{`RANDOM}};
  pht_502 = _RAND_503[1:0];
  _RAND_504 = {1{`RANDOM}};
  pht_503 = _RAND_504[1:0];
  _RAND_505 = {1{`RANDOM}};
  pht_504 = _RAND_505[1:0];
  _RAND_506 = {1{`RANDOM}};
  pht_505 = _RAND_506[1:0];
  _RAND_507 = {1{`RANDOM}};
  pht_506 = _RAND_507[1:0];
  _RAND_508 = {1{`RANDOM}};
  pht_507 = _RAND_508[1:0];
  _RAND_509 = {1{`RANDOM}};
  pht_508 = _RAND_509[1:0];
  _RAND_510 = {1{`RANDOM}};
  pht_509 = _RAND_510[1:0];
  _RAND_511 = {1{`RANDOM}};
  pht_510 = _RAND_511[1:0];
  _RAND_512 = {1{`RANDOM}};
  pht_511 = _RAND_512[1:0];
  _RAND_513 = {2{`RANDOM}};
  btb_0_tag = _RAND_513[36:0];
  _RAND_514 = {2{`RANDOM}};
  btb_0_target = _RAND_514[36:0];
  _RAND_515 = {1{`RANDOM}};
  btb_0_valid = _RAND_515[0:0];
  _RAND_516 = {2{`RANDOM}};
  btb_1_tag = _RAND_516[36:0];
  _RAND_517 = {2{`RANDOM}};
  btb_1_target = _RAND_517[36:0];
  _RAND_518 = {1{`RANDOM}};
  btb_1_valid = _RAND_518[0:0];
  _RAND_519 = {2{`RANDOM}};
  btb_2_tag = _RAND_519[36:0];
  _RAND_520 = {2{`RANDOM}};
  btb_2_target = _RAND_520[36:0];
  _RAND_521 = {1{`RANDOM}};
  btb_2_valid = _RAND_521[0:0];
  _RAND_522 = {2{`RANDOM}};
  btb_3_tag = _RAND_522[36:0];
  _RAND_523 = {2{`RANDOM}};
  btb_3_target = _RAND_523[36:0];
  _RAND_524 = {1{`RANDOM}};
  btb_3_valid = _RAND_524[0:0];
  _RAND_525 = {2{`RANDOM}};
  btb_4_tag = _RAND_525[36:0];
  _RAND_526 = {2{`RANDOM}};
  btb_4_target = _RAND_526[36:0];
  _RAND_527 = {1{`RANDOM}};
  btb_4_valid = _RAND_527[0:0];
  _RAND_528 = {2{`RANDOM}};
  btb_5_tag = _RAND_528[36:0];
  _RAND_529 = {2{`RANDOM}};
  btb_5_target = _RAND_529[36:0];
  _RAND_530 = {1{`RANDOM}};
  btb_5_valid = _RAND_530[0:0];
  _RAND_531 = {2{`RANDOM}};
  btb_6_tag = _RAND_531[36:0];
  _RAND_532 = {2{`RANDOM}};
  btb_6_target = _RAND_532[36:0];
  _RAND_533 = {1{`RANDOM}};
  btb_6_valid = _RAND_533[0:0];
  _RAND_534 = {2{`RANDOM}};
  btb_7_tag = _RAND_534[36:0];
  _RAND_535 = {2{`RANDOM}};
  btb_7_target = _RAND_535[36:0];
  _RAND_536 = {1{`RANDOM}};
  btb_7_valid = _RAND_536[0:0];
  _RAND_537 = {2{`RANDOM}};
  btb_8_tag = _RAND_537[36:0];
  _RAND_538 = {2{`RANDOM}};
  btb_8_target = _RAND_538[36:0];
  _RAND_539 = {1{`RANDOM}};
  btb_8_valid = _RAND_539[0:0];
  _RAND_540 = {2{`RANDOM}};
  btb_9_tag = _RAND_540[36:0];
  _RAND_541 = {2{`RANDOM}};
  btb_9_target = _RAND_541[36:0];
  _RAND_542 = {1{`RANDOM}};
  btb_9_valid = _RAND_542[0:0];
  _RAND_543 = {2{`RANDOM}};
  btb_10_tag = _RAND_543[36:0];
  _RAND_544 = {2{`RANDOM}};
  btb_10_target = _RAND_544[36:0];
  _RAND_545 = {1{`RANDOM}};
  btb_10_valid = _RAND_545[0:0];
  _RAND_546 = {2{`RANDOM}};
  btb_11_tag = _RAND_546[36:0];
  _RAND_547 = {2{`RANDOM}};
  btb_11_target = _RAND_547[36:0];
  _RAND_548 = {1{`RANDOM}};
  btb_11_valid = _RAND_548[0:0];
  _RAND_549 = {2{`RANDOM}};
  btb_12_tag = _RAND_549[36:0];
  _RAND_550 = {2{`RANDOM}};
  btb_12_target = _RAND_550[36:0];
  _RAND_551 = {1{`RANDOM}};
  btb_12_valid = _RAND_551[0:0];
  _RAND_552 = {2{`RANDOM}};
  btb_13_tag = _RAND_552[36:0];
  _RAND_553 = {2{`RANDOM}};
  btb_13_target = _RAND_553[36:0];
  _RAND_554 = {1{`RANDOM}};
  btb_13_valid = _RAND_554[0:0];
  _RAND_555 = {2{`RANDOM}};
  btb_14_tag = _RAND_555[36:0];
  _RAND_556 = {2{`RANDOM}};
  btb_14_target = _RAND_556[36:0];
  _RAND_557 = {1{`RANDOM}};
  btb_14_valid = _RAND_557[0:0];
  _RAND_558 = {2{`RANDOM}};
  btb_15_tag = _RAND_558[36:0];
  _RAND_559 = {2{`RANDOM}};
  btb_15_target = _RAND_559[36:0];
  _RAND_560 = {1{`RANDOM}};
  btb_15_valid = _RAND_560[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IF0(
  input         clock,
  input         reset,
  input         io_jmp_packet_valid,
  input  [63:0] io_jmp_packet_target,
  input         io_jmp_packet_bp_update,
  input         io_jmp_packet_bp_taken,
  input  [63:0] io_jmp_packet_bp_pc,
  input         io_req_ready,
  output        io_req_valid,
  output [38:0] io_req_bits_addr,
  output [38:0] io_req_addr,
  output [63:0] io_bp_npc,
  input         io_stall_b
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  bpu_clock; // @[IFU.scala 21:21]
  wire  bpu_reset; // @[IFU.scala 21:21]
  wire [63:0] bpu_io_pc; // @[IFU.scala 21:21]
  wire [63:0] bpu_io_jmp_packet_target; // @[IFU.scala 21:21]
  wire  bpu_io_jmp_packet_bp_update; // @[IFU.scala 21:21]
  wire  bpu_io_jmp_packet_bp_taken; // @[IFU.scala 21:21]
  wire [63:0] bpu_io_jmp_packet_bp_pc; // @[IFU.scala 21:21]
  wire [63:0] bpu_io_out; // @[IFU.scala 21:21]
  wire  _pc_update_T = io_req_ready & io_req_valid; // @[Decoupled.scala 51:35]
  wire  pc_update = io_jmp_packet_valid | _pc_update_T; // @[IFU.scala 15:41]
  reg [63:0] pc; // @[Reg.scala 35:20]
  wire [63:0] jmp_target = {io_jmp_packet_target[63:2],2'h0}; // @[Cat.scala 33:92]
  wire [63:0] pc_next_raw = bpu_io_out; // @[IFU.scala 19:25 24:23]
  wire [63:0] _io_req_addr_T = io_jmp_packet_valid ? jmp_target : pc; // @[IFU.scala 33:26]
  BPU bpu ( // @[IFU.scala 21:21]
    .clock(bpu_clock),
    .reset(bpu_reset),
    .io_pc(bpu_io_pc),
    .io_jmp_packet_target(bpu_io_jmp_packet_target),
    .io_jmp_packet_bp_update(bpu_io_jmp_packet_bp_update),
    .io_jmp_packet_bp_taken(bpu_io_jmp_packet_bp_taken),
    .io_jmp_packet_bp_pc(bpu_io_jmp_packet_bp_pc),
    .io_out(bpu_io_out)
  );
  assign io_req_valid = io_stall_b; // @[IFU.scala 36:20]
  assign io_req_bits_addr = {io_req_addr[38:3],3'h0}; // @[Cat.scala 33:92]
  assign io_req_addr = _io_req_addr_T[38:0]; // @[IFU.scala 33:20]
  assign io_bp_npc = bpu_io_out; // @[IFU.scala 19:25 24:23]
  assign bpu_clock = clock;
  assign bpu_reset = reset;
  assign bpu_io_pc = io_jmp_packet_valid & _pc_update_T ? jmp_target : pc; // @[IFU.scala 22:29]
  assign bpu_io_jmp_packet_target = io_jmp_packet_target; // @[IFU.scala 23:23]
  assign bpu_io_jmp_packet_bp_update = io_jmp_packet_bp_update; // @[IFU.scala 23:23]
  assign bpu_io_jmp_packet_bp_taken = io_jmp_packet_bp_taken; // @[IFU.scala 23:23]
  assign bpu_io_jmp_packet_bp_pc = io_jmp_packet_bp_pc; // @[IFU.scala 23:23]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 35:20]
      pc <= 64'h10000; // @[Reg.scala 35:20]
    end else if (pc_update) begin // @[Reg.scala 36:18]
      if (io_jmp_packet_valid & ~_pc_update_T) begin // @[IFU.scala 31:20]
        pc <= jmp_target;
      end else begin
        pc <= pc_next_raw;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  pc = _RAND_0[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IF1(
  input   clock,
  input   reset,
  input   io_jmp_packet_valid,
  output  io_resp_ready,
  input   io_resp_valid,
  input   io_stall_b,
  output  io_out_valid,
  input   io_req_fire,
  input   io_pc_queue_empty
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[IFU.scala 51:50]
  wire  _jmp_r_T = io_resp_ready & io_resp_valid; // @[Decoupled.scala 51:35]
  wire  _jmp_r_T_6 = io_jmp_packet_valid & ~_jmp_r_T & state != 2'h2 & ~io_pc_queue_empty; // @[IFU.scala 54:64]
  reg  jmp_r; // @[Utils.scala 36:20]
  wire  _GEN_0 = _jmp_r_T_6 | jmp_r; // @[Utils.scala 41:19 36:20 41:23]
  wire  _state_to_wait_T_1 = ~jmp_r; // @[IFU.scala 58:81]
  wire  _state_to_wait_T_3 = ~io_jmp_packet_valid; // @[IFU.scala 58:91]
  wire [1:0] _state_T = io_jmp_packet_valid ? 2'h0 : 2'h1; // @[IFU.scala 68:21]
  wire [1:0] _GEN_4 = io_jmp_packet_valid ? 2'h0 : state; // @[IFU.scala 72:33 73:15 51:50]
  assign io_resp_ready = (io_stall_b | io_jmp_packet_valid) & state == 2'h1 | state == 2'h0; // @[IFU.scala 78:80]
  assign io_out_valid = _jmp_r_T & _state_to_wait_T_3 & _state_to_wait_T_1; // @[IFU.scala 81:56]
  always @(posedge clock) begin
    if (reset) begin // @[IFU.scala 51:50]
      state <= 2'h0; // @[IFU.scala 51:50]
    end else if (2'h0 == state) begin // @[IFU.scala 60:17]
      if (io_req_fire) begin // @[IFU.scala 62:25]
        state <= 2'h1; // @[IFU.scala 63:15]
      end
    end else if (2'h1 == state) begin // @[IFU.scala 60:17]
      if (_jmp_r_T) begin // @[IFU.scala 67:26]
        state <= _state_T; // @[IFU.scala 68:15]
      end
    end else if (2'h2 == state) begin // @[IFU.scala 60:17]
      state <= _GEN_4;
    end
    if (reset) begin // @[Utils.scala 36:20]
      jmp_r <= 1'h0; // @[Utils.scala 36:20]
    end else if (_jmp_r_T) begin // @[Utils.scala 42:18]
      jmp_r <= 1'h0; // @[Utils.scala 42:22]
    end else begin
      jmp_r <= _GEN_0;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  jmp_r = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [38:0] io_enq_bits,
  input         io_deq_ready,
  output        io_deq_valid,
  output [38:0] io_deq_bits,
  output        io_count
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [38:0] ram [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [38:0] ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [38:0] ram_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_MPORT_en; // @[Decoupled.scala 273:95]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 278:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  assign ram_io_deq_bits_MPORT_en = 1'h1;
  assign ram_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_MPORT_data = io_enq_bits;
  assign ram_MPORT_addr = 1'h0;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = io_deq_ready | empty; // @[Decoupled.scala 303:16 323:{24,39}]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits = ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_count = maybe_full; // @[Decoupled.scala 329:62]
  always @(posedge clock) begin
    if (ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram[initvar] = _RAND_0[38:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  maybe_full = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_1(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [63:0] io_enq_bits,
  input         io_deq_ready,
  output        io_deq_valid,
  output [63:0] io_deq_bits
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] ram [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [63:0] ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [63:0] ram_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_MPORT_en; // @[Decoupled.scala 273:95]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 278:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  assign ram_io_deq_bits_MPORT_en = 1'h1;
  assign ram_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_MPORT_data = io_enq_bits;
  assign ram_MPORT_addr = 1'h0;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = io_deq_ready | empty; // @[Decoupled.scala 303:16 323:{24,39}]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits = ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  always @(posedge clock) begin
    if (ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram[initvar] = _RAND_0[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  maybe_full = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IFU(
  input         clock,
  input         reset,
  input         io_jmp_packet_valid,
  input  [63:0] io_jmp_packet_target,
  input         io_jmp_packet_bp_update,
  input         io_jmp_packet_bp_taken,
  input  [63:0] io_jmp_packet_bp_pc,
  input         io_imem_req_ready,
  output        io_imem_req_valid,
  output [38:0] io_imem_req_bits_addr,
  output        io_imem_resp_ready,
  input         io_imem_resp_valid,
  input  [63:0] io_imem_resp_bits_rdata,
  input         io_imem_resp_bits_page_fault,
  input         io_imem_resp_bits_access_fault,
  output [63:0] io_out_pc,
  output [31:0] io_out_instr,
  output        io_out_valid,
  output        io_out_page_fault,
  output        io_out_access_fault,
  output [63:0] io_out_bp_npc,
  input         io_stall_b
);
  wire  if0_clock; // @[IFU.scala 96:19]
  wire  if0_reset; // @[IFU.scala 96:19]
  wire  if0_io_jmp_packet_valid; // @[IFU.scala 96:19]
  wire [63:0] if0_io_jmp_packet_target; // @[IFU.scala 96:19]
  wire  if0_io_jmp_packet_bp_update; // @[IFU.scala 96:19]
  wire  if0_io_jmp_packet_bp_taken; // @[IFU.scala 96:19]
  wire [63:0] if0_io_jmp_packet_bp_pc; // @[IFU.scala 96:19]
  wire  if0_io_req_ready; // @[IFU.scala 96:19]
  wire  if0_io_req_valid; // @[IFU.scala 96:19]
  wire [38:0] if0_io_req_bits_addr; // @[IFU.scala 96:19]
  wire [38:0] if0_io_req_addr; // @[IFU.scala 96:19]
  wire [63:0] if0_io_bp_npc; // @[IFU.scala 96:19]
  wire  if0_io_stall_b; // @[IFU.scala 96:19]
  wire  if1_clock; // @[IFU.scala 97:19]
  wire  if1_reset; // @[IFU.scala 97:19]
  wire  if1_io_jmp_packet_valid; // @[IFU.scala 97:19]
  wire  if1_io_resp_ready; // @[IFU.scala 97:19]
  wire  if1_io_resp_valid; // @[IFU.scala 97:19]
  wire  if1_io_stall_b; // @[IFU.scala 97:19]
  wire  if1_io_out_valid; // @[IFU.scala 97:19]
  wire  if1_io_req_fire; // @[IFU.scala 97:19]
  wire  if1_io_pc_queue_empty; // @[IFU.scala 97:19]
  wire  pc_queue_clock; // @[IFU.scala 99:28]
  wire  pc_queue_reset; // @[IFU.scala 99:28]
  wire  pc_queue_io_enq_ready; // @[IFU.scala 99:28]
  wire  pc_queue_io_enq_valid; // @[IFU.scala 99:28]
  wire [38:0] pc_queue_io_enq_bits; // @[IFU.scala 99:28]
  wire  pc_queue_io_deq_ready; // @[IFU.scala 99:28]
  wire  pc_queue_io_deq_valid; // @[IFU.scala 99:28]
  wire [38:0] pc_queue_io_deq_bits; // @[IFU.scala 99:28]
  wire  pc_queue_io_count; // @[IFU.scala 99:28]
  wire  bp_npc_queue_clock; // @[IFU.scala 100:28]
  wire  bp_npc_queue_reset; // @[IFU.scala 100:28]
  wire  bp_npc_queue_io_enq_ready; // @[IFU.scala 100:28]
  wire  bp_npc_queue_io_enq_valid; // @[IFU.scala 100:28]
  wire [63:0] bp_npc_queue_io_enq_bits; // @[IFU.scala 100:28]
  wire  bp_npc_queue_io_deq_ready; // @[IFU.scala 100:28]
  wire  bp_npc_queue_io_deq_valid; // @[IFU.scala 100:28]
  wire [63:0] bp_npc_queue_io_deq_bits; // @[IFU.scala 100:28]
  wire [24:0] _io_out_pc_T_2 = pc_queue_io_deq_bits[38] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 77:12]
  IF0 if0 ( // @[IFU.scala 96:19]
    .clock(if0_clock),
    .reset(if0_reset),
    .io_jmp_packet_valid(if0_io_jmp_packet_valid),
    .io_jmp_packet_target(if0_io_jmp_packet_target),
    .io_jmp_packet_bp_update(if0_io_jmp_packet_bp_update),
    .io_jmp_packet_bp_taken(if0_io_jmp_packet_bp_taken),
    .io_jmp_packet_bp_pc(if0_io_jmp_packet_bp_pc),
    .io_req_ready(if0_io_req_ready),
    .io_req_valid(if0_io_req_valid),
    .io_req_bits_addr(if0_io_req_bits_addr),
    .io_req_addr(if0_io_req_addr),
    .io_bp_npc(if0_io_bp_npc),
    .io_stall_b(if0_io_stall_b)
  );
  IF1 if1 ( // @[IFU.scala 97:19]
    .clock(if1_clock),
    .reset(if1_reset),
    .io_jmp_packet_valid(if1_io_jmp_packet_valid),
    .io_resp_ready(if1_io_resp_ready),
    .io_resp_valid(if1_io_resp_valid),
    .io_stall_b(if1_io_stall_b),
    .io_out_valid(if1_io_out_valid),
    .io_req_fire(if1_io_req_fire),
    .io_pc_queue_empty(if1_io_pc_queue_empty)
  );
  Queue pc_queue ( // @[IFU.scala 99:28]
    .clock(pc_queue_clock),
    .reset(pc_queue_reset),
    .io_enq_ready(pc_queue_io_enq_ready),
    .io_enq_valid(pc_queue_io_enq_valid),
    .io_enq_bits(pc_queue_io_enq_bits),
    .io_deq_ready(pc_queue_io_deq_ready),
    .io_deq_valid(pc_queue_io_deq_valid),
    .io_deq_bits(pc_queue_io_deq_bits),
    .io_count(pc_queue_io_count)
  );
  Queue_1 bp_npc_queue ( // @[IFU.scala 100:28]
    .clock(bp_npc_queue_clock),
    .reset(bp_npc_queue_reset),
    .io_enq_ready(bp_npc_queue_io_enq_ready),
    .io_enq_valid(bp_npc_queue_io_enq_valid),
    .io_enq_bits(bp_npc_queue_io_enq_bits),
    .io_deq_ready(bp_npc_queue_io_deq_ready),
    .io_deq_valid(bp_npc_queue_io_deq_valid),
    .io_deq_bits(bp_npc_queue_io_deq_bits)
  );
  assign io_imem_req_valid = if0_io_req_valid; // @[IFU.scala 103:21]
  assign io_imem_req_bits_addr = if0_io_req_bits_addr; // @[IFU.scala 103:21]
  assign io_imem_resp_ready = if1_io_resp_ready; // @[IFU.scala 107:25]
  assign io_out_pc = {_io_out_pc_T_2,pc_queue_io_deq_bits}; // @[Cat.scala 33:92]
  assign io_out_instr = io_out_pc[2] ? io_imem_resp_bits_rdata[63:32] : io_imem_resp_bits_rdata[31:0]; // @[IFU.scala 122:29]
  assign io_out_valid = if1_io_out_valid; // @[IFU.scala 120:23]
  assign io_out_page_fault = io_imem_resp_bits_page_fault; // @[IFU.scala 123:23]
  assign io_out_access_fault = io_imem_resp_bits_access_fault; // @[IFU.scala 124:23]
  assign io_out_bp_npc = bp_npc_queue_io_deq_bits; // @[IFU.scala 125:23]
  assign if0_clock = clock;
  assign if0_reset = reset;
  assign if0_io_jmp_packet_valid = io_jmp_packet_valid; // @[IFU.scala 102:21]
  assign if0_io_jmp_packet_target = io_jmp_packet_target; // @[IFU.scala 102:21]
  assign if0_io_jmp_packet_bp_update = io_jmp_packet_bp_update; // @[IFU.scala 102:21]
  assign if0_io_jmp_packet_bp_taken = io_jmp_packet_bp_taken; // @[IFU.scala 102:21]
  assign if0_io_jmp_packet_bp_pc = io_jmp_packet_bp_pc; // @[IFU.scala 102:21]
  assign if0_io_req_ready = io_imem_req_ready; // @[IFU.scala 103:21]
  assign if0_io_stall_b = pc_queue_io_enq_ready & io_stall_b; // @[IFU.scala 104:46]
  assign if1_clock = clock;
  assign if1_reset = reset;
  assign if1_io_jmp_packet_valid = io_jmp_packet_valid; // @[IFU.scala 106:25]
  assign if1_io_resp_valid = io_imem_resp_valid; // @[IFU.scala 107:25]
  assign if1_io_stall_b = io_stall_b; // @[IFU.scala 108:25]
  assign if1_io_req_fire = io_imem_req_ready & io_imem_req_valid; // @[Decoupled.scala 51:35]
  assign if1_io_pc_queue_empty = ~pc_queue_io_count; // @[IFU.scala 110:47]
  assign pc_queue_clock = clock;
  assign pc_queue_reset = reset;
  assign pc_queue_io_enq_valid = io_imem_req_ready & io_imem_req_valid; // @[Decoupled.scala 51:35]
  assign pc_queue_io_enq_bits = if0_io_req_addr; // @[IFU.scala 112:25]
  assign pc_queue_io_deq_ready = io_imem_resp_ready & io_imem_resp_valid; // @[Decoupled.scala 51:35]
  assign bp_npc_queue_clock = clock;
  assign bp_npc_queue_reset = reset;
  assign bp_npc_queue_io_enq_valid = io_imem_req_ready & io_imem_req_valid; // @[Decoupled.scala 51:35]
  assign bp_npc_queue_io_enq_bits = if0_io_bp_npc; // @[IFU.scala 116:29]
  assign bp_npc_queue_io_deq_ready = io_imem_resp_ready & io_imem_resp_valid; // @[Decoupled.scala 51:35]
endmodule
module MaxPeriodFibonacciLFSR_1(
  input   clock,
  input   reset,
  output  io_out_0,
  output  io_out_1,
  output  io_out_2,
  output  io_out_3,
  output  io_out_4
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg  state_0; // @[PRNG.scala 55:49]
  reg  state_1; // @[PRNG.scala 55:49]
  reg  state_2; // @[PRNG.scala 55:49]
  reg  state_3; // @[PRNG.scala 55:49]
  reg  state_4; // @[PRNG.scala 55:49]
  wire  _T = state_4 ^ state_2; // @[LFSR.scala 15:41]
  assign io_out_0 = state_0; // @[PRNG.scala 78:10]
  assign io_out_1 = state_1; // @[PRNG.scala 78:10]
  assign io_out_2 = state_2; // @[PRNG.scala 78:10]
  assign io_out_3 = state_3; // @[PRNG.scala 78:10]
  assign io_out_4 = state_4; // @[PRNG.scala 78:10]
  always @(posedge clock) begin
    state_0 <= reset | _T; // @[PRNG.scala 55:{49,49}]
    if (reset) begin // @[PRNG.scala 55:49]
      state_1 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_1 <= state_0;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_2 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_2 <= state_1;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_3 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_3 <= state_2;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_4 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_4 <= state_3;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  state_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  state_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  state_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  state_4 = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLB(
  input         clock,
  input         reset,
  input         io_sfence_vma,
  input  [8:0]  io_vaddr_vpn2,
  input  [8:0]  io_vaddr_vpn1,
  input  [8:0]  io_vaddr_vpn0,
  output [1:0]  io_rpte_ppn2,
  output [8:0]  io_rpte_ppn1,
  output [8:0]  io_rpte_ppn0,
  output        io_rpte_flag_d,
  output        io_rpte_flag_a,
  output        io_rpte_flag_u,
  output        io_rpte_flag_x,
  output        io_rpte_flag_w,
  output        io_rpte_flag_r,
  output        io_rpte_flag_v,
  output [1:0]  io_rlevel,
  output        io_hit,
  input         io_wen,
  input  [8:0]  io_wvaddr_vpn2,
  input  [8:0]  io_wvaddr_vpn1,
  input  [8:0]  io_wvaddr_vpn0,
  input  [1:0]  io_wpte_ppn2,
  input  [8:0]  io_wpte_ppn1,
  input  [8:0]  io_wpte_ppn0,
  input         io_wpte_flag_d,
  input         io_wpte_flag_a,
  input         io_wpte_flag_g,
  input         io_wpte_flag_u,
  input         io_wpte_flag_x,
  input         io_wpte_flag_w,
  input         io_wpte_flag_r,
  input         io_wpte_flag_v,
  input  [1:0]  io_wlevel,
  input  [15:0] io_satp_asid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
`endif // RANDOMIZE_REG_INIT
  wire  replace_idx_prng_clock; // @[PRNG.scala 91:22]
  wire  replace_idx_prng_reset; // @[PRNG.scala 91:22]
  wire  replace_idx_prng_io_out_0; // @[PRNG.scala 91:22]
  wire  replace_idx_prng_io_out_1; // @[PRNG.scala 91:22]
  wire  replace_idx_prng_io_out_2; // @[PRNG.scala 91:22]
  wire  replace_idx_prng_io_out_3; // @[PRNG.scala 91:22]
  wire  replace_idx_prng_io_out_4; // @[PRNG.scala 91:22]
  wire  _T_2 = ~reset; // @[TLB.scala 48:9]
  wire [4:0] replace_idx = {replace_idx_prng_io_out_4,replace_idx_prng_io_out_3,replace_idx_prng_io_out_2,
    replace_idx_prng_io_out_1,replace_idx_prng_io_out_0}; // @[PRNG.scala 95:17]
  reg  array4kb_0_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_0_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_0_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_0_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_0_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_0_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_0_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_0_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_0_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_0_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_0_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_0_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_0_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_0_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_0_asid; // @[TLB.scala 64:31]
  reg  array4kb_1_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_1_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_1_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_1_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_1_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_1_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_1_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_1_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_1_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_1_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_1_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_1_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_1_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_1_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_1_asid; // @[TLB.scala 64:31]
  reg  array4kb_2_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_2_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_2_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_2_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_2_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_2_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_2_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_2_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_2_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_2_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_2_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_2_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_2_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_2_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_2_asid; // @[TLB.scala 64:31]
  reg  array4kb_3_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_3_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_3_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_3_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_3_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_3_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_3_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_3_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_3_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_3_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_3_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_3_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_3_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_3_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_3_asid; // @[TLB.scala 64:31]
  reg  array4kb_4_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_4_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_4_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_4_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_4_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_4_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_4_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_4_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_4_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_4_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_4_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_4_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_4_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_4_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_4_asid; // @[TLB.scala 64:31]
  reg  array4kb_5_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_5_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_5_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_5_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_5_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_5_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_5_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_5_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_5_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_5_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_5_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_5_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_5_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_5_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_5_asid; // @[TLB.scala 64:31]
  reg  array4kb_6_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_6_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_6_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_6_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_6_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_6_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_6_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_6_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_6_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_6_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_6_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_6_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_6_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_6_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_6_asid; // @[TLB.scala 64:31]
  reg  array4kb_7_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_7_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_7_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_7_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_7_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_7_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_7_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_7_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_7_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_7_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_7_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_7_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_7_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_7_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_7_asid; // @[TLB.scala 64:31]
  reg  array4kb_8_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_8_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_8_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_8_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_8_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_8_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_8_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_8_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_8_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_8_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_8_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_8_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_8_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_8_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_8_asid; // @[TLB.scala 64:31]
  reg  array4kb_9_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_9_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_9_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_9_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_9_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_9_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_9_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_9_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_9_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_9_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_9_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_9_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_9_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_9_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_9_asid; // @[TLB.scala 64:31]
  reg  array4kb_10_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_10_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_10_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_10_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_10_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_10_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_10_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_10_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_10_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_10_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_10_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_10_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_10_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_10_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_10_asid; // @[TLB.scala 64:31]
  reg  array4kb_11_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_11_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_11_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_11_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_11_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_11_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_11_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_11_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_11_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_11_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_11_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_11_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_11_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_11_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_11_asid; // @[TLB.scala 64:31]
  reg  array4kb_12_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_12_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_12_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_12_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_12_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_12_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_12_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_12_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_12_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_12_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_12_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_12_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_12_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_12_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_12_asid; // @[TLB.scala 64:31]
  reg  array4kb_13_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_13_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_13_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_13_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_13_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_13_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_13_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_13_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_13_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_13_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_13_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_13_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_13_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_13_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_13_asid; // @[TLB.scala 64:31]
  reg  array4kb_14_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_14_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_14_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_14_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_14_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_14_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_14_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_14_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_14_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_14_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_14_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_14_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_14_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_14_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_14_asid; // @[TLB.scala 64:31]
  reg  array4kb_15_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_15_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_15_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_15_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_15_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_15_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_15_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_15_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_15_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_15_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_15_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_15_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_15_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_15_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_15_asid; // @[TLB.scala 64:31]
  reg  array4kb_16_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_16_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_16_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_16_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_16_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_16_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_16_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_16_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_16_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_16_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_16_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_16_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_16_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_16_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_16_asid; // @[TLB.scala 64:31]
  reg  array4kb_17_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_17_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_17_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_17_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_17_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_17_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_17_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_17_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_17_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_17_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_17_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_17_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_17_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_17_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_17_asid; // @[TLB.scala 64:31]
  reg  array4kb_18_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_18_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_18_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_18_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_18_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_18_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_18_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_18_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_18_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_18_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_18_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_18_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_18_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_18_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_18_asid; // @[TLB.scala 64:31]
  reg  array4kb_19_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_19_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_19_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_19_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_19_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_19_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_19_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_19_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_19_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_19_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_19_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_19_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_19_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_19_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_19_asid; // @[TLB.scala 64:31]
  reg  array4kb_20_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_20_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_20_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_20_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_20_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_20_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_20_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_20_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_20_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_20_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_20_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_20_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_20_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_20_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_20_asid; // @[TLB.scala 64:31]
  reg  array4kb_21_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_21_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_21_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_21_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_21_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_21_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_21_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_21_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_21_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_21_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_21_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_21_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_21_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_21_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_21_asid; // @[TLB.scala 64:31]
  reg  array4kb_22_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_22_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_22_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_22_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_22_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_22_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_22_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_22_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_22_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_22_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_22_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_22_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_22_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_22_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_22_asid; // @[TLB.scala 64:31]
  reg  array4kb_23_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_23_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_23_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_23_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_23_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_23_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_23_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_23_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_23_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_23_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_23_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_23_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_23_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_23_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_23_asid; // @[TLB.scala 64:31]
  reg  array4kb_24_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_24_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_24_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_24_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_24_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_24_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_24_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_24_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_24_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_24_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_24_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_24_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_24_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_24_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_24_asid; // @[TLB.scala 64:31]
  reg  array4kb_25_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_25_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_25_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_25_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_25_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_25_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_25_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_25_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_25_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_25_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_25_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_25_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_25_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_25_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_25_asid; // @[TLB.scala 64:31]
  reg  array4kb_26_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_26_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_26_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_26_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_26_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_26_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_26_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_26_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_26_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_26_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_26_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_26_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_26_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_26_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_26_asid; // @[TLB.scala 64:31]
  reg  array4kb_27_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_27_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_27_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_27_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_27_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_27_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_27_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_27_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_27_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_27_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_27_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_27_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_27_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_27_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_27_asid; // @[TLB.scala 64:31]
  reg  array4kb_28_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_28_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_28_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_28_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_28_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_28_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_28_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_28_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_28_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_28_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_28_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_28_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_28_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_28_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_28_asid; // @[TLB.scala 64:31]
  reg  array4kb_29_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_29_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_29_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_29_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_29_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_29_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_29_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_29_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_29_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_29_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_29_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_29_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_29_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_29_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_29_asid; // @[TLB.scala 64:31]
  reg  array4kb_30_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_30_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_30_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_30_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_30_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_30_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_30_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_30_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_30_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_30_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_30_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_30_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_30_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_30_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_30_asid; // @[TLB.scala 64:31]
  reg  array4kb_31_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_31_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_31_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_31_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_31_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_31_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_31_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_31_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_31_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_31_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_31_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_31_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_31_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_31_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_31_asid; // @[TLB.scala 64:31]
  reg  array4kb_valid_0; // @[TLB.scala 65:31]
  reg  array4kb_valid_1; // @[TLB.scala 65:31]
  reg  array4kb_valid_2; // @[TLB.scala 65:31]
  reg  array4kb_valid_3; // @[TLB.scala 65:31]
  reg  array4kb_valid_4; // @[TLB.scala 65:31]
  reg  array4kb_valid_5; // @[TLB.scala 65:31]
  reg  array4kb_valid_6; // @[TLB.scala 65:31]
  reg  array4kb_valid_7; // @[TLB.scala 65:31]
  reg  array4kb_valid_8; // @[TLB.scala 65:31]
  reg  array4kb_valid_9; // @[TLB.scala 65:31]
  reg  array4kb_valid_10; // @[TLB.scala 65:31]
  reg  array4kb_valid_11; // @[TLB.scala 65:31]
  reg  array4kb_valid_12; // @[TLB.scala 65:31]
  reg  array4kb_valid_13; // @[TLB.scala 65:31]
  reg  array4kb_valid_14; // @[TLB.scala 65:31]
  reg  array4kb_valid_15; // @[TLB.scala 65:31]
  reg  array4kb_valid_16; // @[TLB.scala 65:31]
  reg  array4kb_valid_17; // @[TLB.scala 65:31]
  reg  array4kb_valid_18; // @[TLB.scala 65:31]
  reg  array4kb_valid_19; // @[TLB.scala 65:31]
  reg  array4kb_valid_20; // @[TLB.scala 65:31]
  reg  array4kb_valid_21; // @[TLB.scala 65:31]
  reg  array4kb_valid_22; // @[TLB.scala 65:31]
  reg  array4kb_valid_23; // @[TLB.scala 65:31]
  reg  array4kb_valid_24; // @[TLB.scala 65:31]
  reg  array4kb_valid_25; // @[TLB.scala 65:31]
  reg  array4kb_valid_26; // @[TLB.scala 65:31]
  reg  array4kb_valid_27; // @[TLB.scala 65:31]
  reg  array4kb_valid_28; // @[TLB.scala 65:31]
  reg  array4kb_valid_29; // @[TLB.scala 65:31]
  reg  array4kb_valid_30; // @[TLB.scala 65:31]
  reg  array4kb_valid_31; // @[TLB.scala 65:31]
  wire [26:0] _T_8 = {array4kb_0_vpn2,array4kb_0_vpn1,array4kb_0_vpn0}; // @[Cat.scala 33:92]
  wire [17:0] hi_1 = {io_vaddr_vpn2,io_vaddr_vpn1}; // @[Cat.scala 33:92]
  wire [26:0] _T_9 = {io_vaddr_vpn2,io_vaddr_vpn1,io_vaddr_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_0 = array4kb_valid_0 & _T_8 == _T_9 & (array4kb_0_asid == io_satp_asid | array4kb_0_flag_g); // @[TLB.scala 71:71 72:22 68:35]
  wire  _GEN_2 = array4kb_valid_0 & _T_8 == _T_9 & array4kb_0_flag_d; // @[TLB.scala 71:71 73:22 66:35]
  wire  _GEN_3 = array4kb_valid_0 & _T_8 == _T_9 & array4kb_0_flag_a; // @[TLB.scala 71:71 73:22 66:35]
  wire  _GEN_5 = array4kb_valid_0 & _T_8 == _T_9 & array4kb_0_flag_u; // @[TLB.scala 71:71 73:22 66:35]
  wire  _GEN_6 = array4kb_valid_0 & _T_8 == _T_9 & array4kb_0_flag_x; // @[TLB.scala 71:71 73:22 66:35]
  wire  _GEN_7 = array4kb_valid_0 & _T_8 == _T_9 & array4kb_0_flag_w; // @[TLB.scala 71:71 73:22 66:35]
  wire  _GEN_8 = array4kb_valid_0 & _T_8 == _T_9 & array4kb_0_flag_r; // @[TLB.scala 71:71 73:22 66:35]
  wire  _GEN_9 = array4kb_valid_0 & _T_8 == _T_9 & array4kb_0_flag_v; // @[TLB.scala 71:71 73:22 66:35]
  wire [1:0] _GEN_13 = array4kb_valid_0 & _T_8 == _T_9 ? array4kb_0_ppn2 : 2'h0; // @[TLB.scala 71:71 73:22 66:35]
  wire [8:0] _GEN_14 = array4kb_valid_0 & _T_8 == _T_9 ? array4kb_0_ppn1 : 9'h0; // @[TLB.scala 71:71 73:22 66:35]
  wire [8:0] _GEN_15 = array4kb_valid_0 & _T_8 == _T_9 ? array4kb_0_ppn0 : 9'h0; // @[TLB.scala 71:71 73:22 66:35]
  wire [26:0] _T_12 = {array4kb_1_vpn2,array4kb_1_vpn1,array4kb_1_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_17 = array4kb_valid_1 & _T_12 == _T_9 ? array4kb_1_asid == io_satp_asid | array4kb_1_flag_g : _GEN_0; // @[TLB.scala 71:71 72:22]
  wire  _GEN_19 = array4kb_valid_1 & _T_12 == _T_9 ? array4kb_1_flag_d : _GEN_2; // @[TLB.scala 71:71 73:22]
  wire  _GEN_20 = array4kb_valid_1 & _T_12 == _T_9 ? array4kb_1_flag_a : _GEN_3; // @[TLB.scala 71:71 73:22]
  wire  _GEN_22 = array4kb_valid_1 & _T_12 == _T_9 ? array4kb_1_flag_u : _GEN_5; // @[TLB.scala 71:71 73:22]
  wire  _GEN_23 = array4kb_valid_1 & _T_12 == _T_9 ? array4kb_1_flag_x : _GEN_6; // @[TLB.scala 71:71 73:22]
  wire  _GEN_24 = array4kb_valid_1 & _T_12 == _T_9 ? array4kb_1_flag_w : _GEN_7; // @[TLB.scala 71:71 73:22]
  wire  _GEN_25 = array4kb_valid_1 & _T_12 == _T_9 ? array4kb_1_flag_r : _GEN_8; // @[TLB.scala 71:71 73:22]
  wire  _GEN_26 = array4kb_valid_1 & _T_12 == _T_9 ? array4kb_1_flag_v : _GEN_9; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_30 = array4kb_valid_1 & _T_12 == _T_9 ? array4kb_1_ppn2 : _GEN_13; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_31 = array4kb_valid_1 & _T_12 == _T_9 ? array4kb_1_ppn1 : _GEN_14; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_32 = array4kb_valid_1 & _T_12 == _T_9 ? array4kb_1_ppn0 : _GEN_15; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_16 = {array4kb_2_vpn2,array4kb_2_vpn1,array4kb_2_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_34 = array4kb_valid_2 & _T_16 == _T_9 ? array4kb_2_asid == io_satp_asid | array4kb_2_flag_g : _GEN_17; // @[TLB.scala 71:71 72:22]
  wire  _GEN_36 = array4kb_valid_2 & _T_16 == _T_9 ? array4kb_2_flag_d : _GEN_19; // @[TLB.scala 71:71 73:22]
  wire  _GEN_37 = array4kb_valid_2 & _T_16 == _T_9 ? array4kb_2_flag_a : _GEN_20; // @[TLB.scala 71:71 73:22]
  wire  _GEN_39 = array4kb_valid_2 & _T_16 == _T_9 ? array4kb_2_flag_u : _GEN_22; // @[TLB.scala 71:71 73:22]
  wire  _GEN_40 = array4kb_valid_2 & _T_16 == _T_9 ? array4kb_2_flag_x : _GEN_23; // @[TLB.scala 71:71 73:22]
  wire  _GEN_41 = array4kb_valid_2 & _T_16 == _T_9 ? array4kb_2_flag_w : _GEN_24; // @[TLB.scala 71:71 73:22]
  wire  _GEN_42 = array4kb_valid_2 & _T_16 == _T_9 ? array4kb_2_flag_r : _GEN_25; // @[TLB.scala 71:71 73:22]
  wire  _GEN_43 = array4kb_valid_2 & _T_16 == _T_9 ? array4kb_2_flag_v : _GEN_26; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_47 = array4kb_valid_2 & _T_16 == _T_9 ? array4kb_2_ppn2 : _GEN_30; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_48 = array4kb_valid_2 & _T_16 == _T_9 ? array4kb_2_ppn1 : _GEN_31; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_49 = array4kb_valid_2 & _T_16 == _T_9 ? array4kb_2_ppn0 : _GEN_32; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_20 = {array4kb_3_vpn2,array4kb_3_vpn1,array4kb_3_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_51 = array4kb_valid_3 & _T_20 == _T_9 ? array4kb_3_asid == io_satp_asid | array4kb_3_flag_g : _GEN_34; // @[TLB.scala 71:71 72:22]
  wire  _GEN_53 = array4kb_valid_3 & _T_20 == _T_9 ? array4kb_3_flag_d : _GEN_36; // @[TLB.scala 71:71 73:22]
  wire  _GEN_54 = array4kb_valid_3 & _T_20 == _T_9 ? array4kb_3_flag_a : _GEN_37; // @[TLB.scala 71:71 73:22]
  wire  _GEN_56 = array4kb_valid_3 & _T_20 == _T_9 ? array4kb_3_flag_u : _GEN_39; // @[TLB.scala 71:71 73:22]
  wire  _GEN_57 = array4kb_valid_3 & _T_20 == _T_9 ? array4kb_3_flag_x : _GEN_40; // @[TLB.scala 71:71 73:22]
  wire  _GEN_58 = array4kb_valid_3 & _T_20 == _T_9 ? array4kb_3_flag_w : _GEN_41; // @[TLB.scala 71:71 73:22]
  wire  _GEN_59 = array4kb_valid_3 & _T_20 == _T_9 ? array4kb_3_flag_r : _GEN_42; // @[TLB.scala 71:71 73:22]
  wire  _GEN_60 = array4kb_valid_3 & _T_20 == _T_9 ? array4kb_3_flag_v : _GEN_43; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_64 = array4kb_valid_3 & _T_20 == _T_9 ? array4kb_3_ppn2 : _GEN_47; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_65 = array4kb_valid_3 & _T_20 == _T_9 ? array4kb_3_ppn1 : _GEN_48; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_66 = array4kb_valid_3 & _T_20 == _T_9 ? array4kb_3_ppn0 : _GEN_49; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_24 = {array4kb_4_vpn2,array4kb_4_vpn1,array4kb_4_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_68 = array4kb_valid_4 & _T_24 == _T_9 ? array4kb_4_asid == io_satp_asid | array4kb_4_flag_g : _GEN_51; // @[TLB.scala 71:71 72:22]
  wire  _GEN_70 = array4kb_valid_4 & _T_24 == _T_9 ? array4kb_4_flag_d : _GEN_53; // @[TLB.scala 71:71 73:22]
  wire  _GEN_71 = array4kb_valid_4 & _T_24 == _T_9 ? array4kb_4_flag_a : _GEN_54; // @[TLB.scala 71:71 73:22]
  wire  _GEN_73 = array4kb_valid_4 & _T_24 == _T_9 ? array4kb_4_flag_u : _GEN_56; // @[TLB.scala 71:71 73:22]
  wire  _GEN_74 = array4kb_valid_4 & _T_24 == _T_9 ? array4kb_4_flag_x : _GEN_57; // @[TLB.scala 71:71 73:22]
  wire  _GEN_75 = array4kb_valid_4 & _T_24 == _T_9 ? array4kb_4_flag_w : _GEN_58; // @[TLB.scala 71:71 73:22]
  wire  _GEN_76 = array4kb_valid_4 & _T_24 == _T_9 ? array4kb_4_flag_r : _GEN_59; // @[TLB.scala 71:71 73:22]
  wire  _GEN_77 = array4kb_valid_4 & _T_24 == _T_9 ? array4kb_4_flag_v : _GEN_60; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_81 = array4kb_valid_4 & _T_24 == _T_9 ? array4kb_4_ppn2 : _GEN_64; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_82 = array4kb_valid_4 & _T_24 == _T_9 ? array4kb_4_ppn1 : _GEN_65; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_83 = array4kb_valid_4 & _T_24 == _T_9 ? array4kb_4_ppn0 : _GEN_66; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_28 = {array4kb_5_vpn2,array4kb_5_vpn1,array4kb_5_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_85 = array4kb_valid_5 & _T_28 == _T_9 ? array4kb_5_asid == io_satp_asid | array4kb_5_flag_g : _GEN_68; // @[TLB.scala 71:71 72:22]
  wire  _GEN_87 = array4kb_valid_5 & _T_28 == _T_9 ? array4kb_5_flag_d : _GEN_70; // @[TLB.scala 71:71 73:22]
  wire  _GEN_88 = array4kb_valid_5 & _T_28 == _T_9 ? array4kb_5_flag_a : _GEN_71; // @[TLB.scala 71:71 73:22]
  wire  _GEN_90 = array4kb_valid_5 & _T_28 == _T_9 ? array4kb_5_flag_u : _GEN_73; // @[TLB.scala 71:71 73:22]
  wire  _GEN_91 = array4kb_valid_5 & _T_28 == _T_9 ? array4kb_5_flag_x : _GEN_74; // @[TLB.scala 71:71 73:22]
  wire  _GEN_92 = array4kb_valid_5 & _T_28 == _T_9 ? array4kb_5_flag_w : _GEN_75; // @[TLB.scala 71:71 73:22]
  wire  _GEN_93 = array4kb_valid_5 & _T_28 == _T_9 ? array4kb_5_flag_r : _GEN_76; // @[TLB.scala 71:71 73:22]
  wire  _GEN_94 = array4kb_valid_5 & _T_28 == _T_9 ? array4kb_5_flag_v : _GEN_77; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_98 = array4kb_valid_5 & _T_28 == _T_9 ? array4kb_5_ppn2 : _GEN_81; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_99 = array4kb_valid_5 & _T_28 == _T_9 ? array4kb_5_ppn1 : _GEN_82; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_100 = array4kb_valid_5 & _T_28 == _T_9 ? array4kb_5_ppn0 : _GEN_83; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_32 = {array4kb_6_vpn2,array4kb_6_vpn1,array4kb_6_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_102 = array4kb_valid_6 & _T_32 == _T_9 ? array4kb_6_asid == io_satp_asid | array4kb_6_flag_g : _GEN_85; // @[TLB.scala 71:71 72:22]
  wire  _GEN_104 = array4kb_valid_6 & _T_32 == _T_9 ? array4kb_6_flag_d : _GEN_87; // @[TLB.scala 71:71 73:22]
  wire  _GEN_105 = array4kb_valid_6 & _T_32 == _T_9 ? array4kb_6_flag_a : _GEN_88; // @[TLB.scala 71:71 73:22]
  wire  _GEN_107 = array4kb_valid_6 & _T_32 == _T_9 ? array4kb_6_flag_u : _GEN_90; // @[TLB.scala 71:71 73:22]
  wire  _GEN_108 = array4kb_valid_6 & _T_32 == _T_9 ? array4kb_6_flag_x : _GEN_91; // @[TLB.scala 71:71 73:22]
  wire  _GEN_109 = array4kb_valid_6 & _T_32 == _T_9 ? array4kb_6_flag_w : _GEN_92; // @[TLB.scala 71:71 73:22]
  wire  _GEN_110 = array4kb_valid_6 & _T_32 == _T_9 ? array4kb_6_flag_r : _GEN_93; // @[TLB.scala 71:71 73:22]
  wire  _GEN_111 = array4kb_valid_6 & _T_32 == _T_9 ? array4kb_6_flag_v : _GEN_94; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_115 = array4kb_valid_6 & _T_32 == _T_9 ? array4kb_6_ppn2 : _GEN_98; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_116 = array4kb_valid_6 & _T_32 == _T_9 ? array4kb_6_ppn1 : _GEN_99; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_117 = array4kb_valid_6 & _T_32 == _T_9 ? array4kb_6_ppn0 : _GEN_100; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_36 = {array4kb_7_vpn2,array4kb_7_vpn1,array4kb_7_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_119 = array4kb_valid_7 & _T_36 == _T_9 ? array4kb_7_asid == io_satp_asid | array4kb_7_flag_g : _GEN_102; // @[TLB.scala 71:71 72:22]
  wire  _GEN_121 = array4kb_valid_7 & _T_36 == _T_9 ? array4kb_7_flag_d : _GEN_104; // @[TLB.scala 71:71 73:22]
  wire  _GEN_122 = array4kb_valid_7 & _T_36 == _T_9 ? array4kb_7_flag_a : _GEN_105; // @[TLB.scala 71:71 73:22]
  wire  _GEN_124 = array4kb_valid_7 & _T_36 == _T_9 ? array4kb_7_flag_u : _GEN_107; // @[TLB.scala 71:71 73:22]
  wire  _GEN_125 = array4kb_valid_7 & _T_36 == _T_9 ? array4kb_7_flag_x : _GEN_108; // @[TLB.scala 71:71 73:22]
  wire  _GEN_126 = array4kb_valid_7 & _T_36 == _T_9 ? array4kb_7_flag_w : _GEN_109; // @[TLB.scala 71:71 73:22]
  wire  _GEN_127 = array4kb_valid_7 & _T_36 == _T_9 ? array4kb_7_flag_r : _GEN_110; // @[TLB.scala 71:71 73:22]
  wire  _GEN_128 = array4kb_valid_7 & _T_36 == _T_9 ? array4kb_7_flag_v : _GEN_111; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_132 = array4kb_valid_7 & _T_36 == _T_9 ? array4kb_7_ppn2 : _GEN_115; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_133 = array4kb_valid_7 & _T_36 == _T_9 ? array4kb_7_ppn1 : _GEN_116; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_134 = array4kb_valid_7 & _T_36 == _T_9 ? array4kb_7_ppn0 : _GEN_117; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_40 = {array4kb_8_vpn2,array4kb_8_vpn1,array4kb_8_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_136 = array4kb_valid_8 & _T_40 == _T_9 ? array4kb_8_asid == io_satp_asid | array4kb_8_flag_g : _GEN_119; // @[TLB.scala 71:71 72:22]
  wire  _GEN_138 = array4kb_valid_8 & _T_40 == _T_9 ? array4kb_8_flag_d : _GEN_121; // @[TLB.scala 71:71 73:22]
  wire  _GEN_139 = array4kb_valid_8 & _T_40 == _T_9 ? array4kb_8_flag_a : _GEN_122; // @[TLB.scala 71:71 73:22]
  wire  _GEN_141 = array4kb_valid_8 & _T_40 == _T_9 ? array4kb_8_flag_u : _GEN_124; // @[TLB.scala 71:71 73:22]
  wire  _GEN_142 = array4kb_valid_8 & _T_40 == _T_9 ? array4kb_8_flag_x : _GEN_125; // @[TLB.scala 71:71 73:22]
  wire  _GEN_143 = array4kb_valid_8 & _T_40 == _T_9 ? array4kb_8_flag_w : _GEN_126; // @[TLB.scala 71:71 73:22]
  wire  _GEN_144 = array4kb_valid_8 & _T_40 == _T_9 ? array4kb_8_flag_r : _GEN_127; // @[TLB.scala 71:71 73:22]
  wire  _GEN_145 = array4kb_valid_8 & _T_40 == _T_9 ? array4kb_8_flag_v : _GEN_128; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_149 = array4kb_valid_8 & _T_40 == _T_9 ? array4kb_8_ppn2 : _GEN_132; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_150 = array4kb_valid_8 & _T_40 == _T_9 ? array4kb_8_ppn1 : _GEN_133; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_151 = array4kb_valid_8 & _T_40 == _T_9 ? array4kb_8_ppn0 : _GEN_134; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_44 = {array4kb_9_vpn2,array4kb_9_vpn1,array4kb_9_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_153 = array4kb_valid_9 & _T_44 == _T_9 ? array4kb_9_asid == io_satp_asid | array4kb_9_flag_g : _GEN_136; // @[TLB.scala 71:71 72:22]
  wire  _GEN_155 = array4kb_valid_9 & _T_44 == _T_9 ? array4kb_9_flag_d : _GEN_138; // @[TLB.scala 71:71 73:22]
  wire  _GEN_156 = array4kb_valid_9 & _T_44 == _T_9 ? array4kb_9_flag_a : _GEN_139; // @[TLB.scala 71:71 73:22]
  wire  _GEN_158 = array4kb_valid_9 & _T_44 == _T_9 ? array4kb_9_flag_u : _GEN_141; // @[TLB.scala 71:71 73:22]
  wire  _GEN_159 = array4kb_valid_9 & _T_44 == _T_9 ? array4kb_9_flag_x : _GEN_142; // @[TLB.scala 71:71 73:22]
  wire  _GEN_160 = array4kb_valid_9 & _T_44 == _T_9 ? array4kb_9_flag_w : _GEN_143; // @[TLB.scala 71:71 73:22]
  wire  _GEN_161 = array4kb_valid_9 & _T_44 == _T_9 ? array4kb_9_flag_r : _GEN_144; // @[TLB.scala 71:71 73:22]
  wire  _GEN_162 = array4kb_valid_9 & _T_44 == _T_9 ? array4kb_9_flag_v : _GEN_145; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_166 = array4kb_valid_9 & _T_44 == _T_9 ? array4kb_9_ppn2 : _GEN_149; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_167 = array4kb_valid_9 & _T_44 == _T_9 ? array4kb_9_ppn1 : _GEN_150; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_168 = array4kb_valid_9 & _T_44 == _T_9 ? array4kb_9_ppn0 : _GEN_151; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_48 = {array4kb_10_vpn2,array4kb_10_vpn1,array4kb_10_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_170 = array4kb_valid_10 & _T_48 == _T_9 ? array4kb_10_asid == io_satp_asid | array4kb_10_flag_g : _GEN_153; // @[TLB.scala 71:71 72:22]
  wire  _GEN_172 = array4kb_valid_10 & _T_48 == _T_9 ? array4kb_10_flag_d : _GEN_155; // @[TLB.scala 71:71 73:22]
  wire  _GEN_173 = array4kb_valid_10 & _T_48 == _T_9 ? array4kb_10_flag_a : _GEN_156; // @[TLB.scala 71:71 73:22]
  wire  _GEN_175 = array4kb_valid_10 & _T_48 == _T_9 ? array4kb_10_flag_u : _GEN_158; // @[TLB.scala 71:71 73:22]
  wire  _GEN_176 = array4kb_valid_10 & _T_48 == _T_9 ? array4kb_10_flag_x : _GEN_159; // @[TLB.scala 71:71 73:22]
  wire  _GEN_177 = array4kb_valid_10 & _T_48 == _T_9 ? array4kb_10_flag_w : _GEN_160; // @[TLB.scala 71:71 73:22]
  wire  _GEN_178 = array4kb_valid_10 & _T_48 == _T_9 ? array4kb_10_flag_r : _GEN_161; // @[TLB.scala 71:71 73:22]
  wire  _GEN_179 = array4kb_valid_10 & _T_48 == _T_9 ? array4kb_10_flag_v : _GEN_162; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_183 = array4kb_valid_10 & _T_48 == _T_9 ? array4kb_10_ppn2 : _GEN_166; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_184 = array4kb_valid_10 & _T_48 == _T_9 ? array4kb_10_ppn1 : _GEN_167; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_185 = array4kb_valid_10 & _T_48 == _T_9 ? array4kb_10_ppn0 : _GEN_168; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_52 = {array4kb_11_vpn2,array4kb_11_vpn1,array4kb_11_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_187 = array4kb_valid_11 & _T_52 == _T_9 ? array4kb_11_asid == io_satp_asid | array4kb_11_flag_g : _GEN_170; // @[TLB.scala 71:71 72:22]
  wire  _GEN_189 = array4kb_valid_11 & _T_52 == _T_9 ? array4kb_11_flag_d : _GEN_172; // @[TLB.scala 71:71 73:22]
  wire  _GEN_190 = array4kb_valid_11 & _T_52 == _T_9 ? array4kb_11_flag_a : _GEN_173; // @[TLB.scala 71:71 73:22]
  wire  _GEN_192 = array4kb_valid_11 & _T_52 == _T_9 ? array4kb_11_flag_u : _GEN_175; // @[TLB.scala 71:71 73:22]
  wire  _GEN_193 = array4kb_valid_11 & _T_52 == _T_9 ? array4kb_11_flag_x : _GEN_176; // @[TLB.scala 71:71 73:22]
  wire  _GEN_194 = array4kb_valid_11 & _T_52 == _T_9 ? array4kb_11_flag_w : _GEN_177; // @[TLB.scala 71:71 73:22]
  wire  _GEN_195 = array4kb_valid_11 & _T_52 == _T_9 ? array4kb_11_flag_r : _GEN_178; // @[TLB.scala 71:71 73:22]
  wire  _GEN_196 = array4kb_valid_11 & _T_52 == _T_9 ? array4kb_11_flag_v : _GEN_179; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_200 = array4kb_valid_11 & _T_52 == _T_9 ? array4kb_11_ppn2 : _GEN_183; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_201 = array4kb_valid_11 & _T_52 == _T_9 ? array4kb_11_ppn1 : _GEN_184; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_202 = array4kb_valid_11 & _T_52 == _T_9 ? array4kb_11_ppn0 : _GEN_185; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_56 = {array4kb_12_vpn2,array4kb_12_vpn1,array4kb_12_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_204 = array4kb_valid_12 & _T_56 == _T_9 ? array4kb_12_asid == io_satp_asid | array4kb_12_flag_g : _GEN_187; // @[TLB.scala 71:71 72:22]
  wire  _GEN_206 = array4kb_valid_12 & _T_56 == _T_9 ? array4kb_12_flag_d : _GEN_189; // @[TLB.scala 71:71 73:22]
  wire  _GEN_207 = array4kb_valid_12 & _T_56 == _T_9 ? array4kb_12_flag_a : _GEN_190; // @[TLB.scala 71:71 73:22]
  wire  _GEN_209 = array4kb_valid_12 & _T_56 == _T_9 ? array4kb_12_flag_u : _GEN_192; // @[TLB.scala 71:71 73:22]
  wire  _GEN_210 = array4kb_valid_12 & _T_56 == _T_9 ? array4kb_12_flag_x : _GEN_193; // @[TLB.scala 71:71 73:22]
  wire  _GEN_211 = array4kb_valid_12 & _T_56 == _T_9 ? array4kb_12_flag_w : _GEN_194; // @[TLB.scala 71:71 73:22]
  wire  _GEN_212 = array4kb_valid_12 & _T_56 == _T_9 ? array4kb_12_flag_r : _GEN_195; // @[TLB.scala 71:71 73:22]
  wire  _GEN_213 = array4kb_valid_12 & _T_56 == _T_9 ? array4kb_12_flag_v : _GEN_196; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_217 = array4kb_valid_12 & _T_56 == _T_9 ? array4kb_12_ppn2 : _GEN_200; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_218 = array4kb_valid_12 & _T_56 == _T_9 ? array4kb_12_ppn1 : _GEN_201; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_219 = array4kb_valid_12 & _T_56 == _T_9 ? array4kb_12_ppn0 : _GEN_202; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_60 = {array4kb_13_vpn2,array4kb_13_vpn1,array4kb_13_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_221 = array4kb_valid_13 & _T_60 == _T_9 ? array4kb_13_asid == io_satp_asid | array4kb_13_flag_g : _GEN_204; // @[TLB.scala 71:71 72:22]
  wire  _GEN_223 = array4kb_valid_13 & _T_60 == _T_9 ? array4kb_13_flag_d : _GEN_206; // @[TLB.scala 71:71 73:22]
  wire  _GEN_224 = array4kb_valid_13 & _T_60 == _T_9 ? array4kb_13_flag_a : _GEN_207; // @[TLB.scala 71:71 73:22]
  wire  _GEN_226 = array4kb_valid_13 & _T_60 == _T_9 ? array4kb_13_flag_u : _GEN_209; // @[TLB.scala 71:71 73:22]
  wire  _GEN_227 = array4kb_valid_13 & _T_60 == _T_9 ? array4kb_13_flag_x : _GEN_210; // @[TLB.scala 71:71 73:22]
  wire  _GEN_228 = array4kb_valid_13 & _T_60 == _T_9 ? array4kb_13_flag_w : _GEN_211; // @[TLB.scala 71:71 73:22]
  wire  _GEN_229 = array4kb_valid_13 & _T_60 == _T_9 ? array4kb_13_flag_r : _GEN_212; // @[TLB.scala 71:71 73:22]
  wire  _GEN_230 = array4kb_valid_13 & _T_60 == _T_9 ? array4kb_13_flag_v : _GEN_213; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_234 = array4kb_valid_13 & _T_60 == _T_9 ? array4kb_13_ppn2 : _GEN_217; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_235 = array4kb_valid_13 & _T_60 == _T_9 ? array4kb_13_ppn1 : _GEN_218; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_236 = array4kb_valid_13 & _T_60 == _T_9 ? array4kb_13_ppn0 : _GEN_219; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_64 = {array4kb_14_vpn2,array4kb_14_vpn1,array4kb_14_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_238 = array4kb_valid_14 & _T_64 == _T_9 ? array4kb_14_asid == io_satp_asid | array4kb_14_flag_g : _GEN_221; // @[TLB.scala 71:71 72:22]
  wire  _GEN_240 = array4kb_valid_14 & _T_64 == _T_9 ? array4kb_14_flag_d : _GEN_223; // @[TLB.scala 71:71 73:22]
  wire  _GEN_241 = array4kb_valid_14 & _T_64 == _T_9 ? array4kb_14_flag_a : _GEN_224; // @[TLB.scala 71:71 73:22]
  wire  _GEN_243 = array4kb_valid_14 & _T_64 == _T_9 ? array4kb_14_flag_u : _GEN_226; // @[TLB.scala 71:71 73:22]
  wire  _GEN_244 = array4kb_valid_14 & _T_64 == _T_9 ? array4kb_14_flag_x : _GEN_227; // @[TLB.scala 71:71 73:22]
  wire  _GEN_245 = array4kb_valid_14 & _T_64 == _T_9 ? array4kb_14_flag_w : _GEN_228; // @[TLB.scala 71:71 73:22]
  wire  _GEN_246 = array4kb_valid_14 & _T_64 == _T_9 ? array4kb_14_flag_r : _GEN_229; // @[TLB.scala 71:71 73:22]
  wire  _GEN_247 = array4kb_valid_14 & _T_64 == _T_9 ? array4kb_14_flag_v : _GEN_230; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_251 = array4kb_valid_14 & _T_64 == _T_9 ? array4kb_14_ppn2 : _GEN_234; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_252 = array4kb_valid_14 & _T_64 == _T_9 ? array4kb_14_ppn1 : _GEN_235; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_253 = array4kb_valid_14 & _T_64 == _T_9 ? array4kb_14_ppn0 : _GEN_236; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_68 = {array4kb_15_vpn2,array4kb_15_vpn1,array4kb_15_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_255 = array4kb_valid_15 & _T_68 == _T_9 ? array4kb_15_asid == io_satp_asid | array4kb_15_flag_g : _GEN_238; // @[TLB.scala 71:71 72:22]
  wire  _GEN_257 = array4kb_valid_15 & _T_68 == _T_9 ? array4kb_15_flag_d : _GEN_240; // @[TLB.scala 71:71 73:22]
  wire  _GEN_258 = array4kb_valid_15 & _T_68 == _T_9 ? array4kb_15_flag_a : _GEN_241; // @[TLB.scala 71:71 73:22]
  wire  _GEN_260 = array4kb_valid_15 & _T_68 == _T_9 ? array4kb_15_flag_u : _GEN_243; // @[TLB.scala 71:71 73:22]
  wire  _GEN_261 = array4kb_valid_15 & _T_68 == _T_9 ? array4kb_15_flag_x : _GEN_244; // @[TLB.scala 71:71 73:22]
  wire  _GEN_262 = array4kb_valid_15 & _T_68 == _T_9 ? array4kb_15_flag_w : _GEN_245; // @[TLB.scala 71:71 73:22]
  wire  _GEN_263 = array4kb_valid_15 & _T_68 == _T_9 ? array4kb_15_flag_r : _GEN_246; // @[TLB.scala 71:71 73:22]
  wire  _GEN_264 = array4kb_valid_15 & _T_68 == _T_9 ? array4kb_15_flag_v : _GEN_247; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_268 = array4kb_valid_15 & _T_68 == _T_9 ? array4kb_15_ppn2 : _GEN_251; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_269 = array4kb_valid_15 & _T_68 == _T_9 ? array4kb_15_ppn1 : _GEN_252; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_270 = array4kb_valid_15 & _T_68 == _T_9 ? array4kb_15_ppn0 : _GEN_253; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_72 = {array4kb_16_vpn2,array4kb_16_vpn1,array4kb_16_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_272 = array4kb_valid_16 & _T_72 == _T_9 ? array4kb_16_asid == io_satp_asid | array4kb_16_flag_g : _GEN_255; // @[TLB.scala 71:71 72:22]
  wire  _GEN_274 = array4kb_valid_16 & _T_72 == _T_9 ? array4kb_16_flag_d : _GEN_257; // @[TLB.scala 71:71 73:22]
  wire  _GEN_275 = array4kb_valid_16 & _T_72 == _T_9 ? array4kb_16_flag_a : _GEN_258; // @[TLB.scala 71:71 73:22]
  wire  _GEN_277 = array4kb_valid_16 & _T_72 == _T_9 ? array4kb_16_flag_u : _GEN_260; // @[TLB.scala 71:71 73:22]
  wire  _GEN_278 = array4kb_valid_16 & _T_72 == _T_9 ? array4kb_16_flag_x : _GEN_261; // @[TLB.scala 71:71 73:22]
  wire  _GEN_279 = array4kb_valid_16 & _T_72 == _T_9 ? array4kb_16_flag_w : _GEN_262; // @[TLB.scala 71:71 73:22]
  wire  _GEN_280 = array4kb_valid_16 & _T_72 == _T_9 ? array4kb_16_flag_r : _GEN_263; // @[TLB.scala 71:71 73:22]
  wire  _GEN_281 = array4kb_valid_16 & _T_72 == _T_9 ? array4kb_16_flag_v : _GEN_264; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_285 = array4kb_valid_16 & _T_72 == _T_9 ? array4kb_16_ppn2 : _GEN_268; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_286 = array4kb_valid_16 & _T_72 == _T_9 ? array4kb_16_ppn1 : _GEN_269; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_287 = array4kb_valid_16 & _T_72 == _T_9 ? array4kb_16_ppn0 : _GEN_270; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_76 = {array4kb_17_vpn2,array4kb_17_vpn1,array4kb_17_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_289 = array4kb_valid_17 & _T_76 == _T_9 ? array4kb_17_asid == io_satp_asid | array4kb_17_flag_g : _GEN_272; // @[TLB.scala 71:71 72:22]
  wire  _GEN_291 = array4kb_valid_17 & _T_76 == _T_9 ? array4kb_17_flag_d : _GEN_274; // @[TLB.scala 71:71 73:22]
  wire  _GEN_292 = array4kb_valid_17 & _T_76 == _T_9 ? array4kb_17_flag_a : _GEN_275; // @[TLB.scala 71:71 73:22]
  wire  _GEN_294 = array4kb_valid_17 & _T_76 == _T_9 ? array4kb_17_flag_u : _GEN_277; // @[TLB.scala 71:71 73:22]
  wire  _GEN_295 = array4kb_valid_17 & _T_76 == _T_9 ? array4kb_17_flag_x : _GEN_278; // @[TLB.scala 71:71 73:22]
  wire  _GEN_296 = array4kb_valid_17 & _T_76 == _T_9 ? array4kb_17_flag_w : _GEN_279; // @[TLB.scala 71:71 73:22]
  wire  _GEN_297 = array4kb_valid_17 & _T_76 == _T_9 ? array4kb_17_flag_r : _GEN_280; // @[TLB.scala 71:71 73:22]
  wire  _GEN_298 = array4kb_valid_17 & _T_76 == _T_9 ? array4kb_17_flag_v : _GEN_281; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_302 = array4kb_valid_17 & _T_76 == _T_9 ? array4kb_17_ppn2 : _GEN_285; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_303 = array4kb_valid_17 & _T_76 == _T_9 ? array4kb_17_ppn1 : _GEN_286; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_304 = array4kb_valid_17 & _T_76 == _T_9 ? array4kb_17_ppn0 : _GEN_287; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_80 = {array4kb_18_vpn2,array4kb_18_vpn1,array4kb_18_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_306 = array4kb_valid_18 & _T_80 == _T_9 ? array4kb_18_asid == io_satp_asid | array4kb_18_flag_g : _GEN_289; // @[TLB.scala 71:71 72:22]
  wire  _GEN_308 = array4kb_valid_18 & _T_80 == _T_9 ? array4kb_18_flag_d : _GEN_291; // @[TLB.scala 71:71 73:22]
  wire  _GEN_309 = array4kb_valid_18 & _T_80 == _T_9 ? array4kb_18_flag_a : _GEN_292; // @[TLB.scala 71:71 73:22]
  wire  _GEN_311 = array4kb_valid_18 & _T_80 == _T_9 ? array4kb_18_flag_u : _GEN_294; // @[TLB.scala 71:71 73:22]
  wire  _GEN_312 = array4kb_valid_18 & _T_80 == _T_9 ? array4kb_18_flag_x : _GEN_295; // @[TLB.scala 71:71 73:22]
  wire  _GEN_313 = array4kb_valid_18 & _T_80 == _T_9 ? array4kb_18_flag_w : _GEN_296; // @[TLB.scala 71:71 73:22]
  wire  _GEN_314 = array4kb_valid_18 & _T_80 == _T_9 ? array4kb_18_flag_r : _GEN_297; // @[TLB.scala 71:71 73:22]
  wire  _GEN_315 = array4kb_valid_18 & _T_80 == _T_9 ? array4kb_18_flag_v : _GEN_298; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_319 = array4kb_valid_18 & _T_80 == _T_9 ? array4kb_18_ppn2 : _GEN_302; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_320 = array4kb_valid_18 & _T_80 == _T_9 ? array4kb_18_ppn1 : _GEN_303; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_321 = array4kb_valid_18 & _T_80 == _T_9 ? array4kb_18_ppn0 : _GEN_304; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_84 = {array4kb_19_vpn2,array4kb_19_vpn1,array4kb_19_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_323 = array4kb_valid_19 & _T_84 == _T_9 ? array4kb_19_asid == io_satp_asid | array4kb_19_flag_g : _GEN_306; // @[TLB.scala 71:71 72:22]
  wire  _GEN_325 = array4kb_valid_19 & _T_84 == _T_9 ? array4kb_19_flag_d : _GEN_308; // @[TLB.scala 71:71 73:22]
  wire  _GEN_326 = array4kb_valid_19 & _T_84 == _T_9 ? array4kb_19_flag_a : _GEN_309; // @[TLB.scala 71:71 73:22]
  wire  _GEN_328 = array4kb_valid_19 & _T_84 == _T_9 ? array4kb_19_flag_u : _GEN_311; // @[TLB.scala 71:71 73:22]
  wire  _GEN_329 = array4kb_valid_19 & _T_84 == _T_9 ? array4kb_19_flag_x : _GEN_312; // @[TLB.scala 71:71 73:22]
  wire  _GEN_330 = array4kb_valid_19 & _T_84 == _T_9 ? array4kb_19_flag_w : _GEN_313; // @[TLB.scala 71:71 73:22]
  wire  _GEN_331 = array4kb_valid_19 & _T_84 == _T_9 ? array4kb_19_flag_r : _GEN_314; // @[TLB.scala 71:71 73:22]
  wire  _GEN_332 = array4kb_valid_19 & _T_84 == _T_9 ? array4kb_19_flag_v : _GEN_315; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_336 = array4kb_valid_19 & _T_84 == _T_9 ? array4kb_19_ppn2 : _GEN_319; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_337 = array4kb_valid_19 & _T_84 == _T_9 ? array4kb_19_ppn1 : _GEN_320; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_338 = array4kb_valid_19 & _T_84 == _T_9 ? array4kb_19_ppn0 : _GEN_321; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_88 = {array4kb_20_vpn2,array4kb_20_vpn1,array4kb_20_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_340 = array4kb_valid_20 & _T_88 == _T_9 ? array4kb_20_asid == io_satp_asid | array4kb_20_flag_g : _GEN_323; // @[TLB.scala 71:71 72:22]
  wire  _GEN_342 = array4kb_valid_20 & _T_88 == _T_9 ? array4kb_20_flag_d : _GEN_325; // @[TLB.scala 71:71 73:22]
  wire  _GEN_343 = array4kb_valid_20 & _T_88 == _T_9 ? array4kb_20_flag_a : _GEN_326; // @[TLB.scala 71:71 73:22]
  wire  _GEN_345 = array4kb_valid_20 & _T_88 == _T_9 ? array4kb_20_flag_u : _GEN_328; // @[TLB.scala 71:71 73:22]
  wire  _GEN_346 = array4kb_valid_20 & _T_88 == _T_9 ? array4kb_20_flag_x : _GEN_329; // @[TLB.scala 71:71 73:22]
  wire  _GEN_347 = array4kb_valid_20 & _T_88 == _T_9 ? array4kb_20_flag_w : _GEN_330; // @[TLB.scala 71:71 73:22]
  wire  _GEN_348 = array4kb_valid_20 & _T_88 == _T_9 ? array4kb_20_flag_r : _GEN_331; // @[TLB.scala 71:71 73:22]
  wire  _GEN_349 = array4kb_valid_20 & _T_88 == _T_9 ? array4kb_20_flag_v : _GEN_332; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_353 = array4kb_valid_20 & _T_88 == _T_9 ? array4kb_20_ppn2 : _GEN_336; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_354 = array4kb_valid_20 & _T_88 == _T_9 ? array4kb_20_ppn1 : _GEN_337; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_355 = array4kb_valid_20 & _T_88 == _T_9 ? array4kb_20_ppn0 : _GEN_338; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_92 = {array4kb_21_vpn2,array4kb_21_vpn1,array4kb_21_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_357 = array4kb_valid_21 & _T_92 == _T_9 ? array4kb_21_asid == io_satp_asid | array4kb_21_flag_g : _GEN_340; // @[TLB.scala 71:71 72:22]
  wire  _GEN_359 = array4kb_valid_21 & _T_92 == _T_9 ? array4kb_21_flag_d : _GEN_342; // @[TLB.scala 71:71 73:22]
  wire  _GEN_360 = array4kb_valid_21 & _T_92 == _T_9 ? array4kb_21_flag_a : _GEN_343; // @[TLB.scala 71:71 73:22]
  wire  _GEN_362 = array4kb_valid_21 & _T_92 == _T_9 ? array4kb_21_flag_u : _GEN_345; // @[TLB.scala 71:71 73:22]
  wire  _GEN_363 = array4kb_valid_21 & _T_92 == _T_9 ? array4kb_21_flag_x : _GEN_346; // @[TLB.scala 71:71 73:22]
  wire  _GEN_364 = array4kb_valid_21 & _T_92 == _T_9 ? array4kb_21_flag_w : _GEN_347; // @[TLB.scala 71:71 73:22]
  wire  _GEN_365 = array4kb_valid_21 & _T_92 == _T_9 ? array4kb_21_flag_r : _GEN_348; // @[TLB.scala 71:71 73:22]
  wire  _GEN_366 = array4kb_valid_21 & _T_92 == _T_9 ? array4kb_21_flag_v : _GEN_349; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_370 = array4kb_valid_21 & _T_92 == _T_9 ? array4kb_21_ppn2 : _GEN_353; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_371 = array4kb_valid_21 & _T_92 == _T_9 ? array4kb_21_ppn1 : _GEN_354; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_372 = array4kb_valid_21 & _T_92 == _T_9 ? array4kb_21_ppn0 : _GEN_355; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_96 = {array4kb_22_vpn2,array4kb_22_vpn1,array4kb_22_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_374 = array4kb_valid_22 & _T_96 == _T_9 ? array4kb_22_asid == io_satp_asid | array4kb_22_flag_g : _GEN_357; // @[TLB.scala 71:71 72:22]
  wire  _GEN_376 = array4kb_valid_22 & _T_96 == _T_9 ? array4kb_22_flag_d : _GEN_359; // @[TLB.scala 71:71 73:22]
  wire  _GEN_377 = array4kb_valid_22 & _T_96 == _T_9 ? array4kb_22_flag_a : _GEN_360; // @[TLB.scala 71:71 73:22]
  wire  _GEN_379 = array4kb_valid_22 & _T_96 == _T_9 ? array4kb_22_flag_u : _GEN_362; // @[TLB.scala 71:71 73:22]
  wire  _GEN_380 = array4kb_valid_22 & _T_96 == _T_9 ? array4kb_22_flag_x : _GEN_363; // @[TLB.scala 71:71 73:22]
  wire  _GEN_381 = array4kb_valid_22 & _T_96 == _T_9 ? array4kb_22_flag_w : _GEN_364; // @[TLB.scala 71:71 73:22]
  wire  _GEN_382 = array4kb_valid_22 & _T_96 == _T_9 ? array4kb_22_flag_r : _GEN_365; // @[TLB.scala 71:71 73:22]
  wire  _GEN_383 = array4kb_valid_22 & _T_96 == _T_9 ? array4kb_22_flag_v : _GEN_366; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_387 = array4kb_valid_22 & _T_96 == _T_9 ? array4kb_22_ppn2 : _GEN_370; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_388 = array4kb_valid_22 & _T_96 == _T_9 ? array4kb_22_ppn1 : _GEN_371; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_389 = array4kb_valid_22 & _T_96 == _T_9 ? array4kb_22_ppn0 : _GEN_372; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_100 = {array4kb_23_vpn2,array4kb_23_vpn1,array4kb_23_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_391 = array4kb_valid_23 & _T_100 == _T_9 ? array4kb_23_asid == io_satp_asid | array4kb_23_flag_g : _GEN_374
    ; // @[TLB.scala 71:71 72:22]
  wire  _GEN_393 = array4kb_valid_23 & _T_100 == _T_9 ? array4kb_23_flag_d : _GEN_376; // @[TLB.scala 71:71 73:22]
  wire  _GEN_394 = array4kb_valid_23 & _T_100 == _T_9 ? array4kb_23_flag_a : _GEN_377; // @[TLB.scala 71:71 73:22]
  wire  _GEN_396 = array4kb_valid_23 & _T_100 == _T_9 ? array4kb_23_flag_u : _GEN_379; // @[TLB.scala 71:71 73:22]
  wire  _GEN_397 = array4kb_valid_23 & _T_100 == _T_9 ? array4kb_23_flag_x : _GEN_380; // @[TLB.scala 71:71 73:22]
  wire  _GEN_398 = array4kb_valid_23 & _T_100 == _T_9 ? array4kb_23_flag_w : _GEN_381; // @[TLB.scala 71:71 73:22]
  wire  _GEN_399 = array4kb_valid_23 & _T_100 == _T_9 ? array4kb_23_flag_r : _GEN_382; // @[TLB.scala 71:71 73:22]
  wire  _GEN_400 = array4kb_valid_23 & _T_100 == _T_9 ? array4kb_23_flag_v : _GEN_383; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_404 = array4kb_valid_23 & _T_100 == _T_9 ? array4kb_23_ppn2 : _GEN_387; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_405 = array4kb_valid_23 & _T_100 == _T_9 ? array4kb_23_ppn1 : _GEN_388; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_406 = array4kb_valid_23 & _T_100 == _T_9 ? array4kb_23_ppn0 : _GEN_389; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_104 = {array4kb_24_vpn2,array4kb_24_vpn1,array4kb_24_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_408 = array4kb_valid_24 & _T_104 == _T_9 ? array4kb_24_asid == io_satp_asid | array4kb_24_flag_g : _GEN_391
    ; // @[TLB.scala 71:71 72:22]
  wire  _GEN_410 = array4kb_valid_24 & _T_104 == _T_9 ? array4kb_24_flag_d : _GEN_393; // @[TLB.scala 71:71 73:22]
  wire  _GEN_411 = array4kb_valid_24 & _T_104 == _T_9 ? array4kb_24_flag_a : _GEN_394; // @[TLB.scala 71:71 73:22]
  wire  _GEN_413 = array4kb_valid_24 & _T_104 == _T_9 ? array4kb_24_flag_u : _GEN_396; // @[TLB.scala 71:71 73:22]
  wire  _GEN_414 = array4kb_valid_24 & _T_104 == _T_9 ? array4kb_24_flag_x : _GEN_397; // @[TLB.scala 71:71 73:22]
  wire  _GEN_415 = array4kb_valid_24 & _T_104 == _T_9 ? array4kb_24_flag_w : _GEN_398; // @[TLB.scala 71:71 73:22]
  wire  _GEN_416 = array4kb_valid_24 & _T_104 == _T_9 ? array4kb_24_flag_r : _GEN_399; // @[TLB.scala 71:71 73:22]
  wire  _GEN_417 = array4kb_valid_24 & _T_104 == _T_9 ? array4kb_24_flag_v : _GEN_400; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_421 = array4kb_valid_24 & _T_104 == _T_9 ? array4kb_24_ppn2 : _GEN_404; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_422 = array4kb_valid_24 & _T_104 == _T_9 ? array4kb_24_ppn1 : _GEN_405; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_423 = array4kb_valid_24 & _T_104 == _T_9 ? array4kb_24_ppn0 : _GEN_406; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_108 = {array4kb_25_vpn2,array4kb_25_vpn1,array4kb_25_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_425 = array4kb_valid_25 & _T_108 == _T_9 ? array4kb_25_asid == io_satp_asid | array4kb_25_flag_g : _GEN_408
    ; // @[TLB.scala 71:71 72:22]
  wire  _GEN_427 = array4kb_valid_25 & _T_108 == _T_9 ? array4kb_25_flag_d : _GEN_410; // @[TLB.scala 71:71 73:22]
  wire  _GEN_428 = array4kb_valid_25 & _T_108 == _T_9 ? array4kb_25_flag_a : _GEN_411; // @[TLB.scala 71:71 73:22]
  wire  _GEN_430 = array4kb_valid_25 & _T_108 == _T_9 ? array4kb_25_flag_u : _GEN_413; // @[TLB.scala 71:71 73:22]
  wire  _GEN_431 = array4kb_valid_25 & _T_108 == _T_9 ? array4kb_25_flag_x : _GEN_414; // @[TLB.scala 71:71 73:22]
  wire  _GEN_432 = array4kb_valid_25 & _T_108 == _T_9 ? array4kb_25_flag_w : _GEN_415; // @[TLB.scala 71:71 73:22]
  wire  _GEN_433 = array4kb_valid_25 & _T_108 == _T_9 ? array4kb_25_flag_r : _GEN_416; // @[TLB.scala 71:71 73:22]
  wire  _GEN_434 = array4kb_valid_25 & _T_108 == _T_9 ? array4kb_25_flag_v : _GEN_417; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_438 = array4kb_valid_25 & _T_108 == _T_9 ? array4kb_25_ppn2 : _GEN_421; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_439 = array4kb_valid_25 & _T_108 == _T_9 ? array4kb_25_ppn1 : _GEN_422; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_440 = array4kb_valid_25 & _T_108 == _T_9 ? array4kb_25_ppn0 : _GEN_423; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_112 = {array4kb_26_vpn2,array4kb_26_vpn1,array4kb_26_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_442 = array4kb_valid_26 & _T_112 == _T_9 ? array4kb_26_asid == io_satp_asid | array4kb_26_flag_g : _GEN_425
    ; // @[TLB.scala 71:71 72:22]
  wire  _GEN_444 = array4kb_valid_26 & _T_112 == _T_9 ? array4kb_26_flag_d : _GEN_427; // @[TLB.scala 71:71 73:22]
  wire  _GEN_445 = array4kb_valid_26 & _T_112 == _T_9 ? array4kb_26_flag_a : _GEN_428; // @[TLB.scala 71:71 73:22]
  wire  _GEN_447 = array4kb_valid_26 & _T_112 == _T_9 ? array4kb_26_flag_u : _GEN_430; // @[TLB.scala 71:71 73:22]
  wire  _GEN_448 = array4kb_valid_26 & _T_112 == _T_9 ? array4kb_26_flag_x : _GEN_431; // @[TLB.scala 71:71 73:22]
  wire  _GEN_449 = array4kb_valid_26 & _T_112 == _T_9 ? array4kb_26_flag_w : _GEN_432; // @[TLB.scala 71:71 73:22]
  wire  _GEN_450 = array4kb_valid_26 & _T_112 == _T_9 ? array4kb_26_flag_r : _GEN_433; // @[TLB.scala 71:71 73:22]
  wire  _GEN_451 = array4kb_valid_26 & _T_112 == _T_9 ? array4kb_26_flag_v : _GEN_434; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_455 = array4kb_valid_26 & _T_112 == _T_9 ? array4kb_26_ppn2 : _GEN_438; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_456 = array4kb_valid_26 & _T_112 == _T_9 ? array4kb_26_ppn1 : _GEN_439; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_457 = array4kb_valid_26 & _T_112 == _T_9 ? array4kb_26_ppn0 : _GEN_440; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_116 = {array4kb_27_vpn2,array4kb_27_vpn1,array4kb_27_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_459 = array4kb_valid_27 & _T_116 == _T_9 ? array4kb_27_asid == io_satp_asid | array4kb_27_flag_g : _GEN_442
    ; // @[TLB.scala 71:71 72:22]
  wire  _GEN_461 = array4kb_valid_27 & _T_116 == _T_9 ? array4kb_27_flag_d : _GEN_444; // @[TLB.scala 71:71 73:22]
  wire  _GEN_462 = array4kb_valid_27 & _T_116 == _T_9 ? array4kb_27_flag_a : _GEN_445; // @[TLB.scala 71:71 73:22]
  wire  _GEN_464 = array4kb_valid_27 & _T_116 == _T_9 ? array4kb_27_flag_u : _GEN_447; // @[TLB.scala 71:71 73:22]
  wire  _GEN_465 = array4kb_valid_27 & _T_116 == _T_9 ? array4kb_27_flag_x : _GEN_448; // @[TLB.scala 71:71 73:22]
  wire  _GEN_466 = array4kb_valid_27 & _T_116 == _T_9 ? array4kb_27_flag_w : _GEN_449; // @[TLB.scala 71:71 73:22]
  wire  _GEN_467 = array4kb_valid_27 & _T_116 == _T_9 ? array4kb_27_flag_r : _GEN_450; // @[TLB.scala 71:71 73:22]
  wire  _GEN_468 = array4kb_valid_27 & _T_116 == _T_9 ? array4kb_27_flag_v : _GEN_451; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_472 = array4kb_valid_27 & _T_116 == _T_9 ? array4kb_27_ppn2 : _GEN_455; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_473 = array4kb_valid_27 & _T_116 == _T_9 ? array4kb_27_ppn1 : _GEN_456; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_474 = array4kb_valid_27 & _T_116 == _T_9 ? array4kb_27_ppn0 : _GEN_457; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_120 = {array4kb_28_vpn2,array4kb_28_vpn1,array4kb_28_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_476 = array4kb_valid_28 & _T_120 == _T_9 ? array4kb_28_asid == io_satp_asid | array4kb_28_flag_g : _GEN_459
    ; // @[TLB.scala 71:71 72:22]
  wire  _GEN_478 = array4kb_valid_28 & _T_120 == _T_9 ? array4kb_28_flag_d : _GEN_461; // @[TLB.scala 71:71 73:22]
  wire  _GEN_479 = array4kb_valid_28 & _T_120 == _T_9 ? array4kb_28_flag_a : _GEN_462; // @[TLB.scala 71:71 73:22]
  wire  _GEN_481 = array4kb_valid_28 & _T_120 == _T_9 ? array4kb_28_flag_u : _GEN_464; // @[TLB.scala 71:71 73:22]
  wire  _GEN_482 = array4kb_valid_28 & _T_120 == _T_9 ? array4kb_28_flag_x : _GEN_465; // @[TLB.scala 71:71 73:22]
  wire  _GEN_483 = array4kb_valid_28 & _T_120 == _T_9 ? array4kb_28_flag_w : _GEN_466; // @[TLB.scala 71:71 73:22]
  wire  _GEN_484 = array4kb_valid_28 & _T_120 == _T_9 ? array4kb_28_flag_r : _GEN_467; // @[TLB.scala 71:71 73:22]
  wire  _GEN_485 = array4kb_valid_28 & _T_120 == _T_9 ? array4kb_28_flag_v : _GEN_468; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_489 = array4kb_valid_28 & _T_120 == _T_9 ? array4kb_28_ppn2 : _GEN_472; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_490 = array4kb_valid_28 & _T_120 == _T_9 ? array4kb_28_ppn1 : _GEN_473; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_491 = array4kb_valid_28 & _T_120 == _T_9 ? array4kb_28_ppn0 : _GEN_474; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_124 = {array4kb_29_vpn2,array4kb_29_vpn1,array4kb_29_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_493 = array4kb_valid_29 & _T_124 == _T_9 ? array4kb_29_asid == io_satp_asid | array4kb_29_flag_g : _GEN_476
    ; // @[TLB.scala 71:71 72:22]
  wire  _GEN_495 = array4kb_valid_29 & _T_124 == _T_9 ? array4kb_29_flag_d : _GEN_478; // @[TLB.scala 71:71 73:22]
  wire  _GEN_496 = array4kb_valid_29 & _T_124 == _T_9 ? array4kb_29_flag_a : _GEN_479; // @[TLB.scala 71:71 73:22]
  wire  _GEN_498 = array4kb_valid_29 & _T_124 == _T_9 ? array4kb_29_flag_u : _GEN_481; // @[TLB.scala 71:71 73:22]
  wire  _GEN_499 = array4kb_valid_29 & _T_124 == _T_9 ? array4kb_29_flag_x : _GEN_482; // @[TLB.scala 71:71 73:22]
  wire  _GEN_500 = array4kb_valid_29 & _T_124 == _T_9 ? array4kb_29_flag_w : _GEN_483; // @[TLB.scala 71:71 73:22]
  wire  _GEN_501 = array4kb_valid_29 & _T_124 == _T_9 ? array4kb_29_flag_r : _GEN_484; // @[TLB.scala 71:71 73:22]
  wire  _GEN_502 = array4kb_valid_29 & _T_124 == _T_9 ? array4kb_29_flag_v : _GEN_485; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_506 = array4kb_valid_29 & _T_124 == _T_9 ? array4kb_29_ppn2 : _GEN_489; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_507 = array4kb_valid_29 & _T_124 == _T_9 ? array4kb_29_ppn1 : _GEN_490; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_508 = array4kb_valid_29 & _T_124 == _T_9 ? array4kb_29_ppn0 : _GEN_491; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_128 = {array4kb_30_vpn2,array4kb_30_vpn1,array4kb_30_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_510 = array4kb_valid_30 & _T_128 == _T_9 ? array4kb_30_asid == io_satp_asid | array4kb_30_flag_g : _GEN_493
    ; // @[TLB.scala 71:71 72:22]
  wire  _GEN_512 = array4kb_valid_30 & _T_128 == _T_9 ? array4kb_30_flag_d : _GEN_495; // @[TLB.scala 71:71 73:22]
  wire  _GEN_513 = array4kb_valid_30 & _T_128 == _T_9 ? array4kb_30_flag_a : _GEN_496; // @[TLB.scala 71:71 73:22]
  wire  _GEN_515 = array4kb_valid_30 & _T_128 == _T_9 ? array4kb_30_flag_u : _GEN_498; // @[TLB.scala 71:71 73:22]
  wire  _GEN_516 = array4kb_valid_30 & _T_128 == _T_9 ? array4kb_30_flag_x : _GEN_499; // @[TLB.scala 71:71 73:22]
  wire  _GEN_517 = array4kb_valid_30 & _T_128 == _T_9 ? array4kb_30_flag_w : _GEN_500; // @[TLB.scala 71:71 73:22]
  wire  _GEN_518 = array4kb_valid_30 & _T_128 == _T_9 ? array4kb_30_flag_r : _GEN_501; // @[TLB.scala 71:71 73:22]
  wire  _GEN_519 = array4kb_valid_30 & _T_128 == _T_9 ? array4kb_30_flag_v : _GEN_502; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_523 = array4kb_valid_30 & _T_128 == _T_9 ? array4kb_30_ppn2 : _GEN_506; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_524 = array4kb_valid_30 & _T_128 == _T_9 ? array4kb_30_ppn1 : _GEN_507; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_525 = array4kb_valid_30 & _T_128 == _T_9 ? array4kb_30_ppn0 : _GEN_508; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_132 = {array4kb_31_vpn2,array4kb_31_vpn1,array4kb_31_vpn0}; // @[Cat.scala 33:92]
  wire  hit4kb = array4kb_valid_31 & _T_132 == _T_9 ? array4kb_31_asid == io_satp_asid | array4kb_31_flag_g : _GEN_510; // @[TLB.scala 71:71 72:22]
  wire  array4kb_rdata_flag_d = array4kb_valid_31 & _T_132 == _T_9 ? array4kb_31_flag_d : _GEN_512; // @[TLB.scala 71:71 73:22]
  wire  array4kb_rdata_flag_a = array4kb_valid_31 & _T_132 == _T_9 ? array4kb_31_flag_a : _GEN_513; // @[TLB.scala 71:71 73:22]
  wire  array4kb_rdata_flag_u = array4kb_valid_31 & _T_132 == _T_9 ? array4kb_31_flag_u : _GEN_515; // @[TLB.scala 71:71 73:22]
  wire  array4kb_rdata_flag_x = array4kb_valid_31 & _T_132 == _T_9 ? array4kb_31_flag_x : _GEN_516; // @[TLB.scala 71:71 73:22]
  wire  array4kb_rdata_flag_w = array4kb_valid_31 & _T_132 == _T_9 ? array4kb_31_flag_w : _GEN_517; // @[TLB.scala 71:71 73:22]
  wire  array4kb_rdata_flag_r = array4kb_valid_31 & _T_132 == _T_9 ? array4kb_31_flag_r : _GEN_518; // @[TLB.scala 71:71 73:22]
  wire  array4kb_rdata_flag_v = array4kb_valid_31 & _T_132 == _T_9 ? array4kb_31_flag_v : _GEN_519; // @[TLB.scala 71:71 73:22]
  wire [1:0] array4kb_rdata_ppn2 = array4kb_valid_31 & _T_132 == _T_9 ? array4kb_31_ppn2 : _GEN_523; // @[TLB.scala 71:71 73:22]
  wire [8:0] array4kb_rdata_ppn1 = array4kb_valid_31 & _T_132 == _T_9 ? array4kb_31_ppn1 : _GEN_524; // @[TLB.scala 71:71 73:22]
  wire [8:0] array4kb_rdata_ppn0 = array4kb_valid_31 & _T_132 == _T_9 ? array4kb_31_ppn0 : _GEN_525; // @[TLB.scala 71:71 73:22]
  wire  _GEN_1056 = 5'h0 == replace_idx | array4kb_valid_0; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1057 = 5'h1 == replace_idx | array4kb_valid_1; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1058 = 5'h2 == replace_idx | array4kb_valid_2; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1059 = 5'h3 == replace_idx | array4kb_valid_3; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1060 = 5'h4 == replace_idx | array4kb_valid_4; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1061 = 5'h5 == replace_idx | array4kb_valid_5; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1062 = 5'h6 == replace_idx | array4kb_valid_6; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1063 = 5'h7 == replace_idx | array4kb_valid_7; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1064 = 5'h8 == replace_idx | array4kb_valid_8; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1065 = 5'h9 == replace_idx | array4kb_valid_9; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1066 = 5'ha == replace_idx | array4kb_valid_10; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1067 = 5'hb == replace_idx | array4kb_valid_11; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1068 = 5'hc == replace_idx | array4kb_valid_12; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1069 = 5'hd == replace_idx | array4kb_valid_13; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1070 = 5'he == replace_idx | array4kb_valid_14; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1071 = 5'hf == replace_idx | array4kb_valid_15; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1072 = 5'h10 == replace_idx | array4kb_valid_16; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1073 = 5'h11 == replace_idx | array4kb_valid_17; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1074 = 5'h12 == replace_idx | array4kb_valid_18; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1075 = 5'h13 == replace_idx | array4kb_valid_19; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1076 = 5'h14 == replace_idx | array4kb_valid_20; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1077 = 5'h15 == replace_idx | array4kb_valid_21; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1078 = 5'h16 == replace_idx | array4kb_valid_22; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1079 = 5'h17 == replace_idx | array4kb_valid_23; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1080 = 5'h18 == replace_idx | array4kb_valid_24; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1081 = 5'h19 == replace_idx | array4kb_valid_25; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1082 = 5'h1a == replace_idx | array4kb_valid_26; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1083 = 5'h1b == replace_idx | array4kb_valid_27; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1084 = 5'h1c == replace_idx | array4kb_valid_28; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1085 = 5'h1d == replace_idx | array4kb_valid_29; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1086 = 5'h1e == replace_idx | array4kb_valid_30; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1087 = 5'h1f == replace_idx | array4kb_valid_31; // @[TLB.scala 65:31 87:{33,33}]
  reg  array2mb_0_flag_d; // @[TLB.scala 98:31]
  reg  array2mb_0_flag_a; // @[TLB.scala 98:31]
  reg  array2mb_0_flag_g; // @[TLB.scala 98:31]
  reg  array2mb_0_flag_u; // @[TLB.scala 98:31]
  reg  array2mb_0_flag_x; // @[TLB.scala 98:31]
  reg  array2mb_0_flag_w; // @[TLB.scala 98:31]
  reg  array2mb_0_flag_r; // @[TLB.scala 98:31]
  reg  array2mb_0_flag_v; // @[TLB.scala 98:31]
  reg [8:0] array2mb_0_vpn2; // @[TLB.scala 98:31]
  reg [8:0] array2mb_0_vpn1; // @[TLB.scala 98:31]
  reg [1:0] array2mb_0_ppn2; // @[TLB.scala 98:31]
  reg [8:0] array2mb_0_ppn1; // @[TLB.scala 98:31]
  reg [15:0] array2mb_0_asid; // @[TLB.scala 98:31]
  reg  array2mb_1_flag_d; // @[TLB.scala 98:31]
  reg  array2mb_1_flag_a; // @[TLB.scala 98:31]
  reg  array2mb_1_flag_g; // @[TLB.scala 98:31]
  reg  array2mb_1_flag_u; // @[TLB.scala 98:31]
  reg  array2mb_1_flag_x; // @[TLB.scala 98:31]
  reg  array2mb_1_flag_w; // @[TLB.scala 98:31]
  reg  array2mb_1_flag_r; // @[TLB.scala 98:31]
  reg  array2mb_1_flag_v; // @[TLB.scala 98:31]
  reg [8:0] array2mb_1_vpn2; // @[TLB.scala 98:31]
  reg [8:0] array2mb_1_vpn1; // @[TLB.scala 98:31]
  reg [1:0] array2mb_1_ppn2; // @[TLB.scala 98:31]
  reg [8:0] array2mb_1_ppn1; // @[TLB.scala 98:31]
  reg [15:0] array2mb_1_asid; // @[TLB.scala 98:31]
  reg  array2mb_2_flag_d; // @[TLB.scala 98:31]
  reg  array2mb_2_flag_a; // @[TLB.scala 98:31]
  reg  array2mb_2_flag_g; // @[TLB.scala 98:31]
  reg  array2mb_2_flag_u; // @[TLB.scala 98:31]
  reg  array2mb_2_flag_x; // @[TLB.scala 98:31]
  reg  array2mb_2_flag_w; // @[TLB.scala 98:31]
  reg  array2mb_2_flag_r; // @[TLB.scala 98:31]
  reg  array2mb_2_flag_v; // @[TLB.scala 98:31]
  reg [8:0] array2mb_2_vpn2; // @[TLB.scala 98:31]
  reg [8:0] array2mb_2_vpn1; // @[TLB.scala 98:31]
  reg [1:0] array2mb_2_ppn2; // @[TLB.scala 98:31]
  reg [8:0] array2mb_2_ppn1; // @[TLB.scala 98:31]
  reg [15:0] array2mb_2_asid; // @[TLB.scala 98:31]
  reg  array2mb_3_flag_d; // @[TLB.scala 98:31]
  reg  array2mb_3_flag_a; // @[TLB.scala 98:31]
  reg  array2mb_3_flag_g; // @[TLB.scala 98:31]
  reg  array2mb_3_flag_u; // @[TLB.scala 98:31]
  reg  array2mb_3_flag_x; // @[TLB.scala 98:31]
  reg  array2mb_3_flag_w; // @[TLB.scala 98:31]
  reg  array2mb_3_flag_r; // @[TLB.scala 98:31]
  reg  array2mb_3_flag_v; // @[TLB.scala 98:31]
  reg [8:0] array2mb_3_vpn2; // @[TLB.scala 98:31]
  reg [8:0] array2mb_3_vpn1; // @[TLB.scala 98:31]
  reg [1:0] array2mb_3_ppn2; // @[TLB.scala 98:31]
  reg [8:0] array2mb_3_ppn1; // @[TLB.scala 98:31]
  reg [15:0] array2mb_3_asid; // @[TLB.scala 98:31]
  reg  array2mb_4_flag_d; // @[TLB.scala 98:31]
  reg  array2mb_4_flag_a; // @[TLB.scala 98:31]
  reg  array2mb_4_flag_g; // @[TLB.scala 98:31]
  reg  array2mb_4_flag_u; // @[TLB.scala 98:31]
  reg  array2mb_4_flag_x; // @[TLB.scala 98:31]
  reg  array2mb_4_flag_w; // @[TLB.scala 98:31]
  reg  array2mb_4_flag_r; // @[TLB.scala 98:31]
  reg  array2mb_4_flag_v; // @[TLB.scala 98:31]
  reg [8:0] array2mb_4_vpn2; // @[TLB.scala 98:31]
  reg [8:0] array2mb_4_vpn1; // @[TLB.scala 98:31]
  reg [1:0] array2mb_4_ppn2; // @[TLB.scala 98:31]
  reg [8:0] array2mb_4_ppn1; // @[TLB.scala 98:31]
  reg [15:0] array2mb_4_asid; // @[TLB.scala 98:31]
  reg  array2mb_5_flag_d; // @[TLB.scala 98:31]
  reg  array2mb_5_flag_a; // @[TLB.scala 98:31]
  reg  array2mb_5_flag_g; // @[TLB.scala 98:31]
  reg  array2mb_5_flag_u; // @[TLB.scala 98:31]
  reg  array2mb_5_flag_x; // @[TLB.scala 98:31]
  reg  array2mb_5_flag_w; // @[TLB.scala 98:31]
  reg  array2mb_5_flag_r; // @[TLB.scala 98:31]
  reg  array2mb_5_flag_v; // @[TLB.scala 98:31]
  reg [8:0] array2mb_5_vpn2; // @[TLB.scala 98:31]
  reg [8:0] array2mb_5_vpn1; // @[TLB.scala 98:31]
  reg [1:0] array2mb_5_ppn2; // @[TLB.scala 98:31]
  reg [8:0] array2mb_5_ppn1; // @[TLB.scala 98:31]
  reg [15:0] array2mb_5_asid; // @[TLB.scala 98:31]
  reg  array2mb_6_flag_d; // @[TLB.scala 98:31]
  reg  array2mb_6_flag_a; // @[TLB.scala 98:31]
  reg  array2mb_6_flag_g; // @[TLB.scala 98:31]
  reg  array2mb_6_flag_u; // @[TLB.scala 98:31]
  reg  array2mb_6_flag_x; // @[TLB.scala 98:31]
  reg  array2mb_6_flag_w; // @[TLB.scala 98:31]
  reg  array2mb_6_flag_r; // @[TLB.scala 98:31]
  reg  array2mb_6_flag_v; // @[TLB.scala 98:31]
  reg [8:0] array2mb_6_vpn2; // @[TLB.scala 98:31]
  reg [8:0] array2mb_6_vpn1; // @[TLB.scala 98:31]
  reg [1:0] array2mb_6_ppn2; // @[TLB.scala 98:31]
  reg [8:0] array2mb_6_ppn1; // @[TLB.scala 98:31]
  reg [15:0] array2mb_6_asid; // @[TLB.scala 98:31]
  reg  array2mb_7_flag_d; // @[TLB.scala 98:31]
  reg  array2mb_7_flag_a; // @[TLB.scala 98:31]
  reg  array2mb_7_flag_g; // @[TLB.scala 98:31]
  reg  array2mb_7_flag_u; // @[TLB.scala 98:31]
  reg  array2mb_7_flag_x; // @[TLB.scala 98:31]
  reg  array2mb_7_flag_w; // @[TLB.scala 98:31]
  reg  array2mb_7_flag_r; // @[TLB.scala 98:31]
  reg  array2mb_7_flag_v; // @[TLB.scala 98:31]
  reg [8:0] array2mb_7_vpn2; // @[TLB.scala 98:31]
  reg [8:0] array2mb_7_vpn1; // @[TLB.scala 98:31]
  reg [1:0] array2mb_7_ppn2; // @[TLB.scala 98:31]
  reg [8:0] array2mb_7_ppn1; // @[TLB.scala 98:31]
  reg [15:0] array2mb_7_asid; // @[TLB.scala 98:31]
  reg  array2mb_valid_0; // @[TLB.scala 99:31]
  reg  array2mb_valid_1; // @[TLB.scala 99:31]
  reg  array2mb_valid_2; // @[TLB.scala 99:31]
  reg  array2mb_valid_3; // @[TLB.scala 99:31]
  reg  array2mb_valid_4; // @[TLB.scala 99:31]
  reg  array2mb_valid_5; // @[TLB.scala 99:31]
  reg  array2mb_valid_6; // @[TLB.scala 99:31]
  reg  array2mb_valid_7; // @[TLB.scala 99:31]
  wire [17:0] _T_138 = {array2mb_0_vpn2,array2mb_0_vpn1}; // @[Cat.scala 33:92]
  wire  _GEN_1664 = array2mb_valid_0 & _T_138 == hi_1 & (array2mb_0_asid == io_satp_asid | array2mb_0_flag_g); // @[TLB.scala 105:77 106:22 102:35]
  wire  _GEN_1666 = array2mb_valid_0 & _T_138 == hi_1 & array2mb_0_flag_d; // @[TLB.scala 105:77 107:22 100:35]
  wire  _GEN_1667 = array2mb_valid_0 & _T_138 == hi_1 & array2mb_0_flag_a; // @[TLB.scala 105:77 107:22 100:35]
  wire  _GEN_1669 = array2mb_valid_0 & _T_138 == hi_1 & array2mb_0_flag_u; // @[TLB.scala 105:77 107:22 100:35]
  wire  _GEN_1670 = array2mb_valid_0 & _T_138 == hi_1 & array2mb_0_flag_x; // @[TLB.scala 105:77 107:22 100:35]
  wire  _GEN_1671 = array2mb_valid_0 & _T_138 == hi_1 & array2mb_0_flag_w; // @[TLB.scala 105:77 107:22 100:35]
  wire  _GEN_1672 = array2mb_valid_0 & _T_138 == hi_1 & array2mb_0_flag_r; // @[TLB.scala 105:77 107:22 100:35]
  wire  _GEN_1673 = array2mb_valid_0 & _T_138 == hi_1 & array2mb_0_flag_v; // @[TLB.scala 105:77 107:22 100:35]
  wire [1:0] _GEN_1676 = array2mb_valid_0 & _T_138 == hi_1 ? array2mb_0_ppn2 : 2'h0; // @[TLB.scala 105:77 107:22 100:35]
  wire [8:0] _GEN_1677 = array2mb_valid_0 & _T_138 == hi_1 ? array2mb_0_ppn1 : 9'h0; // @[TLB.scala 105:77 107:22 100:35]
  wire [17:0] _T_142 = {array2mb_1_vpn2,array2mb_1_vpn1}; // @[Cat.scala 33:92]
  wire  _GEN_1679 = array2mb_valid_1 & _T_142 == hi_1 ? array2mb_1_asid == io_satp_asid | array2mb_1_flag_g : _GEN_1664; // @[TLB.scala 105:77 106:22]
  wire  _GEN_1681 = array2mb_valid_1 & _T_142 == hi_1 ? array2mb_1_flag_d : _GEN_1666; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1682 = array2mb_valid_1 & _T_142 == hi_1 ? array2mb_1_flag_a : _GEN_1667; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1684 = array2mb_valid_1 & _T_142 == hi_1 ? array2mb_1_flag_u : _GEN_1669; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1685 = array2mb_valid_1 & _T_142 == hi_1 ? array2mb_1_flag_x : _GEN_1670; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1686 = array2mb_valid_1 & _T_142 == hi_1 ? array2mb_1_flag_w : _GEN_1671; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1687 = array2mb_valid_1 & _T_142 == hi_1 ? array2mb_1_flag_r : _GEN_1672; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1688 = array2mb_valid_1 & _T_142 == hi_1 ? array2mb_1_flag_v : _GEN_1673; // @[TLB.scala 105:77 107:22]
  wire [1:0] _GEN_1691 = array2mb_valid_1 & _T_142 == hi_1 ? array2mb_1_ppn2 : _GEN_1676; // @[TLB.scala 105:77 107:22]
  wire [8:0] _GEN_1692 = array2mb_valid_1 & _T_142 == hi_1 ? array2mb_1_ppn1 : _GEN_1677; // @[TLB.scala 105:77 107:22]
  wire [17:0] _T_146 = {array2mb_2_vpn2,array2mb_2_vpn1}; // @[Cat.scala 33:92]
  wire  _GEN_1694 = array2mb_valid_2 & _T_146 == hi_1 ? array2mb_2_asid == io_satp_asid | array2mb_2_flag_g : _GEN_1679; // @[TLB.scala 105:77 106:22]
  wire  _GEN_1696 = array2mb_valid_2 & _T_146 == hi_1 ? array2mb_2_flag_d : _GEN_1681; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1697 = array2mb_valid_2 & _T_146 == hi_1 ? array2mb_2_flag_a : _GEN_1682; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1699 = array2mb_valid_2 & _T_146 == hi_1 ? array2mb_2_flag_u : _GEN_1684; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1700 = array2mb_valid_2 & _T_146 == hi_1 ? array2mb_2_flag_x : _GEN_1685; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1701 = array2mb_valid_2 & _T_146 == hi_1 ? array2mb_2_flag_w : _GEN_1686; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1702 = array2mb_valid_2 & _T_146 == hi_1 ? array2mb_2_flag_r : _GEN_1687; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1703 = array2mb_valid_2 & _T_146 == hi_1 ? array2mb_2_flag_v : _GEN_1688; // @[TLB.scala 105:77 107:22]
  wire [1:0] _GEN_1706 = array2mb_valid_2 & _T_146 == hi_1 ? array2mb_2_ppn2 : _GEN_1691; // @[TLB.scala 105:77 107:22]
  wire [8:0] _GEN_1707 = array2mb_valid_2 & _T_146 == hi_1 ? array2mb_2_ppn1 : _GEN_1692; // @[TLB.scala 105:77 107:22]
  wire [17:0] _T_150 = {array2mb_3_vpn2,array2mb_3_vpn1}; // @[Cat.scala 33:92]
  wire  _GEN_1709 = array2mb_valid_3 & _T_150 == hi_1 ? array2mb_3_asid == io_satp_asid | array2mb_3_flag_g : _GEN_1694; // @[TLB.scala 105:77 106:22]
  wire  _GEN_1711 = array2mb_valid_3 & _T_150 == hi_1 ? array2mb_3_flag_d : _GEN_1696; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1712 = array2mb_valid_3 & _T_150 == hi_1 ? array2mb_3_flag_a : _GEN_1697; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1714 = array2mb_valid_3 & _T_150 == hi_1 ? array2mb_3_flag_u : _GEN_1699; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1715 = array2mb_valid_3 & _T_150 == hi_1 ? array2mb_3_flag_x : _GEN_1700; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1716 = array2mb_valid_3 & _T_150 == hi_1 ? array2mb_3_flag_w : _GEN_1701; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1717 = array2mb_valid_3 & _T_150 == hi_1 ? array2mb_3_flag_r : _GEN_1702; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1718 = array2mb_valid_3 & _T_150 == hi_1 ? array2mb_3_flag_v : _GEN_1703; // @[TLB.scala 105:77 107:22]
  wire [1:0] _GEN_1721 = array2mb_valid_3 & _T_150 == hi_1 ? array2mb_3_ppn2 : _GEN_1706; // @[TLB.scala 105:77 107:22]
  wire [8:0] _GEN_1722 = array2mb_valid_3 & _T_150 == hi_1 ? array2mb_3_ppn1 : _GEN_1707; // @[TLB.scala 105:77 107:22]
  wire [17:0] _T_154 = {array2mb_4_vpn2,array2mb_4_vpn1}; // @[Cat.scala 33:92]
  wire  _GEN_1724 = array2mb_valid_4 & _T_154 == hi_1 ? array2mb_4_asid == io_satp_asid | array2mb_4_flag_g : _GEN_1709; // @[TLB.scala 105:77 106:22]
  wire  _GEN_1726 = array2mb_valid_4 & _T_154 == hi_1 ? array2mb_4_flag_d : _GEN_1711; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1727 = array2mb_valid_4 & _T_154 == hi_1 ? array2mb_4_flag_a : _GEN_1712; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1729 = array2mb_valid_4 & _T_154 == hi_1 ? array2mb_4_flag_u : _GEN_1714; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1730 = array2mb_valid_4 & _T_154 == hi_1 ? array2mb_4_flag_x : _GEN_1715; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1731 = array2mb_valid_4 & _T_154 == hi_1 ? array2mb_4_flag_w : _GEN_1716; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1732 = array2mb_valid_4 & _T_154 == hi_1 ? array2mb_4_flag_r : _GEN_1717; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1733 = array2mb_valid_4 & _T_154 == hi_1 ? array2mb_4_flag_v : _GEN_1718; // @[TLB.scala 105:77 107:22]
  wire [1:0] _GEN_1736 = array2mb_valid_4 & _T_154 == hi_1 ? array2mb_4_ppn2 : _GEN_1721; // @[TLB.scala 105:77 107:22]
  wire [8:0] _GEN_1737 = array2mb_valid_4 & _T_154 == hi_1 ? array2mb_4_ppn1 : _GEN_1722; // @[TLB.scala 105:77 107:22]
  wire [17:0] _T_158 = {array2mb_5_vpn2,array2mb_5_vpn1}; // @[Cat.scala 33:92]
  wire  _GEN_1739 = array2mb_valid_5 & _T_158 == hi_1 ? array2mb_5_asid == io_satp_asid | array2mb_5_flag_g : _GEN_1724; // @[TLB.scala 105:77 106:22]
  wire  _GEN_1741 = array2mb_valid_5 & _T_158 == hi_1 ? array2mb_5_flag_d : _GEN_1726; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1742 = array2mb_valid_5 & _T_158 == hi_1 ? array2mb_5_flag_a : _GEN_1727; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1744 = array2mb_valid_5 & _T_158 == hi_1 ? array2mb_5_flag_u : _GEN_1729; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1745 = array2mb_valid_5 & _T_158 == hi_1 ? array2mb_5_flag_x : _GEN_1730; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1746 = array2mb_valid_5 & _T_158 == hi_1 ? array2mb_5_flag_w : _GEN_1731; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1747 = array2mb_valid_5 & _T_158 == hi_1 ? array2mb_5_flag_r : _GEN_1732; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1748 = array2mb_valid_5 & _T_158 == hi_1 ? array2mb_5_flag_v : _GEN_1733; // @[TLB.scala 105:77 107:22]
  wire [1:0] _GEN_1751 = array2mb_valid_5 & _T_158 == hi_1 ? array2mb_5_ppn2 : _GEN_1736; // @[TLB.scala 105:77 107:22]
  wire [8:0] _GEN_1752 = array2mb_valid_5 & _T_158 == hi_1 ? array2mb_5_ppn1 : _GEN_1737; // @[TLB.scala 105:77 107:22]
  wire [17:0] _T_162 = {array2mb_6_vpn2,array2mb_6_vpn1}; // @[Cat.scala 33:92]
  wire  _GEN_1754 = array2mb_valid_6 & _T_162 == hi_1 ? array2mb_6_asid == io_satp_asid | array2mb_6_flag_g : _GEN_1739; // @[TLB.scala 105:77 106:22]
  wire  _GEN_1756 = array2mb_valid_6 & _T_162 == hi_1 ? array2mb_6_flag_d : _GEN_1741; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1757 = array2mb_valid_6 & _T_162 == hi_1 ? array2mb_6_flag_a : _GEN_1742; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1759 = array2mb_valid_6 & _T_162 == hi_1 ? array2mb_6_flag_u : _GEN_1744; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1760 = array2mb_valid_6 & _T_162 == hi_1 ? array2mb_6_flag_x : _GEN_1745; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1761 = array2mb_valid_6 & _T_162 == hi_1 ? array2mb_6_flag_w : _GEN_1746; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1762 = array2mb_valid_6 & _T_162 == hi_1 ? array2mb_6_flag_r : _GEN_1747; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1763 = array2mb_valid_6 & _T_162 == hi_1 ? array2mb_6_flag_v : _GEN_1748; // @[TLB.scala 105:77 107:22]
  wire [1:0] _GEN_1766 = array2mb_valid_6 & _T_162 == hi_1 ? array2mb_6_ppn2 : _GEN_1751; // @[TLB.scala 105:77 107:22]
  wire [8:0] _GEN_1767 = array2mb_valid_6 & _T_162 == hi_1 ? array2mb_6_ppn1 : _GEN_1752; // @[TLB.scala 105:77 107:22]
  wire [17:0] _T_166 = {array2mb_7_vpn2,array2mb_7_vpn1}; // @[Cat.scala 33:92]
  wire  hit2mb = array2mb_valid_7 & _T_166 == hi_1 ? array2mb_7_asid == io_satp_asid | array2mb_7_flag_g : _GEN_1754; // @[TLB.scala 105:77 106:22]
  wire  array2mb_rdata_flag_d = array2mb_valid_7 & _T_166 == hi_1 ? array2mb_7_flag_d : _GEN_1756; // @[TLB.scala 105:77 107:22]
  wire  array2mb_rdata_flag_a = array2mb_valid_7 & _T_166 == hi_1 ? array2mb_7_flag_a : _GEN_1757; // @[TLB.scala 105:77 107:22]
  wire  array2mb_rdata_flag_u = array2mb_valid_7 & _T_166 == hi_1 ? array2mb_7_flag_u : _GEN_1759; // @[TLB.scala 105:77 107:22]
  wire  array2mb_rdata_flag_x = array2mb_valid_7 & _T_166 == hi_1 ? array2mb_7_flag_x : _GEN_1760; // @[TLB.scala 105:77 107:22]
  wire  array2mb_rdata_flag_w = array2mb_valid_7 & _T_166 == hi_1 ? array2mb_7_flag_w : _GEN_1761; // @[TLB.scala 105:77 107:22]
  wire  array2mb_rdata_flag_r = array2mb_valid_7 & _T_166 == hi_1 ? array2mb_7_flag_r : _GEN_1762; // @[TLB.scala 105:77 107:22]
  wire  array2mb_rdata_flag_v = array2mb_valid_7 & _T_166 == hi_1 ? array2mb_7_flag_v : _GEN_1763; // @[TLB.scala 105:77 107:22]
  wire [1:0] array2mb_rdata_ppn2 = array2mb_valid_7 & _T_166 == hi_1 ? array2mb_7_ppn2 : _GEN_1766; // @[TLB.scala 105:77 107:22]
  wire [8:0] array2mb_rdata_ppn1 = array2mb_valid_7 & _T_166 == hi_1 ? array2mb_7_ppn1 : _GEN_1767; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1896 = 3'h0 == replace_idx[2:0] | array2mb_valid_0; // @[TLB.scala 119:{33,33} 99:31]
  wire  _GEN_1897 = 3'h1 == replace_idx[2:0] | array2mb_valid_1; // @[TLB.scala 119:{33,33} 99:31]
  wire  _GEN_1898 = 3'h2 == replace_idx[2:0] | array2mb_valid_2; // @[TLB.scala 119:{33,33} 99:31]
  wire  _GEN_1899 = 3'h3 == replace_idx[2:0] | array2mb_valid_3; // @[TLB.scala 119:{33,33} 99:31]
  wire  _GEN_1900 = 3'h4 == replace_idx[2:0] | array2mb_valid_4; // @[TLB.scala 119:{33,33} 99:31]
  wire  _GEN_1901 = 3'h5 == replace_idx[2:0] | array2mb_valid_5; // @[TLB.scala 119:{33,33} 99:31]
  wire  _GEN_1902 = 3'h6 == replace_idx[2:0] | array2mb_valid_6; // @[TLB.scala 119:{33,33} 99:31]
  wire  _GEN_1903 = 3'h7 == replace_idx[2:0] | array2mb_valid_7; // @[TLB.scala 119:{33,33} 99:31]
  reg  array1gb_0_flag_d; // @[TLB.scala 130:31]
  reg  array1gb_0_flag_a; // @[TLB.scala 130:31]
  reg  array1gb_0_flag_g; // @[TLB.scala 130:31]
  reg  array1gb_0_flag_u; // @[TLB.scala 130:31]
  reg  array1gb_0_flag_x; // @[TLB.scala 130:31]
  reg  array1gb_0_flag_w; // @[TLB.scala 130:31]
  reg  array1gb_0_flag_r; // @[TLB.scala 130:31]
  reg  array1gb_0_flag_v; // @[TLB.scala 130:31]
  reg [8:0] array1gb_0_vpn2; // @[TLB.scala 130:31]
  reg [1:0] array1gb_0_ppn2; // @[TLB.scala 130:31]
  reg [15:0] array1gb_0_asid; // @[TLB.scala 130:31]
  reg  array1gb_1_flag_d; // @[TLB.scala 130:31]
  reg  array1gb_1_flag_a; // @[TLB.scala 130:31]
  reg  array1gb_1_flag_g; // @[TLB.scala 130:31]
  reg  array1gb_1_flag_u; // @[TLB.scala 130:31]
  reg  array1gb_1_flag_x; // @[TLB.scala 130:31]
  reg  array1gb_1_flag_w; // @[TLB.scala 130:31]
  reg  array1gb_1_flag_r; // @[TLB.scala 130:31]
  reg  array1gb_1_flag_v; // @[TLB.scala 130:31]
  reg [8:0] array1gb_1_vpn2; // @[TLB.scala 130:31]
  reg [1:0] array1gb_1_ppn2; // @[TLB.scala 130:31]
  reg [15:0] array1gb_1_asid; // @[TLB.scala 130:31]
  reg  array1gb_2_flag_d; // @[TLB.scala 130:31]
  reg  array1gb_2_flag_a; // @[TLB.scala 130:31]
  reg  array1gb_2_flag_g; // @[TLB.scala 130:31]
  reg  array1gb_2_flag_u; // @[TLB.scala 130:31]
  reg  array1gb_2_flag_x; // @[TLB.scala 130:31]
  reg  array1gb_2_flag_w; // @[TLB.scala 130:31]
  reg  array1gb_2_flag_r; // @[TLB.scala 130:31]
  reg  array1gb_2_flag_v; // @[TLB.scala 130:31]
  reg [8:0] array1gb_2_vpn2; // @[TLB.scala 130:31]
  reg [1:0] array1gb_2_ppn2; // @[TLB.scala 130:31]
  reg [15:0] array1gb_2_asid; // @[TLB.scala 130:31]
  reg  array1gb_3_flag_d; // @[TLB.scala 130:31]
  reg  array1gb_3_flag_a; // @[TLB.scala 130:31]
  reg  array1gb_3_flag_g; // @[TLB.scala 130:31]
  reg  array1gb_3_flag_u; // @[TLB.scala 130:31]
  reg  array1gb_3_flag_x; // @[TLB.scala 130:31]
  reg  array1gb_3_flag_w; // @[TLB.scala 130:31]
  reg  array1gb_3_flag_r; // @[TLB.scala 130:31]
  reg  array1gb_3_flag_v; // @[TLB.scala 130:31]
  reg [8:0] array1gb_3_vpn2; // @[TLB.scala 130:31]
  reg [1:0] array1gb_3_ppn2; // @[TLB.scala 130:31]
  reg [15:0] array1gb_3_asid; // @[TLB.scala 130:31]
  reg  array1gb_valid_0; // @[TLB.scala 131:31]
  reg  array1gb_valid_1; // @[TLB.scala 131:31]
  reg  array1gb_valid_2; // @[TLB.scala 131:31]
  reg  array1gb_valid_3; // @[TLB.scala 131:31]
  wire  _GEN_2032 = array1gb_valid_0 & array1gb_0_vpn2 == io_vaddr_vpn2 & (array1gb_0_asid == io_satp_asid |
    array1gb_0_flag_g); // @[TLB.scala 137:77 138:22 134:35]
  wire  _GEN_2034 = array1gb_valid_0 & array1gb_0_vpn2 == io_vaddr_vpn2 & array1gb_0_flag_d; // @[TLB.scala 137:77 139:22 132:35]
  wire  _GEN_2035 = array1gb_valid_0 & array1gb_0_vpn2 == io_vaddr_vpn2 & array1gb_0_flag_a; // @[TLB.scala 137:77 139:22 132:35]
  wire  _GEN_2037 = array1gb_valid_0 & array1gb_0_vpn2 == io_vaddr_vpn2 & array1gb_0_flag_u; // @[TLB.scala 137:77 139:22 132:35]
  wire  _GEN_2038 = array1gb_valid_0 & array1gb_0_vpn2 == io_vaddr_vpn2 & array1gb_0_flag_x; // @[TLB.scala 137:77 139:22 132:35]
  wire  _GEN_2039 = array1gb_valid_0 & array1gb_0_vpn2 == io_vaddr_vpn2 & array1gb_0_flag_w; // @[TLB.scala 137:77 139:22 132:35]
  wire  _GEN_2040 = array1gb_valid_0 & array1gb_0_vpn2 == io_vaddr_vpn2 & array1gb_0_flag_r; // @[TLB.scala 137:77 139:22 132:35]
  wire  _GEN_2041 = array1gb_valid_0 & array1gb_0_vpn2 == io_vaddr_vpn2 & array1gb_0_flag_v; // @[TLB.scala 137:77 139:22 132:35]
  wire [1:0] _GEN_2043 = array1gb_valid_0 & array1gb_0_vpn2 == io_vaddr_vpn2 ? array1gb_0_ppn2 : 2'h0; // @[TLB.scala 137:77 139:22 132:35]
  wire  _GEN_2045 = array1gb_valid_1 & array1gb_1_vpn2 == io_vaddr_vpn2 ? array1gb_1_asid == io_satp_asid |
    array1gb_1_flag_g : _GEN_2032; // @[TLB.scala 137:77 138:22]
  wire  _GEN_2047 = array1gb_valid_1 & array1gb_1_vpn2 == io_vaddr_vpn2 ? array1gb_1_flag_d : _GEN_2034; // @[TLB.scala 137:77 139:22]
  wire  _GEN_2048 = array1gb_valid_1 & array1gb_1_vpn2 == io_vaddr_vpn2 ? array1gb_1_flag_a : _GEN_2035; // @[TLB.scala 137:77 139:22]
  wire  _GEN_2050 = array1gb_valid_1 & array1gb_1_vpn2 == io_vaddr_vpn2 ? array1gb_1_flag_u : _GEN_2037; // @[TLB.scala 137:77 139:22]
  wire  _GEN_2051 = array1gb_valid_1 & array1gb_1_vpn2 == io_vaddr_vpn2 ? array1gb_1_flag_x : _GEN_2038; // @[TLB.scala 137:77 139:22]
  wire  _GEN_2052 = array1gb_valid_1 & array1gb_1_vpn2 == io_vaddr_vpn2 ? array1gb_1_flag_w : _GEN_2039; // @[TLB.scala 137:77 139:22]
  wire  _GEN_2053 = array1gb_valid_1 & array1gb_1_vpn2 == io_vaddr_vpn2 ? array1gb_1_flag_r : _GEN_2040; // @[TLB.scala 137:77 139:22]
  wire  _GEN_2054 = array1gb_valid_1 & array1gb_1_vpn2 == io_vaddr_vpn2 ? array1gb_1_flag_v : _GEN_2041; // @[TLB.scala 137:77 139:22]
  wire [1:0] _GEN_2056 = array1gb_valid_1 & array1gb_1_vpn2 == io_vaddr_vpn2 ? array1gb_1_ppn2 : _GEN_2043; // @[TLB.scala 137:77 139:22]
  wire  _GEN_2058 = array1gb_valid_2 & array1gb_2_vpn2 == io_vaddr_vpn2 ? array1gb_2_asid == io_satp_asid |
    array1gb_2_flag_g : _GEN_2045; // @[TLB.scala 137:77 138:22]
  wire  _GEN_2060 = array1gb_valid_2 & array1gb_2_vpn2 == io_vaddr_vpn2 ? array1gb_2_flag_d : _GEN_2047; // @[TLB.scala 137:77 139:22]
  wire  _GEN_2061 = array1gb_valid_2 & array1gb_2_vpn2 == io_vaddr_vpn2 ? array1gb_2_flag_a : _GEN_2048; // @[TLB.scala 137:77 139:22]
  wire  _GEN_2063 = array1gb_valid_2 & array1gb_2_vpn2 == io_vaddr_vpn2 ? array1gb_2_flag_u : _GEN_2050; // @[TLB.scala 137:77 139:22]
  wire  _GEN_2064 = array1gb_valid_2 & array1gb_2_vpn2 == io_vaddr_vpn2 ? array1gb_2_flag_x : _GEN_2051; // @[TLB.scala 137:77 139:22]
  wire  _GEN_2065 = array1gb_valid_2 & array1gb_2_vpn2 == io_vaddr_vpn2 ? array1gb_2_flag_w : _GEN_2052; // @[TLB.scala 137:77 139:22]
  wire  _GEN_2066 = array1gb_valid_2 & array1gb_2_vpn2 == io_vaddr_vpn2 ? array1gb_2_flag_r : _GEN_2053; // @[TLB.scala 137:77 139:22]
  wire  _GEN_2067 = array1gb_valid_2 & array1gb_2_vpn2 == io_vaddr_vpn2 ? array1gb_2_flag_v : _GEN_2054; // @[TLB.scala 137:77 139:22]
  wire [1:0] _GEN_2069 = array1gb_valid_2 & array1gb_2_vpn2 == io_vaddr_vpn2 ? array1gb_2_ppn2 : _GEN_2056; // @[TLB.scala 137:77 139:22]
  wire  hit1gb = array1gb_valid_3 & array1gb_3_vpn2 == io_vaddr_vpn2 ? array1gb_3_asid == io_satp_asid |
    array1gb_3_flag_g : _GEN_2058; // @[TLB.scala 137:77 138:22]
  wire  array1gb_rdata_flag_d = array1gb_valid_3 & array1gb_3_vpn2 == io_vaddr_vpn2 ? array1gb_3_flag_d : _GEN_2060; // @[TLB.scala 137:77 139:22]
  wire  array1gb_rdata_flag_a = array1gb_valid_3 & array1gb_3_vpn2 == io_vaddr_vpn2 ? array1gb_3_flag_a : _GEN_2061; // @[TLB.scala 137:77 139:22]
  wire  array1gb_rdata_flag_u = array1gb_valid_3 & array1gb_3_vpn2 == io_vaddr_vpn2 ? array1gb_3_flag_u : _GEN_2063; // @[TLB.scala 137:77 139:22]
  wire  array1gb_rdata_flag_x = array1gb_valid_3 & array1gb_3_vpn2 == io_vaddr_vpn2 ? array1gb_3_flag_x : _GEN_2064; // @[TLB.scala 137:77 139:22]
  wire  array1gb_rdata_flag_w = array1gb_valid_3 & array1gb_3_vpn2 == io_vaddr_vpn2 ? array1gb_3_flag_w : _GEN_2065; // @[TLB.scala 137:77 139:22]
  wire  array1gb_rdata_flag_r = array1gb_valid_3 & array1gb_3_vpn2 == io_vaddr_vpn2 ? array1gb_3_flag_r : _GEN_2066; // @[TLB.scala 137:77 139:22]
  wire  array1gb_rdata_flag_v = array1gb_valid_3 & array1gb_3_vpn2 == io_vaddr_vpn2 ? array1gb_3_flag_v : _GEN_2067; // @[TLB.scala 137:77 139:22]
  wire [1:0] array1gb_rdata_ppn2 = array1gb_valid_3 & array1gb_3_vpn2 == io_vaddr_vpn2 ? array1gb_3_ppn2 : _GEN_2069; // @[TLB.scala 137:77 139:22]
  wire  _GEN_2132 = 2'h0 == replace_idx[1:0] | array1gb_valid_0; // @[TLB.scala 131:31 149:{33,33}]
  wire  _GEN_2133 = 2'h1 == replace_idx[1:0] | array1gb_valid_1; // @[TLB.scala 131:31 149:{33,33}]
  wire  _GEN_2134 = 2'h2 == replace_idx[1:0] | array1gb_valid_2; // @[TLB.scala 131:31 149:{33,33}]
  wire  _GEN_2135 = 2'h3 == replace_idx[1:0] | array1gb_valid_3; // @[TLB.scala 131:31 149:{33,33}]
  wire  _GEN_2193 = hit1gb & array1gb_rdata_flag_d; // @[TLB.scala 158:13 172:22 173:18]
  wire  _GEN_2194 = hit1gb & array1gb_rdata_flag_a; // @[TLB.scala 158:13 172:22 173:18]
  wire  _GEN_2196 = hit1gb & array1gb_rdata_flag_u; // @[TLB.scala 158:13 172:22 173:18]
  wire  _GEN_2197 = hit1gb & array1gb_rdata_flag_x; // @[TLB.scala 158:13 172:22 173:18]
  wire  _GEN_2198 = hit1gb & array1gb_rdata_flag_w; // @[TLB.scala 158:13 172:22 173:18]
  wire  _GEN_2199 = hit1gb & array1gb_rdata_flag_r; // @[TLB.scala 158:13 172:22 173:18]
  wire  _GEN_2200 = hit1gb & array1gb_rdata_flag_v; // @[TLB.scala 158:13 172:22 173:18]
  wire [1:0] _GEN_2203 = hit1gb ? array1gb_rdata_ppn2 : 2'h0; // @[TLB.scala 158:13 172:22 176:18]
  wire [1:0] _GEN_2204 = hit1gb ? 2'h2 : 2'h0; // @[TLB.scala 159:13 172:22 177:18]
  wire  _GEN_2206 = hit2mb ? array2mb_rdata_flag_d : _GEN_2193; // @[TLB.scala 166:22 167:18]
  wire  _GEN_2207 = hit2mb ? array2mb_rdata_flag_a : _GEN_2194; // @[TLB.scala 166:22 167:18]
  wire  _GEN_2209 = hit2mb ? array2mb_rdata_flag_u : _GEN_2196; // @[TLB.scala 166:22 167:18]
  wire  _GEN_2210 = hit2mb ? array2mb_rdata_flag_x : _GEN_2197; // @[TLB.scala 166:22 167:18]
  wire  _GEN_2211 = hit2mb ? array2mb_rdata_flag_w : _GEN_2198; // @[TLB.scala 166:22 167:18]
  wire  _GEN_2212 = hit2mb ? array2mb_rdata_flag_r : _GEN_2199; // @[TLB.scala 166:22 167:18]
  wire  _GEN_2213 = hit2mb ? array2mb_rdata_flag_v : _GEN_2200; // @[TLB.scala 166:22 167:18]
  wire [8:0] _GEN_2215 = hit2mb ? array2mb_rdata_ppn1 : 9'h0; // @[TLB.scala 166:22 169:18]
  wire [1:0] _GEN_2216 = hit2mb ? array2mb_rdata_ppn2 : _GEN_2203; // @[TLB.scala 166:22 170:18]
  wire [1:0] _GEN_2217 = hit2mb ? 2'h1 : _GEN_2204; // @[TLB.scala 166:22 171:18]
  MaxPeriodFibonacciLFSR_1 replace_idx_prng ( // @[PRNG.scala 91:22]
    .clock(replace_idx_prng_clock),
    .reset(replace_idx_prng_reset),
    .io_out_0(replace_idx_prng_io_out_0),
    .io_out_1(replace_idx_prng_io_out_1),
    .io_out_2(replace_idx_prng_io_out_2),
    .io_out_3(replace_idx_prng_io_out_3),
    .io_out_4(replace_idx_prng_io_out_4)
  );
  assign io_rpte_ppn2 = hit4kb ? array4kb_rdata_ppn2 : _GEN_2216; // @[TLB.scala 161:16 165:18]
  assign io_rpte_ppn1 = hit4kb ? array4kb_rdata_ppn1 : _GEN_2215; // @[TLB.scala 161:16 164:18]
  assign io_rpte_ppn0 = hit4kb ? array4kb_rdata_ppn0 : 9'h0; // @[TLB.scala 161:16 163:18]
  assign io_rpte_flag_d = hit4kb ? array4kb_rdata_flag_d : _GEN_2206; // @[TLB.scala 161:16 162:18]
  assign io_rpte_flag_a = hit4kb ? array4kb_rdata_flag_a : _GEN_2207; // @[TLB.scala 161:16 162:18]
  assign io_rpte_flag_u = hit4kb ? array4kb_rdata_flag_u : _GEN_2209; // @[TLB.scala 161:16 162:18]
  assign io_rpte_flag_x = hit4kb ? array4kb_rdata_flag_x : _GEN_2210; // @[TLB.scala 161:16 162:18]
  assign io_rpte_flag_w = hit4kb ? array4kb_rdata_flag_w : _GEN_2211; // @[TLB.scala 161:16 162:18]
  assign io_rpte_flag_r = hit4kb ? array4kb_rdata_flag_r : _GEN_2212; // @[TLB.scala 161:16 162:18]
  assign io_rpte_flag_v = hit4kb ? array4kb_rdata_flag_v : _GEN_2213; // @[TLB.scala 161:16 162:18]
  assign io_rlevel = hit4kb ? 2'h0 : _GEN_2217; // @[TLB.scala 159:13 161:16]
  assign io_hit = hit4kb | hit2mb | hit1gb; // @[TLB.scala 160:33]
  assign replace_idx_prng_clock = clock;
  assign replace_idx_prng_reset = reset;
  always @(posedge clock) begin
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_0_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h0 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_0_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_0_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h0 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_0_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_0_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h0 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_0_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_0_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h0 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_0_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_0_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h0 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_0_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_0_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h0 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_0_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_0_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h0 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_0_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_0_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h0 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_0_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_0_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h0 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_0_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_0_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h0 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_0_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_0_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h0 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_0_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_0_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h0 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_0_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_0_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h0 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_0_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_0_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h0 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_0_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_0_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h0 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_0_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_1_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_1_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_1_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_1_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_1_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_1_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_1_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_1_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_1_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_1_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_1_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_1_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_1_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_1_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_1_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_1_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_1_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_1_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_1_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_1_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_1_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_1_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_1_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_1_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_1_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_1_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_1_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_1_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_1_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_1_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_2_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h2 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_2_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_2_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h2 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_2_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_2_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h2 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_2_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_2_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h2 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_2_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_2_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h2 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_2_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_2_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h2 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_2_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_2_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h2 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_2_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_2_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h2 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_2_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_2_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h2 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_2_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_2_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h2 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_2_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_2_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h2 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_2_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_2_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h2 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_2_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_2_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h2 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_2_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_2_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h2 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_2_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_2_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h2 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_2_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_3_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h3 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_3_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_3_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h3 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_3_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_3_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h3 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_3_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_3_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h3 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_3_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_3_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h3 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_3_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_3_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h3 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_3_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_3_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h3 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_3_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_3_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h3 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_3_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_3_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h3 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_3_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_3_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h3 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_3_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_3_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h3 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_3_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_3_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h3 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_3_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_3_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h3 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_3_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_3_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h3 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_3_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_3_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h3 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_3_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_4_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h4 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_4_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_4_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h4 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_4_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_4_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h4 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_4_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_4_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h4 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_4_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_4_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h4 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_4_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_4_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h4 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_4_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_4_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h4 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_4_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_4_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h4 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_4_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_4_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h4 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_4_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_4_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h4 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_4_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_4_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h4 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_4_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_4_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h4 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_4_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_4_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h4 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_4_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_4_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h4 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_4_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_4_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h4 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_4_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_5_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h5 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_5_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_5_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h5 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_5_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_5_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h5 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_5_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_5_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h5 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_5_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_5_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h5 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_5_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_5_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h5 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_5_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_5_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h5 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_5_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_5_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h5 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_5_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_5_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h5 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_5_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_5_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h5 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_5_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_5_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h5 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_5_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_5_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h5 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_5_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_5_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h5 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_5_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_5_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h5 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_5_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_5_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h5 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_5_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_6_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h6 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_6_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_6_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h6 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_6_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_6_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h6 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_6_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_6_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h6 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_6_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_6_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h6 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_6_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_6_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h6 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_6_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_6_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h6 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_6_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_6_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h6 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_6_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_6_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h6 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_6_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_6_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h6 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_6_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_6_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h6 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_6_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_6_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h6 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_6_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_6_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h6 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_6_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_6_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h6 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_6_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_6_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h6 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_6_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_7_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h7 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_7_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_7_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h7 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_7_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_7_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h7 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_7_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_7_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h7 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_7_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_7_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h7 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_7_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_7_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h7 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_7_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_7_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h7 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_7_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_7_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h7 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_7_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_7_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h7 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_7_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_7_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h7 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_7_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_7_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h7 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_7_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_7_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h7 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_7_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_7_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h7 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_7_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_7_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h7 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_7_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_7_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h7 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_7_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_8_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h8 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_8_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_8_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h8 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_8_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_8_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h8 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_8_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_8_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h8 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_8_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_8_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h8 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_8_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_8_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h8 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_8_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_8_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h8 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_8_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_8_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h8 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_8_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_8_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h8 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_8_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_8_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h8 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_8_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_8_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h8 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_8_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_8_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h8 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_8_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_8_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h8 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_8_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_8_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h8 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_8_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_8_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h8 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_8_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_9_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h9 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_9_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_9_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h9 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_9_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_9_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h9 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_9_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_9_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h9 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_9_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_9_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h9 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_9_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_9_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h9 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_9_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_9_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h9 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_9_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_9_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h9 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_9_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_9_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h9 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_9_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_9_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h9 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_9_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_9_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h9 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_9_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_9_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h9 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_9_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_9_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h9 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_9_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_9_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h9 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_9_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_9_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h9 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_9_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_10_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'ha == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_10_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_10_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'ha == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_10_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_10_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'ha == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_10_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_10_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'ha == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_10_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_10_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'ha == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_10_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_10_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'ha == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_10_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_10_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'ha == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_10_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_10_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'ha == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_10_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_10_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'ha == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_10_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_10_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'ha == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_10_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_10_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'ha == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_10_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_10_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'ha == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_10_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_10_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'ha == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_10_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_10_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'ha == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_10_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_10_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'ha == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_10_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_11_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hb == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_11_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_11_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hb == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_11_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_11_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hb == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_11_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_11_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hb == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_11_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_11_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hb == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_11_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_11_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hb == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_11_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_11_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hb == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_11_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_11_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hb == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_11_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_11_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hb == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_11_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_11_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hb == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_11_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_11_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hb == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_11_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_11_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hb == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_11_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_11_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hb == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_11_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_11_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hb == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_11_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_11_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hb == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_11_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_12_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hc == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_12_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_12_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hc == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_12_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_12_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hc == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_12_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_12_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hc == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_12_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_12_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hc == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_12_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_12_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hc == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_12_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_12_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hc == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_12_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_12_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hc == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_12_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_12_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hc == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_12_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_12_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hc == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_12_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_12_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hc == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_12_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_12_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hc == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_12_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_12_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hc == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_12_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_12_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hc == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_12_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_12_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hc == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_12_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_13_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hd == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_13_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_13_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hd == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_13_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_13_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hd == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_13_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_13_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hd == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_13_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_13_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hd == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_13_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_13_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hd == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_13_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_13_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hd == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_13_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_13_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hd == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_13_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_13_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hd == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_13_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_13_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hd == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_13_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_13_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hd == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_13_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_13_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hd == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_13_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_13_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hd == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_13_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_13_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hd == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_13_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_13_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hd == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_13_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_14_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'he == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_14_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_14_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'he == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_14_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_14_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'he == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_14_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_14_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'he == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_14_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_14_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'he == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_14_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_14_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'he == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_14_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_14_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'he == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_14_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_14_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'he == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_14_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_14_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'he == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_14_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_14_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'he == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_14_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_14_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'he == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_14_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_14_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'he == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_14_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_14_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'he == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_14_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_14_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'he == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_14_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_14_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'he == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_14_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_15_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hf == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_15_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_15_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hf == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_15_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_15_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hf == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_15_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_15_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hf == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_15_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_15_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hf == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_15_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_15_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hf == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_15_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_15_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hf == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_15_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_15_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hf == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_15_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_15_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hf == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_15_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_15_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hf == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_15_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_15_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hf == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_15_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_15_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hf == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_15_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_15_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hf == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_15_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_15_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hf == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_15_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_15_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hf == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_15_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_16_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h10 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_16_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_16_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h10 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_16_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_16_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h10 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_16_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_16_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h10 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_16_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_16_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h10 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_16_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_16_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h10 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_16_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_16_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h10 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_16_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_16_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h10 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_16_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_16_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h10 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_16_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_16_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h10 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_16_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_16_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h10 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_16_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_16_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h10 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_16_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_16_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h10 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_16_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_16_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h10 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_16_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_16_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h10 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_16_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_17_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h11 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_17_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_17_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h11 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_17_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_17_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h11 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_17_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_17_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h11 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_17_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_17_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h11 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_17_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_17_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h11 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_17_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_17_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h11 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_17_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_17_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h11 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_17_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_17_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h11 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_17_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_17_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h11 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_17_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_17_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h11 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_17_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_17_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h11 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_17_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_17_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h11 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_17_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_17_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h11 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_17_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_17_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h11 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_17_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_18_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h12 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_18_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_18_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h12 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_18_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_18_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h12 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_18_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_18_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h12 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_18_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_18_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h12 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_18_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_18_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h12 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_18_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_18_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h12 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_18_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_18_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h12 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_18_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_18_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h12 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_18_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_18_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h12 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_18_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_18_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h12 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_18_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_18_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h12 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_18_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_18_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h12 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_18_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_18_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h12 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_18_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_18_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h12 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_18_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_19_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h13 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_19_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_19_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h13 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_19_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_19_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h13 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_19_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_19_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h13 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_19_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_19_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h13 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_19_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_19_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h13 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_19_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_19_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h13 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_19_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_19_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h13 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_19_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_19_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h13 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_19_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_19_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h13 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_19_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_19_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h13 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_19_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_19_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h13 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_19_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_19_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h13 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_19_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_19_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h13 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_19_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_19_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h13 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_19_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_20_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h14 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_20_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_20_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h14 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_20_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_20_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h14 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_20_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_20_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h14 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_20_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_20_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h14 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_20_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_20_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h14 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_20_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_20_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h14 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_20_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_20_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h14 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_20_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_20_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h14 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_20_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_20_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h14 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_20_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_20_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h14 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_20_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_20_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h14 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_20_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_20_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h14 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_20_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_20_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h14 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_20_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_20_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h14 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_20_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_21_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h15 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_21_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_21_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h15 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_21_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_21_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h15 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_21_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_21_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h15 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_21_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_21_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h15 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_21_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_21_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h15 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_21_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_21_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h15 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_21_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_21_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h15 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_21_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_21_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h15 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_21_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_21_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h15 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_21_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_21_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h15 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_21_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_21_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h15 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_21_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_21_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h15 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_21_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_21_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h15 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_21_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_21_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h15 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_21_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_22_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h16 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_22_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_22_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h16 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_22_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_22_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h16 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_22_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_22_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h16 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_22_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_22_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h16 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_22_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_22_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h16 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_22_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_22_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h16 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_22_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_22_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h16 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_22_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_22_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h16 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_22_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_22_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h16 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_22_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_22_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h16 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_22_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_22_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h16 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_22_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_22_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h16 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_22_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_22_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h16 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_22_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_22_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h16 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_22_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_23_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h17 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_23_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_23_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h17 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_23_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_23_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h17 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_23_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_23_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h17 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_23_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_23_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h17 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_23_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_23_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h17 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_23_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_23_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h17 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_23_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_23_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h17 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_23_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_23_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h17 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_23_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_23_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h17 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_23_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_23_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h17 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_23_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_23_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h17 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_23_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_23_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h17 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_23_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_23_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h17 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_23_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_23_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h17 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_23_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_24_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h18 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_24_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_24_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h18 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_24_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_24_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h18 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_24_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_24_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h18 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_24_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_24_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h18 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_24_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_24_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h18 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_24_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_24_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h18 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_24_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_24_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h18 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_24_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_24_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h18 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_24_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_24_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h18 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_24_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_24_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h18 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_24_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_24_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h18 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_24_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_24_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h18 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_24_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_24_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h18 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_24_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_24_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h18 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_24_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_25_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h19 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_25_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_25_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h19 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_25_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_25_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h19 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_25_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_25_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h19 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_25_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_25_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h19 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_25_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_25_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h19 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_25_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_25_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h19 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_25_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_25_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h19 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_25_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_25_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h19 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_25_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_25_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h19 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_25_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_25_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h19 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_25_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_25_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h19 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_25_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_25_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h19 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_25_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_25_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h19 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_25_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_25_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h19 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_25_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_26_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1a == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_26_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_26_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1a == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_26_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_26_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1a == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_26_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_26_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1a == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_26_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_26_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1a == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_26_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_26_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1a == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_26_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_26_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1a == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_26_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_26_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1a == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_26_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_26_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1a == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_26_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_26_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1a == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_26_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_26_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1a == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_26_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_26_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1a == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_26_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_26_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1a == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_26_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_26_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1a == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_26_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_26_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1a == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_26_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_27_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1b == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_27_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_27_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1b == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_27_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_27_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1b == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_27_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_27_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1b == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_27_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_27_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1b == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_27_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_27_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1b == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_27_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_27_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1b == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_27_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_27_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1b == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_27_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_27_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1b == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_27_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_27_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1b == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_27_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_27_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1b == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_27_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_27_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1b == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_27_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_27_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1b == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_27_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_27_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1b == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_27_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_27_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1b == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_27_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_28_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1c == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_28_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_28_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1c == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_28_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_28_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1c == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_28_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_28_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1c == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_28_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_28_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1c == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_28_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_28_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1c == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_28_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_28_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1c == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_28_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_28_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1c == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_28_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_28_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1c == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_28_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_28_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1c == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_28_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_28_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1c == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_28_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_28_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1c == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_28_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_28_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1c == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_28_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_28_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1c == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_28_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_28_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1c == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_28_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_29_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1d == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_29_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_29_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1d == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_29_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_29_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1d == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_29_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_29_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1d == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_29_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_29_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1d == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_29_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_29_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1d == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_29_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_29_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1d == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_29_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_29_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1d == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_29_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_29_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1d == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_29_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_29_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1d == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_29_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_29_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1d == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_29_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_29_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1d == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_29_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_29_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1d == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_29_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_29_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1d == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_29_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_29_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1d == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_29_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_30_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1e == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_30_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_30_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1e == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_30_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_30_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1e == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_30_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_30_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1e == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_30_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_30_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1e == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_30_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_30_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1e == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_30_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_30_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1e == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_30_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_30_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1e == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_30_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_30_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1e == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_30_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_30_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1e == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_30_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_30_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1e == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_30_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_30_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1e == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_30_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_30_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1e == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_30_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_30_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1e == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_30_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_30_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1e == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_30_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_31_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1f == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_31_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_31_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1f == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_31_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_31_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1f == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_31_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_31_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1f == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_31_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_31_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1f == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_31_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_31_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1f == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_31_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_31_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1f == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_31_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_31_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1f == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_31_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_31_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1f == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_31_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_31_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1f == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_31_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_31_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1f == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_31_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_31_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1f == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_31_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_31_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1f == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_31_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_31_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1f == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_31_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_31_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1f == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_31_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_0 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_0 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_0 <= _GEN_1056;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_1 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_1 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_1 <= _GEN_1057;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_2 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_2 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_2 <= _GEN_1058;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_3 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_3 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_3 <= _GEN_1059;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_4 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_4 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_4 <= _GEN_1060;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_5 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_5 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_5 <= _GEN_1061;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_6 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_6 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_6 <= _GEN_1062;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_7 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_7 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_7 <= _GEN_1063;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_8 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_8 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_8 <= _GEN_1064;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_9 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_9 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_9 <= _GEN_1065;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_10 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_10 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_10 <= _GEN_1066;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_11 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_11 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_11 <= _GEN_1067;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_12 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_12 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_12 <= _GEN_1068;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_13 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_13 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_13 <= _GEN_1069;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_14 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_14 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_14 <= _GEN_1070;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_15 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_15 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_15 <= _GEN_1071;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_16 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_16 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_16 <= _GEN_1072;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_17 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_17 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_17 <= _GEN_1073;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_18 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_18 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_18 <= _GEN_1074;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_19 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_19 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_19 <= _GEN_1075;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_20 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_20 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_20 <= _GEN_1076;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_21 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_21 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_21 <= _GEN_1077;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_22 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_22 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_22 <= _GEN_1078;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_23 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_23 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_23 <= _GEN_1079;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_24 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_24 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_24 <= _GEN_1080;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_25 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_25 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_25 <= _GEN_1081;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_26 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_26 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_26 <= _GEN_1082;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_27 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_27 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_27 <= _GEN_1083;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_28 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_28 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_28 <= _GEN_1084;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_29 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_29 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_29 <= _GEN_1085;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_30 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_30 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_30 <= _GEN_1086;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_31 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_31 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_31 <= _GEN_1087;
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_0_flag_d <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h0 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_0_flag_d <= io_wpte_flag_d; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_0_flag_a <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h0 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_0_flag_a <= io_wpte_flag_a; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_0_flag_g <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h0 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_0_flag_g <= io_wpte_flag_g; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_0_flag_u <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h0 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_0_flag_u <= io_wpte_flag_u; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_0_flag_x <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h0 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_0_flag_x <= io_wpte_flag_x; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_0_flag_w <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h0 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_0_flag_w <= io_wpte_flag_w; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_0_flag_r <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h0 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_0_flag_r <= io_wpte_flag_r; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_0_flag_v <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h0 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_0_flag_v <= io_wpte_flag_v; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_0_vpn2 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h0 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_0_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_0_vpn1 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h0 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_0_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_0_ppn2 <= 2'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h0 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_0_ppn2 <= io_wpte_ppn2; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_0_ppn1 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h0 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_0_ppn1 <= io_wpte_ppn1; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_0_asid <= 16'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h0 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_0_asid <= io_satp_asid; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_1_flag_d <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h1 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_1_flag_d <= io_wpte_flag_d; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_1_flag_a <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h1 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_1_flag_a <= io_wpte_flag_a; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_1_flag_g <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h1 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_1_flag_g <= io_wpte_flag_g; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_1_flag_u <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h1 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_1_flag_u <= io_wpte_flag_u; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_1_flag_x <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h1 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_1_flag_x <= io_wpte_flag_x; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_1_flag_w <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h1 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_1_flag_w <= io_wpte_flag_w; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_1_flag_r <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h1 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_1_flag_r <= io_wpte_flag_r; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_1_flag_v <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h1 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_1_flag_v <= io_wpte_flag_v; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_1_vpn2 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h1 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_1_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_1_vpn1 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h1 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_1_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_1_ppn2 <= 2'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h1 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_1_ppn2 <= io_wpte_ppn2; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_1_ppn1 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h1 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_1_ppn1 <= io_wpte_ppn1; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_1_asid <= 16'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h1 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_1_asid <= io_satp_asid; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_2_flag_d <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h2 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_2_flag_d <= io_wpte_flag_d; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_2_flag_a <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h2 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_2_flag_a <= io_wpte_flag_a; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_2_flag_g <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h2 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_2_flag_g <= io_wpte_flag_g; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_2_flag_u <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h2 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_2_flag_u <= io_wpte_flag_u; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_2_flag_x <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h2 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_2_flag_x <= io_wpte_flag_x; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_2_flag_w <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h2 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_2_flag_w <= io_wpte_flag_w; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_2_flag_r <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h2 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_2_flag_r <= io_wpte_flag_r; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_2_flag_v <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h2 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_2_flag_v <= io_wpte_flag_v; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_2_vpn2 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h2 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_2_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_2_vpn1 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h2 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_2_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_2_ppn2 <= 2'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h2 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_2_ppn2 <= io_wpte_ppn2; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_2_ppn1 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h2 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_2_ppn1 <= io_wpte_ppn1; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_2_asid <= 16'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h2 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_2_asid <= io_satp_asid; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_3_flag_d <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h3 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_3_flag_d <= io_wpte_flag_d; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_3_flag_a <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h3 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_3_flag_a <= io_wpte_flag_a; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_3_flag_g <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h3 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_3_flag_g <= io_wpte_flag_g; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_3_flag_u <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h3 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_3_flag_u <= io_wpte_flag_u; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_3_flag_x <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h3 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_3_flag_x <= io_wpte_flag_x; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_3_flag_w <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h3 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_3_flag_w <= io_wpte_flag_w; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_3_flag_r <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h3 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_3_flag_r <= io_wpte_flag_r; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_3_flag_v <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h3 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_3_flag_v <= io_wpte_flag_v; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_3_vpn2 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h3 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_3_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_3_vpn1 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h3 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_3_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_3_ppn2 <= 2'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h3 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_3_ppn2 <= io_wpte_ppn2; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_3_ppn1 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h3 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_3_ppn1 <= io_wpte_ppn1; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_3_asid <= 16'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h3 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_3_asid <= io_satp_asid; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_4_flag_d <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h4 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_4_flag_d <= io_wpte_flag_d; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_4_flag_a <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h4 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_4_flag_a <= io_wpte_flag_a; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_4_flag_g <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h4 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_4_flag_g <= io_wpte_flag_g; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_4_flag_u <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h4 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_4_flag_u <= io_wpte_flag_u; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_4_flag_x <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h4 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_4_flag_x <= io_wpte_flag_x; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_4_flag_w <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h4 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_4_flag_w <= io_wpte_flag_w; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_4_flag_r <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h4 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_4_flag_r <= io_wpte_flag_r; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_4_flag_v <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h4 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_4_flag_v <= io_wpte_flag_v; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_4_vpn2 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h4 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_4_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_4_vpn1 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h4 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_4_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_4_ppn2 <= 2'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h4 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_4_ppn2 <= io_wpte_ppn2; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_4_ppn1 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h4 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_4_ppn1 <= io_wpte_ppn1; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_4_asid <= 16'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h4 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_4_asid <= io_satp_asid; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_5_flag_d <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h5 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_5_flag_d <= io_wpte_flag_d; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_5_flag_a <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h5 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_5_flag_a <= io_wpte_flag_a; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_5_flag_g <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h5 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_5_flag_g <= io_wpte_flag_g; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_5_flag_u <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h5 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_5_flag_u <= io_wpte_flag_u; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_5_flag_x <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h5 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_5_flag_x <= io_wpte_flag_x; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_5_flag_w <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h5 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_5_flag_w <= io_wpte_flag_w; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_5_flag_r <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h5 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_5_flag_r <= io_wpte_flag_r; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_5_flag_v <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h5 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_5_flag_v <= io_wpte_flag_v; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_5_vpn2 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h5 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_5_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_5_vpn1 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h5 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_5_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_5_ppn2 <= 2'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h5 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_5_ppn2 <= io_wpte_ppn2; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_5_ppn1 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h5 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_5_ppn1 <= io_wpte_ppn1; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_5_asid <= 16'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h5 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_5_asid <= io_satp_asid; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_6_flag_d <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h6 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_6_flag_d <= io_wpte_flag_d; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_6_flag_a <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h6 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_6_flag_a <= io_wpte_flag_a; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_6_flag_g <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h6 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_6_flag_g <= io_wpte_flag_g; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_6_flag_u <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h6 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_6_flag_u <= io_wpte_flag_u; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_6_flag_x <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h6 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_6_flag_x <= io_wpte_flag_x; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_6_flag_w <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h6 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_6_flag_w <= io_wpte_flag_w; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_6_flag_r <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h6 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_6_flag_r <= io_wpte_flag_r; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_6_flag_v <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h6 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_6_flag_v <= io_wpte_flag_v; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_6_vpn2 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h6 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_6_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_6_vpn1 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h6 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_6_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_6_ppn2 <= 2'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h6 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_6_ppn2 <= io_wpte_ppn2; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_6_ppn1 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h6 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_6_ppn1 <= io_wpte_ppn1; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_6_asid <= 16'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h6 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_6_asid <= io_satp_asid; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_7_flag_d <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h7 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_7_flag_d <= io_wpte_flag_d; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_7_flag_a <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h7 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_7_flag_a <= io_wpte_flag_a; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_7_flag_g <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h7 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_7_flag_g <= io_wpte_flag_g; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_7_flag_u <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h7 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_7_flag_u <= io_wpte_flag_u; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_7_flag_x <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h7 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_7_flag_x <= io_wpte_flag_x; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_7_flag_w <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h7 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_7_flag_w <= io_wpte_flag_w; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_7_flag_r <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h7 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_7_flag_r <= io_wpte_flag_r; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_7_flag_v <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h7 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_7_flag_v <= io_wpte_flag_v; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_7_vpn2 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h7 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_7_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_7_vpn1 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h7 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_7_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_7_ppn2 <= 2'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h7 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_7_ppn2 <= io_wpte_ppn2; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_7_ppn1 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h7 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_7_ppn1 <= io_wpte_ppn1; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_7_asid <= 16'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h7 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_7_asid <= io_satp_asid; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 99:31]
      array2mb_valid_0 <= 1'h0; // @[TLB.scala 99:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 121:23]
      array2mb_valid_0 <= 1'h0; // @[TLB.scala 123:25]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      array2mb_valid_0 <= _GEN_1896;
    end
    if (reset) begin // @[TLB.scala 99:31]
      array2mb_valid_1 <= 1'h0; // @[TLB.scala 99:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 121:23]
      array2mb_valid_1 <= 1'h0; // @[TLB.scala 123:25]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      array2mb_valid_1 <= _GEN_1897;
    end
    if (reset) begin // @[TLB.scala 99:31]
      array2mb_valid_2 <= 1'h0; // @[TLB.scala 99:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 121:23]
      array2mb_valid_2 <= 1'h0; // @[TLB.scala 123:25]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      array2mb_valid_2 <= _GEN_1898;
    end
    if (reset) begin // @[TLB.scala 99:31]
      array2mb_valid_3 <= 1'h0; // @[TLB.scala 99:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 121:23]
      array2mb_valid_3 <= 1'h0; // @[TLB.scala 123:25]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      array2mb_valid_3 <= _GEN_1899;
    end
    if (reset) begin // @[TLB.scala 99:31]
      array2mb_valid_4 <= 1'h0; // @[TLB.scala 99:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 121:23]
      array2mb_valid_4 <= 1'h0; // @[TLB.scala 123:25]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      array2mb_valid_4 <= _GEN_1900;
    end
    if (reset) begin // @[TLB.scala 99:31]
      array2mb_valid_5 <= 1'h0; // @[TLB.scala 99:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 121:23]
      array2mb_valid_5 <= 1'h0; // @[TLB.scala 123:25]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      array2mb_valid_5 <= _GEN_1901;
    end
    if (reset) begin // @[TLB.scala 99:31]
      array2mb_valid_6 <= 1'h0; // @[TLB.scala 99:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 121:23]
      array2mb_valid_6 <= 1'h0; // @[TLB.scala 123:25]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      array2mb_valid_6 <= _GEN_1902;
    end
    if (reset) begin // @[TLB.scala 99:31]
      array2mb_valid_7 <= 1'h0; // @[TLB.scala 99:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 121:23]
      array2mb_valid_7 <= 1'h0; // @[TLB.scala 123:25]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      array2mb_valid_7 <= _GEN_1903;
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_0_flag_d <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h0 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_0_flag_d <= io_wpte_flag_d; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_0_flag_a <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h0 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_0_flag_a <= io_wpte_flag_a; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_0_flag_g <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h0 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_0_flag_g <= io_wpte_flag_g; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_0_flag_u <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h0 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_0_flag_u <= io_wpte_flag_u; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_0_flag_x <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h0 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_0_flag_x <= io_wpte_flag_x; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_0_flag_w <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h0 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_0_flag_w <= io_wpte_flag_w; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_0_flag_r <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h0 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_0_flag_r <= io_wpte_flag_r; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_0_flag_v <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h0 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_0_flag_v <= io_wpte_flag_v; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_0_vpn2 <= 9'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h0 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_0_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_0_ppn2 <= 2'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h0 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_0_ppn2 <= io_wpte_ppn2; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_0_asid <= 16'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h0 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_0_asid <= io_satp_asid; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_1_flag_d <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h1 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_1_flag_d <= io_wpte_flag_d; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_1_flag_a <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h1 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_1_flag_a <= io_wpte_flag_a; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_1_flag_g <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h1 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_1_flag_g <= io_wpte_flag_g; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_1_flag_u <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h1 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_1_flag_u <= io_wpte_flag_u; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_1_flag_x <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h1 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_1_flag_x <= io_wpte_flag_x; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_1_flag_w <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h1 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_1_flag_w <= io_wpte_flag_w; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_1_flag_r <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h1 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_1_flag_r <= io_wpte_flag_r; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_1_flag_v <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h1 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_1_flag_v <= io_wpte_flag_v; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_1_vpn2 <= 9'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h1 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_1_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_1_ppn2 <= 2'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h1 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_1_ppn2 <= io_wpte_ppn2; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_1_asid <= 16'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h1 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_1_asid <= io_satp_asid; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_2_flag_d <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h2 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_2_flag_d <= io_wpte_flag_d; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_2_flag_a <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h2 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_2_flag_a <= io_wpte_flag_a; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_2_flag_g <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h2 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_2_flag_g <= io_wpte_flag_g; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_2_flag_u <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h2 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_2_flag_u <= io_wpte_flag_u; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_2_flag_x <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h2 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_2_flag_x <= io_wpte_flag_x; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_2_flag_w <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h2 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_2_flag_w <= io_wpte_flag_w; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_2_flag_r <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h2 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_2_flag_r <= io_wpte_flag_r; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_2_flag_v <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h2 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_2_flag_v <= io_wpte_flag_v; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_2_vpn2 <= 9'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h2 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_2_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_2_ppn2 <= 2'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h2 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_2_ppn2 <= io_wpte_ppn2; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_2_asid <= 16'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h2 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_2_asid <= io_satp_asid; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_3_flag_d <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h3 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_3_flag_d <= io_wpte_flag_d; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_3_flag_a <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h3 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_3_flag_a <= io_wpte_flag_a; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_3_flag_g <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h3 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_3_flag_g <= io_wpte_flag_g; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_3_flag_u <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h3 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_3_flag_u <= io_wpte_flag_u; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_3_flag_x <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h3 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_3_flag_x <= io_wpte_flag_x; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_3_flag_w <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h3 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_3_flag_w <= io_wpte_flag_w; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_3_flag_r <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h3 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_3_flag_r <= io_wpte_flag_r; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_3_flag_v <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h3 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_3_flag_v <= io_wpte_flag_v; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_3_vpn2 <= 9'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h3 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_3_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_3_ppn2 <= 2'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h3 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_3_ppn2 <= io_wpte_ppn2; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_3_asid <= 16'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h3 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_3_asid <= io_satp_asid; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 131:31]
      array1gb_valid_0 <= 1'h0; // @[TLB.scala 131:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 151:23]
      array1gb_valid_0 <= 1'h0; // @[TLB.scala 153:25]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      array1gb_valid_0 <= _GEN_2132;
    end
    if (reset) begin // @[TLB.scala 131:31]
      array1gb_valid_1 <= 1'h0; // @[TLB.scala 131:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 151:23]
      array1gb_valid_1 <= 1'h0; // @[TLB.scala 153:25]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      array1gb_valid_1 <= _GEN_2133;
    end
    if (reset) begin // @[TLB.scala 131:31]
      array1gb_valid_2 <= 1'h0; // @[TLB.scala 131:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 151:23]
      array1gb_valid_2 <= 1'h0; // @[TLB.scala 153:25]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      array1gb_valid_2 <= _GEN_2134;
    end
    if (reset) begin // @[TLB.scala 131:31]
      array1gb_valid_3 <= 1'h0; // @[TLB.scala 131:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 151:23]
      array1gb_valid_3 <= 1'h0; // @[TLB.scala 153:25]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      array1gb_valid_3 <= _GEN_2135;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_rlevel != 2'h3)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at TLB.scala:48 assert(io.rlevel =/= 3.U)\n"); // @[TLB.scala 48:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_rlevel != 2'h3)) begin
          $fatal; // @[TLB.scala 48:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(io_wlevel != 2'h3)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at TLB.scala:49 assert(io.wlevel =/= 3.U)\n"); // @[TLB.scala 49:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(io_wlevel != 2'h3)) begin
          $fatal; // @[TLB.scala 49:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  array4kb_0_flag_d = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  array4kb_0_flag_a = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  array4kb_0_flag_g = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  array4kb_0_flag_u = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  array4kb_0_flag_x = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  array4kb_0_flag_w = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  array4kb_0_flag_r = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  array4kb_0_flag_v = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  array4kb_0_vpn2 = _RAND_8[8:0];
  _RAND_9 = {1{`RANDOM}};
  array4kb_0_vpn1 = _RAND_9[8:0];
  _RAND_10 = {1{`RANDOM}};
  array4kb_0_vpn0 = _RAND_10[8:0];
  _RAND_11 = {1{`RANDOM}};
  array4kb_0_ppn2 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  array4kb_0_ppn1 = _RAND_12[8:0];
  _RAND_13 = {1{`RANDOM}};
  array4kb_0_ppn0 = _RAND_13[8:0];
  _RAND_14 = {1{`RANDOM}};
  array4kb_0_asid = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  array4kb_1_flag_d = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  array4kb_1_flag_a = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  array4kb_1_flag_g = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  array4kb_1_flag_u = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  array4kb_1_flag_x = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  array4kb_1_flag_w = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  array4kb_1_flag_r = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  array4kb_1_flag_v = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  array4kb_1_vpn2 = _RAND_23[8:0];
  _RAND_24 = {1{`RANDOM}};
  array4kb_1_vpn1 = _RAND_24[8:0];
  _RAND_25 = {1{`RANDOM}};
  array4kb_1_vpn0 = _RAND_25[8:0];
  _RAND_26 = {1{`RANDOM}};
  array4kb_1_ppn2 = _RAND_26[1:0];
  _RAND_27 = {1{`RANDOM}};
  array4kb_1_ppn1 = _RAND_27[8:0];
  _RAND_28 = {1{`RANDOM}};
  array4kb_1_ppn0 = _RAND_28[8:0];
  _RAND_29 = {1{`RANDOM}};
  array4kb_1_asid = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  array4kb_2_flag_d = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  array4kb_2_flag_a = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  array4kb_2_flag_g = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  array4kb_2_flag_u = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  array4kb_2_flag_x = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  array4kb_2_flag_w = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  array4kb_2_flag_r = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  array4kb_2_flag_v = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  array4kb_2_vpn2 = _RAND_38[8:0];
  _RAND_39 = {1{`RANDOM}};
  array4kb_2_vpn1 = _RAND_39[8:0];
  _RAND_40 = {1{`RANDOM}};
  array4kb_2_vpn0 = _RAND_40[8:0];
  _RAND_41 = {1{`RANDOM}};
  array4kb_2_ppn2 = _RAND_41[1:0];
  _RAND_42 = {1{`RANDOM}};
  array4kb_2_ppn1 = _RAND_42[8:0];
  _RAND_43 = {1{`RANDOM}};
  array4kb_2_ppn0 = _RAND_43[8:0];
  _RAND_44 = {1{`RANDOM}};
  array4kb_2_asid = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  array4kb_3_flag_d = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  array4kb_3_flag_a = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  array4kb_3_flag_g = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  array4kb_3_flag_u = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  array4kb_3_flag_x = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  array4kb_3_flag_w = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  array4kb_3_flag_r = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  array4kb_3_flag_v = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  array4kb_3_vpn2 = _RAND_53[8:0];
  _RAND_54 = {1{`RANDOM}};
  array4kb_3_vpn1 = _RAND_54[8:0];
  _RAND_55 = {1{`RANDOM}};
  array4kb_3_vpn0 = _RAND_55[8:0];
  _RAND_56 = {1{`RANDOM}};
  array4kb_3_ppn2 = _RAND_56[1:0];
  _RAND_57 = {1{`RANDOM}};
  array4kb_3_ppn1 = _RAND_57[8:0];
  _RAND_58 = {1{`RANDOM}};
  array4kb_3_ppn0 = _RAND_58[8:0];
  _RAND_59 = {1{`RANDOM}};
  array4kb_3_asid = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  array4kb_4_flag_d = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  array4kb_4_flag_a = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  array4kb_4_flag_g = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  array4kb_4_flag_u = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  array4kb_4_flag_x = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  array4kb_4_flag_w = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  array4kb_4_flag_r = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  array4kb_4_flag_v = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  array4kb_4_vpn2 = _RAND_68[8:0];
  _RAND_69 = {1{`RANDOM}};
  array4kb_4_vpn1 = _RAND_69[8:0];
  _RAND_70 = {1{`RANDOM}};
  array4kb_4_vpn0 = _RAND_70[8:0];
  _RAND_71 = {1{`RANDOM}};
  array4kb_4_ppn2 = _RAND_71[1:0];
  _RAND_72 = {1{`RANDOM}};
  array4kb_4_ppn1 = _RAND_72[8:0];
  _RAND_73 = {1{`RANDOM}};
  array4kb_4_ppn0 = _RAND_73[8:0];
  _RAND_74 = {1{`RANDOM}};
  array4kb_4_asid = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  array4kb_5_flag_d = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  array4kb_5_flag_a = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  array4kb_5_flag_g = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  array4kb_5_flag_u = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  array4kb_5_flag_x = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  array4kb_5_flag_w = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  array4kb_5_flag_r = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  array4kb_5_flag_v = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  array4kb_5_vpn2 = _RAND_83[8:0];
  _RAND_84 = {1{`RANDOM}};
  array4kb_5_vpn1 = _RAND_84[8:0];
  _RAND_85 = {1{`RANDOM}};
  array4kb_5_vpn0 = _RAND_85[8:0];
  _RAND_86 = {1{`RANDOM}};
  array4kb_5_ppn2 = _RAND_86[1:0];
  _RAND_87 = {1{`RANDOM}};
  array4kb_5_ppn1 = _RAND_87[8:0];
  _RAND_88 = {1{`RANDOM}};
  array4kb_5_ppn0 = _RAND_88[8:0];
  _RAND_89 = {1{`RANDOM}};
  array4kb_5_asid = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  array4kb_6_flag_d = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  array4kb_6_flag_a = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  array4kb_6_flag_g = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  array4kb_6_flag_u = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  array4kb_6_flag_x = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  array4kb_6_flag_w = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  array4kb_6_flag_r = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  array4kb_6_flag_v = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  array4kb_6_vpn2 = _RAND_98[8:0];
  _RAND_99 = {1{`RANDOM}};
  array4kb_6_vpn1 = _RAND_99[8:0];
  _RAND_100 = {1{`RANDOM}};
  array4kb_6_vpn0 = _RAND_100[8:0];
  _RAND_101 = {1{`RANDOM}};
  array4kb_6_ppn2 = _RAND_101[1:0];
  _RAND_102 = {1{`RANDOM}};
  array4kb_6_ppn1 = _RAND_102[8:0];
  _RAND_103 = {1{`RANDOM}};
  array4kb_6_ppn0 = _RAND_103[8:0];
  _RAND_104 = {1{`RANDOM}};
  array4kb_6_asid = _RAND_104[15:0];
  _RAND_105 = {1{`RANDOM}};
  array4kb_7_flag_d = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  array4kb_7_flag_a = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  array4kb_7_flag_g = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  array4kb_7_flag_u = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  array4kb_7_flag_x = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  array4kb_7_flag_w = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  array4kb_7_flag_r = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  array4kb_7_flag_v = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  array4kb_7_vpn2 = _RAND_113[8:0];
  _RAND_114 = {1{`RANDOM}};
  array4kb_7_vpn1 = _RAND_114[8:0];
  _RAND_115 = {1{`RANDOM}};
  array4kb_7_vpn0 = _RAND_115[8:0];
  _RAND_116 = {1{`RANDOM}};
  array4kb_7_ppn2 = _RAND_116[1:0];
  _RAND_117 = {1{`RANDOM}};
  array4kb_7_ppn1 = _RAND_117[8:0];
  _RAND_118 = {1{`RANDOM}};
  array4kb_7_ppn0 = _RAND_118[8:0];
  _RAND_119 = {1{`RANDOM}};
  array4kb_7_asid = _RAND_119[15:0];
  _RAND_120 = {1{`RANDOM}};
  array4kb_8_flag_d = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  array4kb_8_flag_a = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  array4kb_8_flag_g = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  array4kb_8_flag_u = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  array4kb_8_flag_x = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  array4kb_8_flag_w = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  array4kb_8_flag_r = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  array4kb_8_flag_v = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  array4kb_8_vpn2 = _RAND_128[8:0];
  _RAND_129 = {1{`RANDOM}};
  array4kb_8_vpn1 = _RAND_129[8:0];
  _RAND_130 = {1{`RANDOM}};
  array4kb_8_vpn0 = _RAND_130[8:0];
  _RAND_131 = {1{`RANDOM}};
  array4kb_8_ppn2 = _RAND_131[1:0];
  _RAND_132 = {1{`RANDOM}};
  array4kb_8_ppn1 = _RAND_132[8:0];
  _RAND_133 = {1{`RANDOM}};
  array4kb_8_ppn0 = _RAND_133[8:0];
  _RAND_134 = {1{`RANDOM}};
  array4kb_8_asid = _RAND_134[15:0];
  _RAND_135 = {1{`RANDOM}};
  array4kb_9_flag_d = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  array4kb_9_flag_a = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  array4kb_9_flag_g = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  array4kb_9_flag_u = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  array4kb_9_flag_x = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  array4kb_9_flag_w = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  array4kb_9_flag_r = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  array4kb_9_flag_v = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  array4kb_9_vpn2 = _RAND_143[8:0];
  _RAND_144 = {1{`RANDOM}};
  array4kb_9_vpn1 = _RAND_144[8:0];
  _RAND_145 = {1{`RANDOM}};
  array4kb_9_vpn0 = _RAND_145[8:0];
  _RAND_146 = {1{`RANDOM}};
  array4kb_9_ppn2 = _RAND_146[1:0];
  _RAND_147 = {1{`RANDOM}};
  array4kb_9_ppn1 = _RAND_147[8:0];
  _RAND_148 = {1{`RANDOM}};
  array4kb_9_ppn0 = _RAND_148[8:0];
  _RAND_149 = {1{`RANDOM}};
  array4kb_9_asid = _RAND_149[15:0];
  _RAND_150 = {1{`RANDOM}};
  array4kb_10_flag_d = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  array4kb_10_flag_a = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  array4kb_10_flag_g = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  array4kb_10_flag_u = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  array4kb_10_flag_x = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  array4kb_10_flag_w = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  array4kb_10_flag_r = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  array4kb_10_flag_v = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  array4kb_10_vpn2 = _RAND_158[8:0];
  _RAND_159 = {1{`RANDOM}};
  array4kb_10_vpn1 = _RAND_159[8:0];
  _RAND_160 = {1{`RANDOM}};
  array4kb_10_vpn0 = _RAND_160[8:0];
  _RAND_161 = {1{`RANDOM}};
  array4kb_10_ppn2 = _RAND_161[1:0];
  _RAND_162 = {1{`RANDOM}};
  array4kb_10_ppn1 = _RAND_162[8:0];
  _RAND_163 = {1{`RANDOM}};
  array4kb_10_ppn0 = _RAND_163[8:0];
  _RAND_164 = {1{`RANDOM}};
  array4kb_10_asid = _RAND_164[15:0];
  _RAND_165 = {1{`RANDOM}};
  array4kb_11_flag_d = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  array4kb_11_flag_a = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  array4kb_11_flag_g = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  array4kb_11_flag_u = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  array4kb_11_flag_x = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  array4kb_11_flag_w = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  array4kb_11_flag_r = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  array4kb_11_flag_v = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  array4kb_11_vpn2 = _RAND_173[8:0];
  _RAND_174 = {1{`RANDOM}};
  array4kb_11_vpn1 = _RAND_174[8:0];
  _RAND_175 = {1{`RANDOM}};
  array4kb_11_vpn0 = _RAND_175[8:0];
  _RAND_176 = {1{`RANDOM}};
  array4kb_11_ppn2 = _RAND_176[1:0];
  _RAND_177 = {1{`RANDOM}};
  array4kb_11_ppn1 = _RAND_177[8:0];
  _RAND_178 = {1{`RANDOM}};
  array4kb_11_ppn0 = _RAND_178[8:0];
  _RAND_179 = {1{`RANDOM}};
  array4kb_11_asid = _RAND_179[15:0];
  _RAND_180 = {1{`RANDOM}};
  array4kb_12_flag_d = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  array4kb_12_flag_a = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  array4kb_12_flag_g = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  array4kb_12_flag_u = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  array4kb_12_flag_x = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  array4kb_12_flag_w = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  array4kb_12_flag_r = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  array4kb_12_flag_v = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  array4kb_12_vpn2 = _RAND_188[8:0];
  _RAND_189 = {1{`RANDOM}};
  array4kb_12_vpn1 = _RAND_189[8:0];
  _RAND_190 = {1{`RANDOM}};
  array4kb_12_vpn0 = _RAND_190[8:0];
  _RAND_191 = {1{`RANDOM}};
  array4kb_12_ppn2 = _RAND_191[1:0];
  _RAND_192 = {1{`RANDOM}};
  array4kb_12_ppn1 = _RAND_192[8:0];
  _RAND_193 = {1{`RANDOM}};
  array4kb_12_ppn0 = _RAND_193[8:0];
  _RAND_194 = {1{`RANDOM}};
  array4kb_12_asid = _RAND_194[15:0];
  _RAND_195 = {1{`RANDOM}};
  array4kb_13_flag_d = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  array4kb_13_flag_a = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  array4kb_13_flag_g = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  array4kb_13_flag_u = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  array4kb_13_flag_x = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  array4kb_13_flag_w = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  array4kb_13_flag_r = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  array4kb_13_flag_v = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  array4kb_13_vpn2 = _RAND_203[8:0];
  _RAND_204 = {1{`RANDOM}};
  array4kb_13_vpn1 = _RAND_204[8:0];
  _RAND_205 = {1{`RANDOM}};
  array4kb_13_vpn0 = _RAND_205[8:0];
  _RAND_206 = {1{`RANDOM}};
  array4kb_13_ppn2 = _RAND_206[1:0];
  _RAND_207 = {1{`RANDOM}};
  array4kb_13_ppn1 = _RAND_207[8:0];
  _RAND_208 = {1{`RANDOM}};
  array4kb_13_ppn0 = _RAND_208[8:0];
  _RAND_209 = {1{`RANDOM}};
  array4kb_13_asid = _RAND_209[15:0];
  _RAND_210 = {1{`RANDOM}};
  array4kb_14_flag_d = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  array4kb_14_flag_a = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  array4kb_14_flag_g = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  array4kb_14_flag_u = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  array4kb_14_flag_x = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  array4kb_14_flag_w = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  array4kb_14_flag_r = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  array4kb_14_flag_v = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  array4kb_14_vpn2 = _RAND_218[8:0];
  _RAND_219 = {1{`RANDOM}};
  array4kb_14_vpn1 = _RAND_219[8:0];
  _RAND_220 = {1{`RANDOM}};
  array4kb_14_vpn0 = _RAND_220[8:0];
  _RAND_221 = {1{`RANDOM}};
  array4kb_14_ppn2 = _RAND_221[1:0];
  _RAND_222 = {1{`RANDOM}};
  array4kb_14_ppn1 = _RAND_222[8:0];
  _RAND_223 = {1{`RANDOM}};
  array4kb_14_ppn0 = _RAND_223[8:0];
  _RAND_224 = {1{`RANDOM}};
  array4kb_14_asid = _RAND_224[15:0];
  _RAND_225 = {1{`RANDOM}};
  array4kb_15_flag_d = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  array4kb_15_flag_a = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  array4kb_15_flag_g = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  array4kb_15_flag_u = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  array4kb_15_flag_x = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  array4kb_15_flag_w = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  array4kb_15_flag_r = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  array4kb_15_flag_v = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  array4kb_15_vpn2 = _RAND_233[8:0];
  _RAND_234 = {1{`RANDOM}};
  array4kb_15_vpn1 = _RAND_234[8:0];
  _RAND_235 = {1{`RANDOM}};
  array4kb_15_vpn0 = _RAND_235[8:0];
  _RAND_236 = {1{`RANDOM}};
  array4kb_15_ppn2 = _RAND_236[1:0];
  _RAND_237 = {1{`RANDOM}};
  array4kb_15_ppn1 = _RAND_237[8:0];
  _RAND_238 = {1{`RANDOM}};
  array4kb_15_ppn0 = _RAND_238[8:0];
  _RAND_239 = {1{`RANDOM}};
  array4kb_15_asid = _RAND_239[15:0];
  _RAND_240 = {1{`RANDOM}};
  array4kb_16_flag_d = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  array4kb_16_flag_a = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  array4kb_16_flag_g = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  array4kb_16_flag_u = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  array4kb_16_flag_x = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  array4kb_16_flag_w = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  array4kb_16_flag_r = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  array4kb_16_flag_v = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  array4kb_16_vpn2 = _RAND_248[8:0];
  _RAND_249 = {1{`RANDOM}};
  array4kb_16_vpn1 = _RAND_249[8:0];
  _RAND_250 = {1{`RANDOM}};
  array4kb_16_vpn0 = _RAND_250[8:0];
  _RAND_251 = {1{`RANDOM}};
  array4kb_16_ppn2 = _RAND_251[1:0];
  _RAND_252 = {1{`RANDOM}};
  array4kb_16_ppn1 = _RAND_252[8:0];
  _RAND_253 = {1{`RANDOM}};
  array4kb_16_ppn0 = _RAND_253[8:0];
  _RAND_254 = {1{`RANDOM}};
  array4kb_16_asid = _RAND_254[15:0];
  _RAND_255 = {1{`RANDOM}};
  array4kb_17_flag_d = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  array4kb_17_flag_a = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  array4kb_17_flag_g = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  array4kb_17_flag_u = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  array4kb_17_flag_x = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  array4kb_17_flag_w = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  array4kb_17_flag_r = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  array4kb_17_flag_v = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  array4kb_17_vpn2 = _RAND_263[8:0];
  _RAND_264 = {1{`RANDOM}};
  array4kb_17_vpn1 = _RAND_264[8:0];
  _RAND_265 = {1{`RANDOM}};
  array4kb_17_vpn0 = _RAND_265[8:0];
  _RAND_266 = {1{`RANDOM}};
  array4kb_17_ppn2 = _RAND_266[1:0];
  _RAND_267 = {1{`RANDOM}};
  array4kb_17_ppn1 = _RAND_267[8:0];
  _RAND_268 = {1{`RANDOM}};
  array4kb_17_ppn0 = _RAND_268[8:0];
  _RAND_269 = {1{`RANDOM}};
  array4kb_17_asid = _RAND_269[15:0];
  _RAND_270 = {1{`RANDOM}};
  array4kb_18_flag_d = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  array4kb_18_flag_a = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  array4kb_18_flag_g = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  array4kb_18_flag_u = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  array4kb_18_flag_x = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  array4kb_18_flag_w = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  array4kb_18_flag_r = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  array4kb_18_flag_v = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  array4kb_18_vpn2 = _RAND_278[8:0];
  _RAND_279 = {1{`RANDOM}};
  array4kb_18_vpn1 = _RAND_279[8:0];
  _RAND_280 = {1{`RANDOM}};
  array4kb_18_vpn0 = _RAND_280[8:0];
  _RAND_281 = {1{`RANDOM}};
  array4kb_18_ppn2 = _RAND_281[1:0];
  _RAND_282 = {1{`RANDOM}};
  array4kb_18_ppn1 = _RAND_282[8:0];
  _RAND_283 = {1{`RANDOM}};
  array4kb_18_ppn0 = _RAND_283[8:0];
  _RAND_284 = {1{`RANDOM}};
  array4kb_18_asid = _RAND_284[15:0];
  _RAND_285 = {1{`RANDOM}};
  array4kb_19_flag_d = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  array4kb_19_flag_a = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  array4kb_19_flag_g = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  array4kb_19_flag_u = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  array4kb_19_flag_x = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  array4kb_19_flag_w = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  array4kb_19_flag_r = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  array4kb_19_flag_v = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  array4kb_19_vpn2 = _RAND_293[8:0];
  _RAND_294 = {1{`RANDOM}};
  array4kb_19_vpn1 = _RAND_294[8:0];
  _RAND_295 = {1{`RANDOM}};
  array4kb_19_vpn0 = _RAND_295[8:0];
  _RAND_296 = {1{`RANDOM}};
  array4kb_19_ppn2 = _RAND_296[1:0];
  _RAND_297 = {1{`RANDOM}};
  array4kb_19_ppn1 = _RAND_297[8:0];
  _RAND_298 = {1{`RANDOM}};
  array4kb_19_ppn0 = _RAND_298[8:0];
  _RAND_299 = {1{`RANDOM}};
  array4kb_19_asid = _RAND_299[15:0];
  _RAND_300 = {1{`RANDOM}};
  array4kb_20_flag_d = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  array4kb_20_flag_a = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  array4kb_20_flag_g = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  array4kb_20_flag_u = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  array4kb_20_flag_x = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  array4kb_20_flag_w = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  array4kb_20_flag_r = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  array4kb_20_flag_v = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  array4kb_20_vpn2 = _RAND_308[8:0];
  _RAND_309 = {1{`RANDOM}};
  array4kb_20_vpn1 = _RAND_309[8:0];
  _RAND_310 = {1{`RANDOM}};
  array4kb_20_vpn0 = _RAND_310[8:0];
  _RAND_311 = {1{`RANDOM}};
  array4kb_20_ppn2 = _RAND_311[1:0];
  _RAND_312 = {1{`RANDOM}};
  array4kb_20_ppn1 = _RAND_312[8:0];
  _RAND_313 = {1{`RANDOM}};
  array4kb_20_ppn0 = _RAND_313[8:0];
  _RAND_314 = {1{`RANDOM}};
  array4kb_20_asid = _RAND_314[15:0];
  _RAND_315 = {1{`RANDOM}};
  array4kb_21_flag_d = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  array4kb_21_flag_a = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  array4kb_21_flag_g = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  array4kb_21_flag_u = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  array4kb_21_flag_x = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  array4kb_21_flag_w = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  array4kb_21_flag_r = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  array4kb_21_flag_v = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  array4kb_21_vpn2 = _RAND_323[8:0];
  _RAND_324 = {1{`RANDOM}};
  array4kb_21_vpn1 = _RAND_324[8:0];
  _RAND_325 = {1{`RANDOM}};
  array4kb_21_vpn0 = _RAND_325[8:0];
  _RAND_326 = {1{`RANDOM}};
  array4kb_21_ppn2 = _RAND_326[1:0];
  _RAND_327 = {1{`RANDOM}};
  array4kb_21_ppn1 = _RAND_327[8:0];
  _RAND_328 = {1{`RANDOM}};
  array4kb_21_ppn0 = _RAND_328[8:0];
  _RAND_329 = {1{`RANDOM}};
  array4kb_21_asid = _RAND_329[15:0];
  _RAND_330 = {1{`RANDOM}};
  array4kb_22_flag_d = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  array4kb_22_flag_a = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  array4kb_22_flag_g = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  array4kb_22_flag_u = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  array4kb_22_flag_x = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  array4kb_22_flag_w = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  array4kb_22_flag_r = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  array4kb_22_flag_v = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  array4kb_22_vpn2 = _RAND_338[8:0];
  _RAND_339 = {1{`RANDOM}};
  array4kb_22_vpn1 = _RAND_339[8:0];
  _RAND_340 = {1{`RANDOM}};
  array4kb_22_vpn0 = _RAND_340[8:0];
  _RAND_341 = {1{`RANDOM}};
  array4kb_22_ppn2 = _RAND_341[1:0];
  _RAND_342 = {1{`RANDOM}};
  array4kb_22_ppn1 = _RAND_342[8:0];
  _RAND_343 = {1{`RANDOM}};
  array4kb_22_ppn0 = _RAND_343[8:0];
  _RAND_344 = {1{`RANDOM}};
  array4kb_22_asid = _RAND_344[15:0];
  _RAND_345 = {1{`RANDOM}};
  array4kb_23_flag_d = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  array4kb_23_flag_a = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  array4kb_23_flag_g = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  array4kb_23_flag_u = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  array4kb_23_flag_x = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  array4kb_23_flag_w = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  array4kb_23_flag_r = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  array4kb_23_flag_v = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  array4kb_23_vpn2 = _RAND_353[8:0];
  _RAND_354 = {1{`RANDOM}};
  array4kb_23_vpn1 = _RAND_354[8:0];
  _RAND_355 = {1{`RANDOM}};
  array4kb_23_vpn0 = _RAND_355[8:0];
  _RAND_356 = {1{`RANDOM}};
  array4kb_23_ppn2 = _RAND_356[1:0];
  _RAND_357 = {1{`RANDOM}};
  array4kb_23_ppn1 = _RAND_357[8:0];
  _RAND_358 = {1{`RANDOM}};
  array4kb_23_ppn0 = _RAND_358[8:0];
  _RAND_359 = {1{`RANDOM}};
  array4kb_23_asid = _RAND_359[15:0];
  _RAND_360 = {1{`RANDOM}};
  array4kb_24_flag_d = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  array4kb_24_flag_a = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  array4kb_24_flag_g = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  array4kb_24_flag_u = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  array4kb_24_flag_x = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  array4kb_24_flag_w = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  array4kb_24_flag_r = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  array4kb_24_flag_v = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  array4kb_24_vpn2 = _RAND_368[8:0];
  _RAND_369 = {1{`RANDOM}};
  array4kb_24_vpn1 = _RAND_369[8:0];
  _RAND_370 = {1{`RANDOM}};
  array4kb_24_vpn0 = _RAND_370[8:0];
  _RAND_371 = {1{`RANDOM}};
  array4kb_24_ppn2 = _RAND_371[1:0];
  _RAND_372 = {1{`RANDOM}};
  array4kb_24_ppn1 = _RAND_372[8:0];
  _RAND_373 = {1{`RANDOM}};
  array4kb_24_ppn0 = _RAND_373[8:0];
  _RAND_374 = {1{`RANDOM}};
  array4kb_24_asid = _RAND_374[15:0];
  _RAND_375 = {1{`RANDOM}};
  array4kb_25_flag_d = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  array4kb_25_flag_a = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  array4kb_25_flag_g = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  array4kb_25_flag_u = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  array4kb_25_flag_x = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  array4kb_25_flag_w = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  array4kb_25_flag_r = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  array4kb_25_flag_v = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  array4kb_25_vpn2 = _RAND_383[8:0];
  _RAND_384 = {1{`RANDOM}};
  array4kb_25_vpn1 = _RAND_384[8:0];
  _RAND_385 = {1{`RANDOM}};
  array4kb_25_vpn0 = _RAND_385[8:0];
  _RAND_386 = {1{`RANDOM}};
  array4kb_25_ppn2 = _RAND_386[1:0];
  _RAND_387 = {1{`RANDOM}};
  array4kb_25_ppn1 = _RAND_387[8:0];
  _RAND_388 = {1{`RANDOM}};
  array4kb_25_ppn0 = _RAND_388[8:0];
  _RAND_389 = {1{`RANDOM}};
  array4kb_25_asid = _RAND_389[15:0];
  _RAND_390 = {1{`RANDOM}};
  array4kb_26_flag_d = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  array4kb_26_flag_a = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  array4kb_26_flag_g = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  array4kb_26_flag_u = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  array4kb_26_flag_x = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  array4kb_26_flag_w = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  array4kb_26_flag_r = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  array4kb_26_flag_v = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  array4kb_26_vpn2 = _RAND_398[8:0];
  _RAND_399 = {1{`RANDOM}};
  array4kb_26_vpn1 = _RAND_399[8:0];
  _RAND_400 = {1{`RANDOM}};
  array4kb_26_vpn0 = _RAND_400[8:0];
  _RAND_401 = {1{`RANDOM}};
  array4kb_26_ppn2 = _RAND_401[1:0];
  _RAND_402 = {1{`RANDOM}};
  array4kb_26_ppn1 = _RAND_402[8:0];
  _RAND_403 = {1{`RANDOM}};
  array4kb_26_ppn0 = _RAND_403[8:0];
  _RAND_404 = {1{`RANDOM}};
  array4kb_26_asid = _RAND_404[15:0];
  _RAND_405 = {1{`RANDOM}};
  array4kb_27_flag_d = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  array4kb_27_flag_a = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  array4kb_27_flag_g = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  array4kb_27_flag_u = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  array4kb_27_flag_x = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  array4kb_27_flag_w = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  array4kb_27_flag_r = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  array4kb_27_flag_v = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  array4kb_27_vpn2 = _RAND_413[8:0];
  _RAND_414 = {1{`RANDOM}};
  array4kb_27_vpn1 = _RAND_414[8:0];
  _RAND_415 = {1{`RANDOM}};
  array4kb_27_vpn0 = _RAND_415[8:0];
  _RAND_416 = {1{`RANDOM}};
  array4kb_27_ppn2 = _RAND_416[1:0];
  _RAND_417 = {1{`RANDOM}};
  array4kb_27_ppn1 = _RAND_417[8:0];
  _RAND_418 = {1{`RANDOM}};
  array4kb_27_ppn0 = _RAND_418[8:0];
  _RAND_419 = {1{`RANDOM}};
  array4kb_27_asid = _RAND_419[15:0];
  _RAND_420 = {1{`RANDOM}};
  array4kb_28_flag_d = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  array4kb_28_flag_a = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  array4kb_28_flag_g = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  array4kb_28_flag_u = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  array4kb_28_flag_x = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  array4kb_28_flag_w = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  array4kb_28_flag_r = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  array4kb_28_flag_v = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  array4kb_28_vpn2 = _RAND_428[8:0];
  _RAND_429 = {1{`RANDOM}};
  array4kb_28_vpn1 = _RAND_429[8:0];
  _RAND_430 = {1{`RANDOM}};
  array4kb_28_vpn0 = _RAND_430[8:0];
  _RAND_431 = {1{`RANDOM}};
  array4kb_28_ppn2 = _RAND_431[1:0];
  _RAND_432 = {1{`RANDOM}};
  array4kb_28_ppn1 = _RAND_432[8:0];
  _RAND_433 = {1{`RANDOM}};
  array4kb_28_ppn0 = _RAND_433[8:0];
  _RAND_434 = {1{`RANDOM}};
  array4kb_28_asid = _RAND_434[15:0];
  _RAND_435 = {1{`RANDOM}};
  array4kb_29_flag_d = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  array4kb_29_flag_a = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  array4kb_29_flag_g = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  array4kb_29_flag_u = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  array4kb_29_flag_x = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  array4kb_29_flag_w = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  array4kb_29_flag_r = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  array4kb_29_flag_v = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  array4kb_29_vpn2 = _RAND_443[8:0];
  _RAND_444 = {1{`RANDOM}};
  array4kb_29_vpn1 = _RAND_444[8:0];
  _RAND_445 = {1{`RANDOM}};
  array4kb_29_vpn0 = _RAND_445[8:0];
  _RAND_446 = {1{`RANDOM}};
  array4kb_29_ppn2 = _RAND_446[1:0];
  _RAND_447 = {1{`RANDOM}};
  array4kb_29_ppn1 = _RAND_447[8:0];
  _RAND_448 = {1{`RANDOM}};
  array4kb_29_ppn0 = _RAND_448[8:0];
  _RAND_449 = {1{`RANDOM}};
  array4kb_29_asid = _RAND_449[15:0];
  _RAND_450 = {1{`RANDOM}};
  array4kb_30_flag_d = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  array4kb_30_flag_a = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  array4kb_30_flag_g = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  array4kb_30_flag_u = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  array4kb_30_flag_x = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  array4kb_30_flag_w = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  array4kb_30_flag_r = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  array4kb_30_flag_v = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  array4kb_30_vpn2 = _RAND_458[8:0];
  _RAND_459 = {1{`RANDOM}};
  array4kb_30_vpn1 = _RAND_459[8:0];
  _RAND_460 = {1{`RANDOM}};
  array4kb_30_vpn0 = _RAND_460[8:0];
  _RAND_461 = {1{`RANDOM}};
  array4kb_30_ppn2 = _RAND_461[1:0];
  _RAND_462 = {1{`RANDOM}};
  array4kb_30_ppn1 = _RAND_462[8:0];
  _RAND_463 = {1{`RANDOM}};
  array4kb_30_ppn0 = _RAND_463[8:0];
  _RAND_464 = {1{`RANDOM}};
  array4kb_30_asid = _RAND_464[15:0];
  _RAND_465 = {1{`RANDOM}};
  array4kb_31_flag_d = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  array4kb_31_flag_a = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  array4kb_31_flag_g = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  array4kb_31_flag_u = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  array4kb_31_flag_x = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  array4kb_31_flag_w = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  array4kb_31_flag_r = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  array4kb_31_flag_v = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  array4kb_31_vpn2 = _RAND_473[8:0];
  _RAND_474 = {1{`RANDOM}};
  array4kb_31_vpn1 = _RAND_474[8:0];
  _RAND_475 = {1{`RANDOM}};
  array4kb_31_vpn0 = _RAND_475[8:0];
  _RAND_476 = {1{`RANDOM}};
  array4kb_31_ppn2 = _RAND_476[1:0];
  _RAND_477 = {1{`RANDOM}};
  array4kb_31_ppn1 = _RAND_477[8:0];
  _RAND_478 = {1{`RANDOM}};
  array4kb_31_ppn0 = _RAND_478[8:0];
  _RAND_479 = {1{`RANDOM}};
  array4kb_31_asid = _RAND_479[15:0];
  _RAND_480 = {1{`RANDOM}};
  array4kb_valid_0 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  array4kb_valid_1 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  array4kb_valid_2 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  array4kb_valid_3 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  array4kb_valid_4 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  array4kb_valid_5 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  array4kb_valid_6 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  array4kb_valid_7 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  array4kb_valid_8 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  array4kb_valid_9 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  array4kb_valid_10 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  array4kb_valid_11 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  array4kb_valid_12 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  array4kb_valid_13 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  array4kb_valid_14 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  array4kb_valid_15 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  array4kb_valid_16 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  array4kb_valid_17 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  array4kb_valid_18 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  array4kb_valid_19 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  array4kb_valid_20 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  array4kb_valid_21 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  array4kb_valid_22 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  array4kb_valid_23 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  array4kb_valid_24 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  array4kb_valid_25 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  array4kb_valid_26 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  array4kb_valid_27 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  array4kb_valid_28 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  array4kb_valid_29 = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  array4kb_valid_30 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  array4kb_valid_31 = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  array2mb_0_flag_d = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  array2mb_0_flag_a = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  array2mb_0_flag_g = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  array2mb_0_flag_u = _RAND_515[0:0];
  _RAND_516 = {1{`RANDOM}};
  array2mb_0_flag_x = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  array2mb_0_flag_w = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  array2mb_0_flag_r = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  array2mb_0_flag_v = _RAND_519[0:0];
  _RAND_520 = {1{`RANDOM}};
  array2mb_0_vpn2 = _RAND_520[8:0];
  _RAND_521 = {1{`RANDOM}};
  array2mb_0_vpn1 = _RAND_521[8:0];
  _RAND_522 = {1{`RANDOM}};
  array2mb_0_ppn2 = _RAND_522[1:0];
  _RAND_523 = {1{`RANDOM}};
  array2mb_0_ppn1 = _RAND_523[8:0];
  _RAND_524 = {1{`RANDOM}};
  array2mb_0_asid = _RAND_524[15:0];
  _RAND_525 = {1{`RANDOM}};
  array2mb_1_flag_d = _RAND_525[0:0];
  _RAND_526 = {1{`RANDOM}};
  array2mb_1_flag_a = _RAND_526[0:0];
  _RAND_527 = {1{`RANDOM}};
  array2mb_1_flag_g = _RAND_527[0:0];
  _RAND_528 = {1{`RANDOM}};
  array2mb_1_flag_u = _RAND_528[0:0];
  _RAND_529 = {1{`RANDOM}};
  array2mb_1_flag_x = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  array2mb_1_flag_w = _RAND_530[0:0];
  _RAND_531 = {1{`RANDOM}};
  array2mb_1_flag_r = _RAND_531[0:0];
  _RAND_532 = {1{`RANDOM}};
  array2mb_1_flag_v = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  array2mb_1_vpn2 = _RAND_533[8:0];
  _RAND_534 = {1{`RANDOM}};
  array2mb_1_vpn1 = _RAND_534[8:0];
  _RAND_535 = {1{`RANDOM}};
  array2mb_1_ppn2 = _RAND_535[1:0];
  _RAND_536 = {1{`RANDOM}};
  array2mb_1_ppn1 = _RAND_536[8:0];
  _RAND_537 = {1{`RANDOM}};
  array2mb_1_asid = _RAND_537[15:0];
  _RAND_538 = {1{`RANDOM}};
  array2mb_2_flag_d = _RAND_538[0:0];
  _RAND_539 = {1{`RANDOM}};
  array2mb_2_flag_a = _RAND_539[0:0];
  _RAND_540 = {1{`RANDOM}};
  array2mb_2_flag_g = _RAND_540[0:0];
  _RAND_541 = {1{`RANDOM}};
  array2mb_2_flag_u = _RAND_541[0:0];
  _RAND_542 = {1{`RANDOM}};
  array2mb_2_flag_x = _RAND_542[0:0];
  _RAND_543 = {1{`RANDOM}};
  array2mb_2_flag_w = _RAND_543[0:0];
  _RAND_544 = {1{`RANDOM}};
  array2mb_2_flag_r = _RAND_544[0:0];
  _RAND_545 = {1{`RANDOM}};
  array2mb_2_flag_v = _RAND_545[0:0];
  _RAND_546 = {1{`RANDOM}};
  array2mb_2_vpn2 = _RAND_546[8:0];
  _RAND_547 = {1{`RANDOM}};
  array2mb_2_vpn1 = _RAND_547[8:0];
  _RAND_548 = {1{`RANDOM}};
  array2mb_2_ppn2 = _RAND_548[1:0];
  _RAND_549 = {1{`RANDOM}};
  array2mb_2_ppn1 = _RAND_549[8:0];
  _RAND_550 = {1{`RANDOM}};
  array2mb_2_asid = _RAND_550[15:0];
  _RAND_551 = {1{`RANDOM}};
  array2mb_3_flag_d = _RAND_551[0:0];
  _RAND_552 = {1{`RANDOM}};
  array2mb_3_flag_a = _RAND_552[0:0];
  _RAND_553 = {1{`RANDOM}};
  array2mb_3_flag_g = _RAND_553[0:0];
  _RAND_554 = {1{`RANDOM}};
  array2mb_3_flag_u = _RAND_554[0:0];
  _RAND_555 = {1{`RANDOM}};
  array2mb_3_flag_x = _RAND_555[0:0];
  _RAND_556 = {1{`RANDOM}};
  array2mb_3_flag_w = _RAND_556[0:0];
  _RAND_557 = {1{`RANDOM}};
  array2mb_3_flag_r = _RAND_557[0:0];
  _RAND_558 = {1{`RANDOM}};
  array2mb_3_flag_v = _RAND_558[0:0];
  _RAND_559 = {1{`RANDOM}};
  array2mb_3_vpn2 = _RAND_559[8:0];
  _RAND_560 = {1{`RANDOM}};
  array2mb_3_vpn1 = _RAND_560[8:0];
  _RAND_561 = {1{`RANDOM}};
  array2mb_3_ppn2 = _RAND_561[1:0];
  _RAND_562 = {1{`RANDOM}};
  array2mb_3_ppn1 = _RAND_562[8:0];
  _RAND_563 = {1{`RANDOM}};
  array2mb_3_asid = _RAND_563[15:0];
  _RAND_564 = {1{`RANDOM}};
  array2mb_4_flag_d = _RAND_564[0:0];
  _RAND_565 = {1{`RANDOM}};
  array2mb_4_flag_a = _RAND_565[0:0];
  _RAND_566 = {1{`RANDOM}};
  array2mb_4_flag_g = _RAND_566[0:0];
  _RAND_567 = {1{`RANDOM}};
  array2mb_4_flag_u = _RAND_567[0:0];
  _RAND_568 = {1{`RANDOM}};
  array2mb_4_flag_x = _RAND_568[0:0];
  _RAND_569 = {1{`RANDOM}};
  array2mb_4_flag_w = _RAND_569[0:0];
  _RAND_570 = {1{`RANDOM}};
  array2mb_4_flag_r = _RAND_570[0:0];
  _RAND_571 = {1{`RANDOM}};
  array2mb_4_flag_v = _RAND_571[0:0];
  _RAND_572 = {1{`RANDOM}};
  array2mb_4_vpn2 = _RAND_572[8:0];
  _RAND_573 = {1{`RANDOM}};
  array2mb_4_vpn1 = _RAND_573[8:0];
  _RAND_574 = {1{`RANDOM}};
  array2mb_4_ppn2 = _RAND_574[1:0];
  _RAND_575 = {1{`RANDOM}};
  array2mb_4_ppn1 = _RAND_575[8:0];
  _RAND_576 = {1{`RANDOM}};
  array2mb_4_asid = _RAND_576[15:0];
  _RAND_577 = {1{`RANDOM}};
  array2mb_5_flag_d = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  array2mb_5_flag_a = _RAND_578[0:0];
  _RAND_579 = {1{`RANDOM}};
  array2mb_5_flag_g = _RAND_579[0:0];
  _RAND_580 = {1{`RANDOM}};
  array2mb_5_flag_u = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  array2mb_5_flag_x = _RAND_581[0:0];
  _RAND_582 = {1{`RANDOM}};
  array2mb_5_flag_w = _RAND_582[0:0];
  _RAND_583 = {1{`RANDOM}};
  array2mb_5_flag_r = _RAND_583[0:0];
  _RAND_584 = {1{`RANDOM}};
  array2mb_5_flag_v = _RAND_584[0:0];
  _RAND_585 = {1{`RANDOM}};
  array2mb_5_vpn2 = _RAND_585[8:0];
  _RAND_586 = {1{`RANDOM}};
  array2mb_5_vpn1 = _RAND_586[8:0];
  _RAND_587 = {1{`RANDOM}};
  array2mb_5_ppn2 = _RAND_587[1:0];
  _RAND_588 = {1{`RANDOM}};
  array2mb_5_ppn1 = _RAND_588[8:0];
  _RAND_589 = {1{`RANDOM}};
  array2mb_5_asid = _RAND_589[15:0];
  _RAND_590 = {1{`RANDOM}};
  array2mb_6_flag_d = _RAND_590[0:0];
  _RAND_591 = {1{`RANDOM}};
  array2mb_6_flag_a = _RAND_591[0:0];
  _RAND_592 = {1{`RANDOM}};
  array2mb_6_flag_g = _RAND_592[0:0];
  _RAND_593 = {1{`RANDOM}};
  array2mb_6_flag_u = _RAND_593[0:0];
  _RAND_594 = {1{`RANDOM}};
  array2mb_6_flag_x = _RAND_594[0:0];
  _RAND_595 = {1{`RANDOM}};
  array2mb_6_flag_w = _RAND_595[0:0];
  _RAND_596 = {1{`RANDOM}};
  array2mb_6_flag_r = _RAND_596[0:0];
  _RAND_597 = {1{`RANDOM}};
  array2mb_6_flag_v = _RAND_597[0:0];
  _RAND_598 = {1{`RANDOM}};
  array2mb_6_vpn2 = _RAND_598[8:0];
  _RAND_599 = {1{`RANDOM}};
  array2mb_6_vpn1 = _RAND_599[8:0];
  _RAND_600 = {1{`RANDOM}};
  array2mb_6_ppn2 = _RAND_600[1:0];
  _RAND_601 = {1{`RANDOM}};
  array2mb_6_ppn1 = _RAND_601[8:0];
  _RAND_602 = {1{`RANDOM}};
  array2mb_6_asid = _RAND_602[15:0];
  _RAND_603 = {1{`RANDOM}};
  array2mb_7_flag_d = _RAND_603[0:0];
  _RAND_604 = {1{`RANDOM}};
  array2mb_7_flag_a = _RAND_604[0:0];
  _RAND_605 = {1{`RANDOM}};
  array2mb_7_flag_g = _RAND_605[0:0];
  _RAND_606 = {1{`RANDOM}};
  array2mb_7_flag_u = _RAND_606[0:0];
  _RAND_607 = {1{`RANDOM}};
  array2mb_7_flag_x = _RAND_607[0:0];
  _RAND_608 = {1{`RANDOM}};
  array2mb_7_flag_w = _RAND_608[0:0];
  _RAND_609 = {1{`RANDOM}};
  array2mb_7_flag_r = _RAND_609[0:0];
  _RAND_610 = {1{`RANDOM}};
  array2mb_7_flag_v = _RAND_610[0:0];
  _RAND_611 = {1{`RANDOM}};
  array2mb_7_vpn2 = _RAND_611[8:0];
  _RAND_612 = {1{`RANDOM}};
  array2mb_7_vpn1 = _RAND_612[8:0];
  _RAND_613 = {1{`RANDOM}};
  array2mb_7_ppn2 = _RAND_613[1:0];
  _RAND_614 = {1{`RANDOM}};
  array2mb_7_ppn1 = _RAND_614[8:0];
  _RAND_615 = {1{`RANDOM}};
  array2mb_7_asid = _RAND_615[15:0];
  _RAND_616 = {1{`RANDOM}};
  array2mb_valid_0 = _RAND_616[0:0];
  _RAND_617 = {1{`RANDOM}};
  array2mb_valid_1 = _RAND_617[0:0];
  _RAND_618 = {1{`RANDOM}};
  array2mb_valid_2 = _RAND_618[0:0];
  _RAND_619 = {1{`RANDOM}};
  array2mb_valid_3 = _RAND_619[0:0];
  _RAND_620 = {1{`RANDOM}};
  array2mb_valid_4 = _RAND_620[0:0];
  _RAND_621 = {1{`RANDOM}};
  array2mb_valid_5 = _RAND_621[0:0];
  _RAND_622 = {1{`RANDOM}};
  array2mb_valid_6 = _RAND_622[0:0];
  _RAND_623 = {1{`RANDOM}};
  array2mb_valid_7 = _RAND_623[0:0];
  _RAND_624 = {1{`RANDOM}};
  array1gb_0_flag_d = _RAND_624[0:0];
  _RAND_625 = {1{`RANDOM}};
  array1gb_0_flag_a = _RAND_625[0:0];
  _RAND_626 = {1{`RANDOM}};
  array1gb_0_flag_g = _RAND_626[0:0];
  _RAND_627 = {1{`RANDOM}};
  array1gb_0_flag_u = _RAND_627[0:0];
  _RAND_628 = {1{`RANDOM}};
  array1gb_0_flag_x = _RAND_628[0:0];
  _RAND_629 = {1{`RANDOM}};
  array1gb_0_flag_w = _RAND_629[0:0];
  _RAND_630 = {1{`RANDOM}};
  array1gb_0_flag_r = _RAND_630[0:0];
  _RAND_631 = {1{`RANDOM}};
  array1gb_0_flag_v = _RAND_631[0:0];
  _RAND_632 = {1{`RANDOM}};
  array1gb_0_vpn2 = _RAND_632[8:0];
  _RAND_633 = {1{`RANDOM}};
  array1gb_0_ppn2 = _RAND_633[1:0];
  _RAND_634 = {1{`RANDOM}};
  array1gb_0_asid = _RAND_634[15:0];
  _RAND_635 = {1{`RANDOM}};
  array1gb_1_flag_d = _RAND_635[0:0];
  _RAND_636 = {1{`RANDOM}};
  array1gb_1_flag_a = _RAND_636[0:0];
  _RAND_637 = {1{`RANDOM}};
  array1gb_1_flag_g = _RAND_637[0:0];
  _RAND_638 = {1{`RANDOM}};
  array1gb_1_flag_u = _RAND_638[0:0];
  _RAND_639 = {1{`RANDOM}};
  array1gb_1_flag_x = _RAND_639[0:0];
  _RAND_640 = {1{`RANDOM}};
  array1gb_1_flag_w = _RAND_640[0:0];
  _RAND_641 = {1{`RANDOM}};
  array1gb_1_flag_r = _RAND_641[0:0];
  _RAND_642 = {1{`RANDOM}};
  array1gb_1_flag_v = _RAND_642[0:0];
  _RAND_643 = {1{`RANDOM}};
  array1gb_1_vpn2 = _RAND_643[8:0];
  _RAND_644 = {1{`RANDOM}};
  array1gb_1_ppn2 = _RAND_644[1:0];
  _RAND_645 = {1{`RANDOM}};
  array1gb_1_asid = _RAND_645[15:0];
  _RAND_646 = {1{`RANDOM}};
  array1gb_2_flag_d = _RAND_646[0:0];
  _RAND_647 = {1{`RANDOM}};
  array1gb_2_flag_a = _RAND_647[0:0];
  _RAND_648 = {1{`RANDOM}};
  array1gb_2_flag_g = _RAND_648[0:0];
  _RAND_649 = {1{`RANDOM}};
  array1gb_2_flag_u = _RAND_649[0:0];
  _RAND_650 = {1{`RANDOM}};
  array1gb_2_flag_x = _RAND_650[0:0];
  _RAND_651 = {1{`RANDOM}};
  array1gb_2_flag_w = _RAND_651[0:0];
  _RAND_652 = {1{`RANDOM}};
  array1gb_2_flag_r = _RAND_652[0:0];
  _RAND_653 = {1{`RANDOM}};
  array1gb_2_flag_v = _RAND_653[0:0];
  _RAND_654 = {1{`RANDOM}};
  array1gb_2_vpn2 = _RAND_654[8:0];
  _RAND_655 = {1{`RANDOM}};
  array1gb_2_ppn2 = _RAND_655[1:0];
  _RAND_656 = {1{`RANDOM}};
  array1gb_2_asid = _RAND_656[15:0];
  _RAND_657 = {1{`RANDOM}};
  array1gb_3_flag_d = _RAND_657[0:0];
  _RAND_658 = {1{`RANDOM}};
  array1gb_3_flag_a = _RAND_658[0:0];
  _RAND_659 = {1{`RANDOM}};
  array1gb_3_flag_g = _RAND_659[0:0];
  _RAND_660 = {1{`RANDOM}};
  array1gb_3_flag_u = _RAND_660[0:0];
  _RAND_661 = {1{`RANDOM}};
  array1gb_3_flag_x = _RAND_661[0:0];
  _RAND_662 = {1{`RANDOM}};
  array1gb_3_flag_w = _RAND_662[0:0];
  _RAND_663 = {1{`RANDOM}};
  array1gb_3_flag_r = _RAND_663[0:0];
  _RAND_664 = {1{`RANDOM}};
  array1gb_3_flag_v = _RAND_664[0:0];
  _RAND_665 = {1{`RANDOM}};
  array1gb_3_vpn2 = _RAND_665[8:0];
  _RAND_666 = {1{`RANDOM}};
  array1gb_3_ppn2 = _RAND_666[1:0];
  _RAND_667 = {1{`RANDOM}};
  array1gb_3_asid = _RAND_667[15:0];
  _RAND_668 = {1{`RANDOM}};
  array1gb_valid_0 = _RAND_668[0:0];
  _RAND_669 = {1{`RANDOM}};
  array1gb_valid_1 = _RAND_669[0:0];
  _RAND_670 = {1{`RANDOM}};
  array1gb_valid_2 = _RAND_670[0:0];
  _RAND_671 = {1{`RANDOM}};
  array1gb_valid_3 = _RAND_671[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CachePortProxy(
  input         clock,
  input         reset,
  input  [1:0]  io_prv,
  input         io_sv39_en,
  input  [15:0] io_satp_asid,
  input  [43:0] io_satp_ppn,
  input         io_sfence_vma,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [38:0] io_in_req_bits_addr,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [63:0] io_in_resp_bits_rdata,
  output        io_in_resp_bits_page_fault,
  output        io_in_resp_bits_access_fault,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [38:0] io_out_req_bits_addr,
  output        io_out_resp_ready,
  input         io_out_resp_valid,
  input  [63:0] io_out_resp_bits_rdata,
  input         io_ptw_req_ready,
  output        io_ptw_req_valid,
  output [38:0] io_ptw_req_bits_addr,
  output        io_ptw_resp_ready,
  input         io_ptw_resp_valid,
  input  [63:0] io_ptw_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  wire  tlb_clock; // @[CachePortProxy.scala 28:19]
  wire  tlb_reset; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_sfence_vma; // @[CachePortProxy.scala 28:19]
  wire [8:0] tlb_io_vaddr_vpn2; // @[CachePortProxy.scala 28:19]
  wire [8:0] tlb_io_vaddr_vpn1; // @[CachePortProxy.scala 28:19]
  wire [8:0] tlb_io_vaddr_vpn0; // @[CachePortProxy.scala 28:19]
  wire [1:0] tlb_io_rpte_ppn2; // @[CachePortProxy.scala 28:19]
  wire [8:0] tlb_io_rpte_ppn1; // @[CachePortProxy.scala 28:19]
  wire [8:0] tlb_io_rpte_ppn0; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_rpte_flag_d; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_rpte_flag_a; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_rpte_flag_u; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_rpte_flag_x; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_rpte_flag_w; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_rpte_flag_r; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_rpte_flag_v; // @[CachePortProxy.scala 28:19]
  wire [1:0] tlb_io_rlevel; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_hit; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_wen; // @[CachePortProxy.scala 28:19]
  wire [8:0] tlb_io_wvaddr_vpn2; // @[CachePortProxy.scala 28:19]
  wire [8:0] tlb_io_wvaddr_vpn1; // @[CachePortProxy.scala 28:19]
  wire [8:0] tlb_io_wvaddr_vpn0; // @[CachePortProxy.scala 28:19]
  wire [1:0] tlb_io_wpte_ppn2; // @[CachePortProxy.scala 28:19]
  wire [8:0] tlb_io_wpte_ppn1; // @[CachePortProxy.scala 28:19]
  wire [8:0] tlb_io_wpte_ppn0; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_wpte_flag_d; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_wpte_flag_a; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_wpte_flag_g; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_wpte_flag_u; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_wpte_flag_x; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_wpte_flag_w; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_wpte_flag_r; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_wpte_flag_v; // @[CachePortProxy.scala 28:19]
  wire [1:0] tlb_io_wlevel; // @[CachePortProxy.scala 28:19]
  wire [15:0] tlb_io_satp_asid; // @[CachePortProxy.scala 28:19]
  reg [2:0] state; // @[CachePortProxy.scala 21:93]
  wire  _in_req_bits_T = state == 3'h0; // @[CachePortProxy.scala 24:54]
  reg [38:0] in_req_bits_r_addr; // @[Reg.scala 35:20]
  wire [38:0] _GEN_0 = _in_req_bits_T ? io_in_req_bits_addr : in_req_bits_r_addr; // @[Reg.scala 36:18 35:20 36:22]
  wire [11:0] in_vaddr_offset = _GEN_0[11:0]; // @[CachePortProxy.scala 25:46]
  wire [8:0] in_vaddr_vpn0 = _GEN_0[20:12]; // @[CachePortProxy.scala 25:46]
  wire [8:0] in_vaddr_vpn1 = _GEN_0[29:21]; // @[CachePortProxy.scala 25:46]
  wire [8:0] in_vaddr_vpn2 = _GEN_0[38:30]; // @[CachePortProxy.scala 25:46]
  wire  _atp_en_T_1 = io_prv != 2'h3 & io_sv39_en; // @[CachePortProxy.scala 38:48]
  reg  atp_en_r; // @[Reg.scala 35:20]
  wire  _GEN_7 = _in_req_bits_T ? _atp_en_T_1 : atp_en_r; // @[Reg.scala 36:18 35:20 36:22]
  wire  in_addr_boot = io_in_req_bits_addr >= 39'h10000 & io_in_req_bits_addr <= 39'h30000; // @[CachePortProxy.scala 42:50]
  wire  in_addr_clint = io_in_req_bits_addr >= 39'h2000000 & io_in_req_bits_addr <= 39'h200ffff; // @[CachePortProxy.scala 43:50]
  wire  in_addr_plic = io_in_req_bits_addr >= 39'hc000000 & io_in_req_bits_addr <= 39'hfffffff; // @[CachePortProxy.scala 44:50]
  wire  in_addr_uart = io_in_req_bits_addr >= 39'h10000000 & io_in_req_bits_addr <= 39'h1000ffff; // @[CachePortProxy.scala 45:50]
  wire  _access_fault_T_3 = ~_GEN_7; // @[CachePortProxy.scala 46:70]
  wire  _access_fault_T_9 = ~(in_addr_boot | in_addr_clint | in_addr_plic | in_addr_uart); // @[CachePortProxy.scala 47:5]
  wire  access_fault = ~io_in_req_bits_addr[31] & (io_prv == 2'h3 | ~_GEN_7) & _access_fault_T_9; // @[CachePortProxy.scala 46:79]
  reg [1:0] ptw_level; // @[CachePortProxy.scala 50:29]
  wire  ptw_pte_flag_v = io_ptw_resp_bits_rdata[0]; // @[CachePortProxy.scala 51:53]
  wire  ptw_pte_flag_r = io_ptw_resp_bits_rdata[1]; // @[CachePortProxy.scala 51:53]
  wire  ptw_pte_flag_w = io_ptw_resp_bits_rdata[2]; // @[CachePortProxy.scala 51:53]
  wire  ptw_pte_flag_x = io_ptw_resp_bits_rdata[3]; // @[CachePortProxy.scala 51:53]
  wire  ptw_pte_flag_u = io_ptw_resp_bits_rdata[4]; // @[CachePortProxy.scala 51:53]
  wire  ptw_pte_flag_g = io_ptw_resp_bits_rdata[5]; // @[CachePortProxy.scala 51:53]
  wire  ptw_pte_flag_a = io_ptw_resp_bits_rdata[6]; // @[CachePortProxy.scala 51:53]
  wire  ptw_pte_flag_d = io_ptw_resp_bits_rdata[7]; // @[CachePortProxy.scala 51:53]
  wire [8:0] ptw_pte_ppn0 = io_ptw_resp_bits_rdata[18:10]; // @[CachePortProxy.scala 51:53]
  wire [8:0] ptw_pte_ppn1 = io_ptw_resp_bits_rdata[27:19]; // @[CachePortProxy.scala 51:53]
  wire [1:0] ptw_pte_ppn2 = io_ptw_resp_bits_rdata[29:28]; // @[CachePortProxy.scala 51:53]
  wire  _ptw_pte_reg_T = io_ptw_resp_ready & io_ptw_resp_valid; // @[Decoupled.scala 51:35]
  reg [1:0] ptw_pte_reg_ppn2; // @[Reg.scala 35:20]
  reg [8:0] ptw_pte_reg_ppn1; // @[Reg.scala 35:20]
  reg [8:0] ptw_pte_reg_ppn0; // @[Reg.scala 35:20]
  reg  ptw_pte_reg_flag_d; // @[Reg.scala 35:20]
  reg  ptw_pte_reg_flag_a; // @[Reg.scala 35:20]
  reg  ptw_pte_reg_flag_g; // @[Reg.scala 35:20]
  reg  ptw_pte_reg_flag_u; // @[Reg.scala 35:20]
  reg  ptw_pte_reg_flag_x; // @[Reg.scala 35:20]
  reg  ptw_pte_reg_flag_w; // @[Reg.scala 35:20]
  reg  ptw_pte_reg_flag_r; // @[Reg.scala 35:20]
  reg  ptw_pte_reg_flag_v; // @[Reg.scala 35:20]
  wire  _ptw_complete_T_4 = ptw_pte_flag_r | ptw_pte_flag_x; // @[CachePortProxy.scala 7:37]
  wire  ptw_complete = ~ptw_pte_flag_v | ~ptw_pte_flag_r & ptw_pte_flag_w | _ptw_complete_T_4 | ptw_level == 2'h0; // @[CachePortProxy.scala 53:96]
  wire  _T_1 = io_in_req_ready & io_in_req_valid; // @[Decoupled.scala 51:35]
  wire  _T_2 = ~tlb_io_hit; // @[CachePortProxy.scala 59:24]
  wire [2:0] _GEN_20 = _GEN_7 & ~tlb_io_hit ? 3'h1 : state; // @[CachePortProxy.scala 59:37 60:17 21:93]
  wire [2:0] _GEN_21 = _T_1 ? _GEN_20 : state; // @[CachePortProxy.scala 58:28 21:93]
  wire  _T_7 = io_ptw_req_ready & io_ptw_req_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _ptw_level_T_1 = ptw_level - 2'h1; // @[CachePortProxy.scala 81:34]
  wire [2:0] _GEN_25 = ptw_complete ? 3'h3 : 3'h1; // @[CachePortProxy.scala 77:28 78:17 80:21]
  wire [1:0] _GEN_26 = ptw_complete ? ptw_level : _ptw_level_T_1; // @[CachePortProxy.scala 77:28 50:29 81:21]
  wire [2:0] _GEN_27 = _ptw_pte_reg_T ? _GEN_25 : state; // @[CachePortProxy.scala 76:30 21:93]
  wire [1:0] _GEN_28 = _ptw_pte_reg_T ? _GEN_26 : ptw_level; // @[CachePortProxy.scala 50:29 76:30]
  wire  _T_11 = io_out_req_ready & io_out_req_valid; // @[Decoupled.scala 51:35]
  wire  pte_flag_v = _in_req_bits_T ? tlb_io_rpte_flag_v : ptw_pte_reg_flag_v; // @[CachePortProxy.scala 121:18]
  wire  pte_flag_r = _in_req_bits_T ? tlb_io_rpte_flag_r : ptw_pte_reg_flag_r; // @[CachePortProxy.scala 121:18]
  wire  pte_flag_w = _in_req_bits_T ? tlb_io_rpte_flag_w : ptw_pte_reg_flag_w; // @[CachePortProxy.scala 121:18]
  wire  pf1 = ~pte_flag_v | ~pte_flag_r & pte_flag_w; // @[CachePortProxy.scala 136:20]
  wire  pte_flag_x = _in_req_bits_T ? tlb_io_rpte_flag_x : ptw_pte_reg_flag_x; // @[CachePortProxy.scala 121:18]
  wire  _T_19 = pte_flag_r | pte_flag_x; // @[CachePortProxy.scala 7:37]
  wire  pte_flag_a = _in_req_bits_T ? tlb_io_rpte_flag_a : ptw_pte_reg_flag_a; // @[CachePortProxy.scala 121:18]
  wire  _T_20 = ~pte_flag_a; // @[CachePortProxy.scala 140:10]
  wire  pf2 = _T_19 & _T_20; // @[CachePortProxy.scala 139:21 132:24]
  reg [1:0] prv_r; // @[Reg.scala 35:20]
  wire [1:0] prv = _in_req_bits_T ? io_prv : prv_r; // @[Utils.scala 50:8]
  wire  pte_flag_u = _in_req_bits_T ? tlb_io_rpte_flag_u : ptw_pte_reg_flag_u; // @[CachePortProxy.scala 121:18]
  wire  _T_23 = prv == 2'h0 & ~pte_flag_u; // @[CachePortProxy.scala 143:26]
  wire  pf3 = _T_19 & _T_23; // @[CachePortProxy.scala 139:21 133:24]
  wire  _T_24 = ~pte_flag_x; // @[CachePortProxy.scala 147:12]
  wire  pf4 = _T_19 & _T_24; // @[CachePortProxy.scala 139:21 134:24]
  wire  _T_25 = state == 3'h3; // @[CachePortProxy.scala 156:16]
  wire [8:0] pte_ppn1 = _in_req_bits_T ? tlb_io_rpte_ppn1 : ptw_pte_reg_ppn1; // @[CachePortProxy.scala 121:18]
  wire [8:0] pte_ppn0 = _in_req_bits_T ? tlb_io_rpte_ppn0 : ptw_pte_reg_ppn0; // @[CachePortProxy.scala 121:18]
  wire [17:0] _T_27 = {pte_ppn1,pte_ppn0}; // @[Cat.scala 33:92]
  wire  _T_33 = ptw_level == 2'h2 & _T_27 != 18'h0 | ptw_level == 2'h1 & pte_ppn0 != 9'h0; // @[CachePortProxy.scala 157:67]
  wire  _GEN_45 = state == 3'h3 & _T_33; // @[CachePortProxy.scala 135:24 156:36]
  wire  pf5 = _T_19 & _GEN_45; // @[CachePortProxy.scala 139:21 135:24]
  wire  page_fault = pf1 | pf2 | pf3 | pf4 | pf5; // @[CachePortProxy.scala 162:42]
  wire [2:0] _GEN_29 = _T_11 | page_fault ? 3'h0 : state; // @[CachePortProxy.scala 86:43 87:15 21:93]
  wire  _T_14 = io_in_resp_ready & io_in_resp_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_30 = _T_14 ? 3'h0 : state; // @[CachePortProxy.scala 91:29 92:15 21:93]
  wire [2:0] _GEN_31 = 3'h4 == state ? _GEN_30 : state; // @[CachePortProxy.scala 56:17 21:93]
  wire [2:0] _GEN_32 = 3'h3 == state ? _GEN_29 : _GEN_31; // @[CachePortProxy.scala 56:17]
  wire [55:0] _l2_addr_T = {io_satp_ppn,in_vaddr_vpn2,3'h0}; // @[Cat.scala 33:92]
  wire [31:0] l1_addr = {ptw_pte_reg_ppn2,ptw_pte_reg_ppn1,ptw_pte_reg_ppn0,in_vaddr_vpn1,3'h0}; // @[Cat.scala 33:92]
  wire [31:0] l0_addr = {ptw_pte_reg_ppn2,ptw_pte_reg_ppn1,ptw_pte_reg_ppn0,in_vaddr_vpn0,3'h0}; // @[Cat.scala 33:92]
  wire [31:0] l2_addr = _l2_addr_T[31:0]; // @[CachePortProxy.scala 102:11 98:21]
  wire [31:0] _io_ptw_req_bits_addr_T_1 = 2'h2 == ptw_level ? l2_addr : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] _io_ptw_req_bits_addr_T_3 = 2'h1 == ptw_level ? l1_addr : _io_ptw_req_bits_addr_T_1; // @[Mux.scala 81:58]
  wire [31:0] _io_ptw_req_bits_addr_T_5 = 2'h0 == ptw_level ? l0_addr : _io_ptw_req_bits_addr_T_3; // @[Mux.scala 81:58]
  wire [1:0] pte_ppn2 = _in_req_bits_T ? tlb_io_rpte_ppn2 : ptw_pte_reg_ppn2; // @[CachePortProxy.scala 121:18]
  wire [1:0] level = _in_req_bits_T ? tlb_io_rlevel : ptw_level; // @[CachePortProxy.scala 122:18]
  wire  _tlb_io_wen_T_1 = ~page_fault; // @[CachePortProxy.scala 125:50]
  wire  _tlb_io_wen_T_2 = _T_25 & ~page_fault; // @[CachePortProxy.scala 125:47]
  wire [8:0] paddr_ppn0 = level > 2'h0 ? in_vaddr_vpn0 : pte_ppn0; // @[CachePortProxy.scala 167:22]
  wire [8:0] paddr_ppn1 = level > 2'h1 ? in_vaddr_vpn1 : pte_ppn1; // @[CachePortProxy.scala 168:22]
  wire [31:0] _io_out_req_bits_addr_T = {pte_ppn2,paddr_ppn1,paddr_ppn0,in_vaddr_offset}; // @[CachePortProxy.scala 177:43]
  wire [38:0] _io_out_req_bits_addr_WIRE = {{7'd0}, _io_out_req_bits_addr_T}; // @[CachePortProxy.scala 177:{43,43}]
  wire  _page_fault_reg_T_7 = page_fault & _GEN_7 & (_in_req_bits_T & tlb_io_hit & _T_1 | _T_25); // @[CachePortProxy.scala 182:26]
  reg  page_fault_reg; // @[Utils.scala 36:20]
  wire  _GEN_51 = _page_fault_reg_T_7 | page_fault_reg; // @[Utils.scala 41:19 36:20 41:23]
  TLB tlb ( // @[CachePortProxy.scala 28:19]
    .clock(tlb_clock),
    .reset(tlb_reset),
    .io_sfence_vma(tlb_io_sfence_vma),
    .io_vaddr_vpn2(tlb_io_vaddr_vpn2),
    .io_vaddr_vpn1(tlb_io_vaddr_vpn1),
    .io_vaddr_vpn0(tlb_io_vaddr_vpn0),
    .io_rpte_ppn2(tlb_io_rpte_ppn2),
    .io_rpte_ppn1(tlb_io_rpte_ppn1),
    .io_rpte_ppn0(tlb_io_rpte_ppn0),
    .io_rpte_flag_d(tlb_io_rpte_flag_d),
    .io_rpte_flag_a(tlb_io_rpte_flag_a),
    .io_rpte_flag_u(tlb_io_rpte_flag_u),
    .io_rpte_flag_x(tlb_io_rpte_flag_x),
    .io_rpte_flag_w(tlb_io_rpte_flag_w),
    .io_rpte_flag_r(tlb_io_rpte_flag_r),
    .io_rpte_flag_v(tlb_io_rpte_flag_v),
    .io_rlevel(tlb_io_rlevel),
    .io_hit(tlb_io_hit),
    .io_wen(tlb_io_wen),
    .io_wvaddr_vpn2(tlb_io_wvaddr_vpn2),
    .io_wvaddr_vpn1(tlb_io_wvaddr_vpn1),
    .io_wvaddr_vpn0(tlb_io_wvaddr_vpn0),
    .io_wpte_ppn2(tlb_io_wpte_ppn2),
    .io_wpte_ppn1(tlb_io_wpte_ppn1),
    .io_wpte_ppn0(tlb_io_wpte_ppn0),
    .io_wpte_flag_d(tlb_io_wpte_flag_d),
    .io_wpte_flag_a(tlb_io_wpte_flag_a),
    .io_wpte_flag_g(tlb_io_wpte_flag_g),
    .io_wpte_flag_u(tlb_io_wpte_flag_u),
    .io_wpte_flag_x(tlb_io_wpte_flag_x),
    .io_wpte_flag_w(tlb_io_wpte_flag_w),
    .io_wpte_flag_r(tlb_io_wpte_flag_r),
    .io_wpte_flag_v(tlb_io_wpte_flag_v),
    .io_wlevel(tlb_io_wlevel),
    .io_satp_asid(tlb_io_satp_asid)
  );
  assign io_in_req_ready = _in_req_bits_T & (io_out_req_ready | access_fault | _GEN_7 & (_T_2 | page_fault)); // @[CachePortProxy.scala 172:41]
  assign io_in_resp_valid = io_out_resp_valid | io_in_resp_bits_page_fault | io_in_resp_bits_access_fault; // @[CachePortProxy.scala 189:83]
  assign io_in_resp_bits_rdata = io_out_resp_bits_rdata; // @[CachePortProxy.scala 185:32]
  assign io_in_resp_bits_page_fault = page_fault_reg; // @[CachePortProxy.scala 186:32]
  assign io_in_resp_bits_access_fault = state == 3'h4; // @[CachePortProxy.scala 187:42]
  assign io_out_req_valid = _in_req_bits_T & (tlb_io_hit & _tlb_io_wen_T_1 | _access_fault_T_3 & ~access_fault) &
    io_in_req_valid | _tlb_io_wen_T_2; // @[CachePortProxy.scala 173:126]
  assign io_out_req_bits_addr = _GEN_7 ? _io_out_req_bits_addr_WIRE : _GEN_0; // @[CachePortProxy.scala 176:16 175:19 177:26]
  assign io_out_resp_ready = io_in_resp_ready; // @[CachePortProxy.scala 190:32]
  assign io_ptw_req_valid = state == 3'h1; // @[CachePortProxy.scala 117:31]
  assign io_ptw_req_bits_addr = {{7'd0}, _io_ptw_req_bits_addr_T_5}; // @[CachePortProxy.scala 108:24]
  assign io_ptw_resp_ready = state == 3'h2; // @[CachePortProxy.scala 118:31]
  assign tlb_clock = clock;
  assign tlb_reset = reset;
  assign tlb_io_sfence_vma = io_sfence_vma; // @[CachePortProxy.scala 31:21]
  assign tlb_io_vaddr_vpn2 = io_in_req_bits_addr[38:30]; // @[CachePortProxy.scala 32:52]
  assign tlb_io_vaddr_vpn1 = io_in_req_bits_addr[29:21]; // @[CachePortProxy.scala 32:52]
  assign tlb_io_vaddr_vpn0 = io_in_req_bits_addr[20:12]; // @[CachePortProxy.scala 32:52]
  assign tlb_io_wen = _T_25 & ~page_fault; // @[CachePortProxy.scala 125:47]
  assign tlb_io_wvaddr_vpn2 = _GEN_0[38:30]; // @[CachePortProxy.scala 25:46]
  assign tlb_io_wvaddr_vpn1 = _GEN_0[29:21]; // @[CachePortProxy.scala 25:46]
  assign tlb_io_wvaddr_vpn0 = _GEN_0[20:12]; // @[CachePortProxy.scala 25:46]
  assign tlb_io_wpte_ppn2 = ptw_pte_reg_ppn2; // @[CachePortProxy.scala 127:17]
  assign tlb_io_wpte_ppn1 = ptw_pte_reg_ppn1; // @[CachePortProxy.scala 127:17]
  assign tlb_io_wpte_ppn0 = ptw_pte_reg_ppn0; // @[CachePortProxy.scala 127:17]
  assign tlb_io_wpte_flag_d = ptw_pte_reg_flag_d; // @[CachePortProxy.scala 127:17]
  assign tlb_io_wpte_flag_a = ptw_pte_reg_flag_a; // @[CachePortProxy.scala 127:17]
  assign tlb_io_wpte_flag_g = ptw_pte_reg_flag_g; // @[CachePortProxy.scala 127:17]
  assign tlb_io_wpte_flag_u = ptw_pte_reg_flag_u; // @[CachePortProxy.scala 127:17]
  assign tlb_io_wpte_flag_x = ptw_pte_reg_flag_x; // @[CachePortProxy.scala 127:17]
  assign tlb_io_wpte_flag_w = ptw_pte_reg_flag_w; // @[CachePortProxy.scala 127:17]
  assign tlb_io_wpte_flag_r = ptw_pte_reg_flag_r; // @[CachePortProxy.scala 127:17]
  assign tlb_io_wpte_flag_v = ptw_pte_reg_flag_v; // @[CachePortProxy.scala 127:17]
  assign tlb_io_wlevel = ptw_level; // @[CachePortProxy.scala 128:17]
  assign tlb_io_satp_asid = io_satp_asid; // @[CachePortProxy.scala 30:21]
  always @(posedge clock) begin
    if (reset) begin // @[CachePortProxy.scala 21:93]
      state <= 3'h0; // @[CachePortProxy.scala 21:93]
    end else if (3'h0 == state) begin // @[CachePortProxy.scala 56:17]
      if (io_in_req_valid) begin // @[CachePortProxy.scala 63:29]
        if (_access_fault_T_3 & access_fault) begin // @[CachePortProxy.scala 64:39]
          state <= 3'h4; // @[CachePortProxy.scala 65:17]
        end else begin
          state <= _GEN_21;
        end
      end else begin
        state <= _GEN_21;
      end
    end else if (3'h1 == state) begin // @[CachePortProxy.scala 56:17]
      if (_T_7) begin // @[CachePortProxy.scala 71:29]
        state <= 3'h2; // @[CachePortProxy.scala 72:15]
      end
    end else if (3'h2 == state) begin // @[CachePortProxy.scala 56:17]
      state <= _GEN_27;
    end else begin
      state <= _GEN_32;
    end
    if (reset) begin // @[Reg.scala 35:20]
      in_req_bits_r_addr <= 39'h0; // @[Reg.scala 35:20]
    end else if (_in_req_bits_T) begin // @[Reg.scala 36:18]
      in_req_bits_r_addr <= io_in_req_bits_addr; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      atp_en_r <= 1'h0; // @[Reg.scala 35:20]
    end else if (_in_req_bits_T) begin // @[Reg.scala 36:18]
      atp_en_r <= _atp_en_T_1; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[CachePortProxy.scala 50:29]
      ptw_level <= 2'h0; // @[CachePortProxy.scala 50:29]
    end else if (3'h0 == state) begin // @[CachePortProxy.scala 56:17]
      ptw_level <= 2'h2; // @[CachePortProxy.scala 68:17]
    end else if (!(3'h1 == state)) begin // @[CachePortProxy.scala 56:17]
      if (3'h2 == state) begin // @[CachePortProxy.scala 56:17]
        ptw_level <= _GEN_28;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      ptw_pte_reg_ppn2 <= 2'h0; // @[Reg.scala 35:20]
    end else if (_ptw_pte_reg_T) begin // @[Reg.scala 36:18]
      ptw_pte_reg_ppn2 <= ptw_pte_ppn2; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ptw_pte_reg_ppn1 <= 9'h0; // @[Reg.scala 35:20]
    end else if (_ptw_pte_reg_T) begin // @[Reg.scala 36:18]
      ptw_pte_reg_ppn1 <= ptw_pte_ppn1; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ptw_pte_reg_ppn0 <= 9'h0; // @[Reg.scala 35:20]
    end else if (_ptw_pte_reg_T) begin // @[Reg.scala 36:18]
      ptw_pte_reg_ppn0 <= ptw_pte_ppn0; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ptw_pte_reg_flag_d <= 1'h0; // @[Reg.scala 35:20]
    end else if (_ptw_pte_reg_T) begin // @[Reg.scala 36:18]
      ptw_pte_reg_flag_d <= ptw_pte_flag_d; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ptw_pte_reg_flag_a <= 1'h0; // @[Reg.scala 35:20]
    end else if (_ptw_pte_reg_T) begin // @[Reg.scala 36:18]
      ptw_pte_reg_flag_a <= ptw_pte_flag_a; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ptw_pte_reg_flag_g <= 1'h0; // @[Reg.scala 35:20]
    end else if (_ptw_pte_reg_T) begin // @[Reg.scala 36:18]
      ptw_pte_reg_flag_g <= ptw_pte_flag_g; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ptw_pte_reg_flag_u <= 1'h0; // @[Reg.scala 35:20]
    end else if (_ptw_pte_reg_T) begin // @[Reg.scala 36:18]
      ptw_pte_reg_flag_u <= ptw_pte_flag_u; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ptw_pte_reg_flag_x <= 1'h0; // @[Reg.scala 35:20]
    end else if (_ptw_pte_reg_T) begin // @[Reg.scala 36:18]
      ptw_pte_reg_flag_x <= ptw_pte_flag_x; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ptw_pte_reg_flag_w <= 1'h0; // @[Reg.scala 35:20]
    end else if (_ptw_pte_reg_T) begin // @[Reg.scala 36:18]
      ptw_pte_reg_flag_w <= ptw_pte_flag_w; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ptw_pte_reg_flag_r <= 1'h0; // @[Reg.scala 35:20]
    end else if (_ptw_pte_reg_T) begin // @[Reg.scala 36:18]
      ptw_pte_reg_flag_r <= ptw_pte_flag_r; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ptw_pte_reg_flag_v <= 1'h0; // @[Reg.scala 35:20]
    end else if (_ptw_pte_reg_T) begin // @[Reg.scala 36:18]
      ptw_pte_reg_flag_v <= ptw_pte_flag_v; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      prv_r <= 2'h0; // @[Reg.scala 35:20]
    end else if (_in_req_bits_T) begin // @[Utils.scala 50:8]
      prv_r <= io_prv;
    end
    if (reset) begin // @[Utils.scala 36:20]
      page_fault_reg <= 1'h0; // @[Utils.scala 36:20]
    end else if (_T_14) begin // @[Utils.scala 42:18]
      page_fault_reg <= 1'h0; // @[Utils.scala 42:22]
    end else begin
      page_fault_reg <= _GEN_51;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {2{`RANDOM}};
  in_req_bits_r_addr = _RAND_1[38:0];
  _RAND_2 = {1{`RANDOM}};
  atp_en_r = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  ptw_level = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  ptw_pte_reg_ppn2 = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  ptw_pte_reg_ppn1 = _RAND_5[8:0];
  _RAND_6 = {1{`RANDOM}};
  ptw_pte_reg_ppn0 = _RAND_6[8:0];
  _RAND_7 = {1{`RANDOM}};
  ptw_pte_reg_flag_d = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  ptw_pte_reg_flag_a = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  ptw_pte_reg_flag_g = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  ptw_pte_reg_flag_u = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  ptw_pte_reg_flag_x = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  ptw_pte_reg_flag_w = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  ptw_pte_reg_flag_r = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  ptw_pte_reg_flag_v = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  prv_r = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  page_fault_reg = _RAND_16[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_2(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [63:0] io_enq_bits_pc,
  input  [31:0] io_enq_bits_instr,
  input         io_enq_bits_page_fault,
  input         io_enq_bits_access_fault,
  input  [63:0] io_enq_bits_bp_npc,
  input         io_deq_ready,
  output        io_deq_valid,
  output [63:0] io_deq_bits_pc,
  output [31:0] io_deq_bits_instr,
  output        io_deq_bits_page_fault,
  output        io_deq_bits_access_fault,
  output [63:0] io_deq_bits_bp_npc,
  input         io_flush
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] ram_pc [0:3]; // @[Decoupled.scala 273:95]
  wire  ram_pc_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire [1:0] ram_pc_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [63:0] ram_pc_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [63:0] ram_pc_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_pc_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_pc_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_pc_MPORT_en; // @[Decoupled.scala 273:95]
  reg [31:0] ram_instr [0:3]; // @[Decoupled.scala 273:95]
  wire  ram_instr_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire [1:0] ram_instr_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [31:0] ram_instr_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [31:0] ram_instr_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_instr_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_instr_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_instr_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_page_fault [0:3]; // @[Decoupled.scala 273:95]
  wire  ram_page_fault_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire [1:0] ram_page_fault_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_page_fault_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_page_fault_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_page_fault_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_page_fault_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_page_fault_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_access_fault [0:3]; // @[Decoupled.scala 273:95]
  wire  ram_access_fault_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire [1:0] ram_access_fault_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_access_fault_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_access_fault_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_access_fault_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_access_fault_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_access_fault_MPORT_en; // @[Decoupled.scala 273:95]
  reg [63:0] ram_bp_npc [0:3]; // @[Decoupled.scala 273:95]
  wire  ram_bp_npc_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire [1:0] ram_bp_npc_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [63:0] ram_bp_npc_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [63:0] ram_bp_npc_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_bp_npc_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_bp_npc_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_bp_npc_MPORT_en; // @[Decoupled.scala 273:95]
  reg [1:0] enq_ptr_value; // @[Counter.scala 61:40]
  reg [1:0] deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _value_T_1 = enq_ptr_value + 2'h1; // @[Counter.scala 77:24]
  wire [1:0] _value_T_3 = deq_ptr_value + 2'h1; // @[Counter.scala 77:24]
  assign ram_pc_io_deq_bits_MPORT_en = 1'h1;
  assign ram_pc_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_pc_io_deq_bits_MPORT_data = ram_pc[ram_pc_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_pc_MPORT_data = io_enq_bits_pc;
  assign ram_pc_MPORT_addr = enq_ptr_value;
  assign ram_pc_MPORT_mask = 1'h1;
  assign ram_pc_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_instr_io_deq_bits_MPORT_en = 1'h1;
  assign ram_instr_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_instr_io_deq_bits_MPORT_data = ram_instr[ram_instr_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_instr_MPORT_data = io_enq_bits_instr;
  assign ram_instr_MPORT_addr = enq_ptr_value;
  assign ram_instr_MPORT_mask = 1'h1;
  assign ram_instr_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_page_fault_io_deq_bits_MPORT_en = 1'h1;
  assign ram_page_fault_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_page_fault_io_deq_bits_MPORT_data = ram_page_fault[ram_page_fault_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_page_fault_MPORT_data = io_enq_bits_page_fault;
  assign ram_page_fault_MPORT_addr = enq_ptr_value;
  assign ram_page_fault_MPORT_mask = 1'h1;
  assign ram_page_fault_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_access_fault_io_deq_bits_MPORT_en = 1'h1;
  assign ram_access_fault_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_access_fault_io_deq_bits_MPORT_data = ram_access_fault[ram_access_fault_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_access_fault_MPORT_data = io_enq_bits_access_fault;
  assign ram_access_fault_MPORT_addr = enq_ptr_value;
  assign ram_access_fault_MPORT_mask = 1'h1;
  assign ram_access_fault_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_bp_npc_io_deq_bits_MPORT_en = 1'h1;
  assign ram_bp_npc_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_bp_npc_io_deq_bits_MPORT_data = ram_bp_npc[ram_bp_npc_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_bp_npc_MPORT_data = io_enq_bits_bp_npc;
  assign ram_bp_npc_MPORT_addr = enq_ptr_value;
  assign ram_bp_npc_MPORT_mask = 1'h1;
  assign ram_bp_npc_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = io_deq_ready | ~full; // @[Decoupled.scala 303:16 323:{24,39}]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits_pc = ram_pc_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_instr = ram_instr_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_page_fault = ram_page_fault_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_access_fault = ram_access_fault_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_bp_npc = ram_bp_npc_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  always @(posedge clock) begin
    if (ram_pc_MPORT_en & ram_pc_MPORT_mask) begin
      ram_pc[ram_pc_MPORT_addr] <= ram_pc_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_instr_MPORT_en & ram_instr_MPORT_mask) begin
      ram_instr[ram_instr_MPORT_addr] <= ram_instr_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_page_fault_MPORT_en & ram_page_fault_MPORT_mask) begin
      ram_page_fault[ram_page_fault_MPORT_addr] <= ram_page_fault_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_access_fault_MPORT_en & ram_access_fault_MPORT_mask) begin
      ram_access_fault[ram_access_fault_MPORT_addr] <= ram_access_fault_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_bp_npc_MPORT_en & ram_bp_npc_MPORT_mask) begin
      ram_bp_npc[ram_bp_npc_MPORT_addr] <= ram_bp_npc_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 2'h0; // @[Counter.scala 61:40]
    end else if (io_flush) begin // @[Decoupled.scala 296:15]
      enq_ptr_value <= 2'h0; // @[Counter.scala 98:11]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 2'h0; // @[Counter.scala 61:40]
    end else if (io_flush) begin // @[Decoupled.scala 296:15]
      deq_ptr_value <= 2'h0; // @[Counter.scala 98:11]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (io_flush) begin // @[Decoupled.scala 296:15]
      maybe_full <= 1'h0; // @[Decoupled.scala 299:16]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_pc[initvar] = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_instr[initvar] = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_page_fault[initvar] = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_access_fault[initvar] = _RAND_3[0:0];
  _RAND_4 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_bp_npc[initvar] = _RAND_4[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  enq_ptr_value = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  deq_ptr_value = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  maybe_full = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Decode(
  input  [63:0] io_in_pc,
  input  [31:0] io_in_instr,
  input         io_in_valid,
  input         io_in_page_fault,
  input         io_in_access_fault,
  output        io_out_valid,
  output [2:0]  io_out_exc,
  output [63:0] io_out_pc,
  output [63:0] io_out_npc,
  output [31:0] io_out_instr,
  output [2:0]  io_out_fu,
  output [3:0]  io_out_alu_op,
  output [1:0]  io_out_jmp_op,
  output [3:0]  io_out_mdu_op,
  output [4:0]  io_out_lsu_op,
  output [1:0]  io_out_mem_len,
  output [1:0]  io_out_csr_op,
  output [2:0]  io_out_sys_op,
  output [1:0]  io_out_rs1_src,
  output [1:0]  io_out_rs2_src,
  output [4:0]  io_out_rs1_index,
  output [4:0]  io_out_rs2_index,
  output [4:0]  io_out_rd_index,
  output        io_out_rd_wen,
  output [31:0] io_out_imm,
  output        io_out_dw
);
  wire [63:0] uop_npc = io_in_pc + 64'h4; // @[Decode.scala 16:29]
  wire [4:0] uop_rs1_index = io_in_instr[19:15]; // @[Decode.scala 18:25]
  wire [4:0] uop_rs2_index = io_in_instr[24:20]; // @[Decode.scala 19:25]
  wire [4:0] uop_rd_index = io_in_instr[11:7]; // @[Decode.scala 20:25]
  wire [31:0] decode_result_invInputs = ~io_in_instr; // @[pla.scala 78:21]
  wire  decode_result_andMatrixInput_0 = decode_result_invInputs[2]; // @[pla.scala 91:29]
  wire  decode_result_andMatrixInput_1 = decode_result_invInputs[5]; // @[pla.scala 91:29]
  wire [1:0] _decode_result_T = {decode_result_andMatrixInput_0,decode_result_andMatrixInput_1}; // @[Cat.scala 33:92]
  wire  _decode_result_T_1 = &_decode_result_T; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_1_1 = decode_result_invInputs[4]; // @[pla.scala 91:29]
  wire [2:0] _decode_result_T_2 = {decode_result_andMatrixInput_0,decode_result_andMatrixInput_1_1,
    decode_result_andMatrixInput_1}; // @[Cat.scala 33:92]
  wire  _decode_result_T_3 = &_decode_result_T_2; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_1_2 = decode_result_invInputs[6]; // @[pla.scala 91:29]
  wire [1:0] _decode_result_T_4 = {decode_result_andMatrixInput_0,decode_result_andMatrixInput_1_2}; // @[Cat.scala 33:92]
  wire  _decode_result_T_5 = &_decode_result_T_4; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_0_3 = io_in_instr[0]; // @[pla.scala 90:45]
  wire  decode_result_andMatrixInput_1_3 = io_in_instr[1]; // @[pla.scala 90:45]
  wire  decode_result_andMatrixInput_3 = decode_result_invInputs[3]; // @[pla.scala 91:29]
  wire  decode_result_andMatrixInput_6 = decode_result_invInputs[12]; // @[pla.scala 91:29]
  wire [6:0] _decode_result_T_6 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3,decode_result_andMatrixInput_1,
    decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_6}; // @[Cat.scala 33:92]
  wire  _decode_result_T_7 = &_decode_result_T_6; // @[pla.scala 98:74]
  wire [7:0] _decode_result_T_8 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3,decode_result_andMatrixInput_1_1,
    decode_result_andMatrixInput_1,decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_6}; // @[Cat.scala 33:92]
  wire  _decode_result_T_9 = &_decode_result_T_8; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_7_1 = decode_result_invInputs[13]; // @[pla.scala 91:29]
  wire [7:0] _decode_result_T_10 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3,decode_result_andMatrixInput_1_1,
    decode_result_andMatrixInput_1,decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_7_1}; // @[Cat.scala 33:92]
  wire  _decode_result_T_11 = &_decode_result_T_10; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_6_3 = decode_result_invInputs[14]; // @[pla.scala 91:29]
  wire [6:0] _decode_result_T_12 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3,decode_result_andMatrixInput_1_1,
    decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_6_3}; // @[Cat.scala 33:92]
  wire  _decode_result_T_13 = &_decode_result_T_12; // @[pla.scala 98:74]
  wire [7:0] _decode_result_T_14 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3,decode_result_andMatrixInput_1_1,
    decode_result_andMatrixInput_1,decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_6_3}; // @[Cat.scala 33:92]
  wire  _decode_result_T_15 = &_decode_result_T_14; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_8 = decode_result_invInputs[25]; // @[pla.scala 91:29]
  wire  decode_result_andMatrixInput_9 = decode_result_invInputs[26]; // @[pla.scala 91:29]
  wire  decode_result_andMatrixInput_10 = decode_result_invInputs[27]; // @[pla.scala 91:29]
  wire  decode_result_andMatrixInput_11 = decode_result_invInputs[28]; // @[pla.scala 91:29]
  wire  decode_result_andMatrixInput_12 = decode_result_invInputs[29]; // @[pla.scala 91:29]
  wire  decode_result_andMatrixInput_13 = decode_result_invInputs[31]; // @[pla.scala 91:29]
  wire [6:0] decode_result_lo_5 = {decode_result_andMatrixInput_6_3,decode_result_andMatrixInput_8,
    decode_result_andMatrixInput_9,decode_result_andMatrixInput_10,decode_result_andMatrixInput_11,
    decode_result_andMatrixInput_12,decode_result_andMatrixInput_13}; // @[Cat.scala 33:92]
  wire [13:0] _decode_result_T_16 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3,decode_result_andMatrixInput_1_2,
    decode_result_andMatrixInput_6,decode_result_andMatrixInput_7_1,decode_result_lo_5}; // @[Cat.scala 33:92]
  wire  _decode_result_T_17 = &_decode_result_T_16; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_0_9 = io_in_instr[2]; // @[pla.scala 90:45]
  wire [2:0] _decode_result_T_18 = {decode_result_andMatrixInput_0_9,decode_result_andMatrixInput_3,
    decode_result_andMatrixInput_1_1}; // @[Cat.scala 33:92]
  wire  _decode_result_T_19 = &_decode_result_T_18; // @[pla.scala 98:74]
  wire [2:0] _decode_result_T_20 = {decode_result_andMatrixInput_0_9,decode_result_andMatrixInput_3,
    decode_result_andMatrixInput_1}; // @[Cat.scala 33:92]
  wire  _decode_result_T_21 = &_decode_result_T_20; // @[pla.scala 98:74]
  wire [2:0] _decode_result_T_22 = {decode_result_andMatrixInput_0_9,decode_result_andMatrixInput_1_1,
    decode_result_andMatrixInput_1}; // @[Cat.scala 33:92]
  wire  _decode_result_T_23 = &_decode_result_T_22; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_1_12 = io_in_instr[3]; // @[pla.scala 90:45]
  wire [1:0] _decode_result_T_24 = {decode_result_andMatrixInput_0,decode_result_andMatrixInput_1_12}; // @[Cat.scala 33:92]
  wire  _decode_result_T_25 = &_decode_result_T_24; // @[pla.scala 98:74]
  wire [8:0] _decode_result_T_26 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0_9,decode_result_andMatrixInput_1_12,decode_result_andMatrixInput_1_1,
    decode_result_andMatrixInput_1,decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_7_1,
    decode_result_andMatrixInput_6_3}; // @[Cat.scala 33:92]
  wire  _decode_result_T_27 = &_decode_result_T_26; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_3_7 = io_in_instr[4]; // @[pla.scala 90:45]
  wire [8:0] _decode_result_T_28 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3_7,decode_result_andMatrixInput_1,
    decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_6,decode_result_andMatrixInput_7_1,
    decode_result_andMatrixInput_6_3}; // @[Cat.scala 33:92]
  wire  _decode_result_T_29 = &_decode_result_T_28; // @[pla.scala 98:74]
  wire [13:0] _decode_result_T_30 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3_7,decode_result_andMatrixInput_1_2,
    decode_result_andMatrixInput_6,decode_result_andMatrixInput_7_1,decode_result_lo_5}; // @[Cat.scala 33:92]
  wire  _decode_result_T_31 = &_decode_result_T_30; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_9_2 = decode_result_invInputs[30]; // @[pla.scala 91:29]
  wire [4:0] decode_result_lo_9 = {decode_result_andMatrixInput_10,decode_result_andMatrixInput_11,
    decode_result_andMatrixInput_12,decode_result_andMatrixInput_9_2,decode_result_andMatrixInput_13}; // @[Cat.scala 33:92]
  wire [10:0] _decode_result_T_32 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_3,decode_result_andMatrixInput_3_7,decode_result_andMatrixInput_1_2,
    decode_result_andMatrixInput_9,decode_result_lo_9}; // @[Cat.scala 33:92]
  wire  _decode_result_T_33 = &_decode_result_T_32; // @[pla.scala 98:74]
  wire [1:0] _decode_result_T_34 = {decode_result_andMatrixInput_0_9,decode_result_andMatrixInput_3_7}; // @[Cat.scala 33:92]
  wire  _decode_result_T_35 = &_decode_result_T_34; // @[pla.scala 98:74]
  wire [5:0] _decode_result_T_36 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0_9,decode_result_andMatrixInput_3,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_1_2}; // @[Cat.scala 33:92]
  wire  _decode_result_T_37 = &_decode_result_T_36; // @[pla.scala 98:74]
  wire [9:0] _decode_result_T_38 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_1_12,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_1,decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_6,
    decode_result_andMatrixInput_7_1,decode_result_andMatrixInput_6_3}; // @[Cat.scala 33:92]
  wire  _decode_result_T_39 = &_decode_result_T_38; // @[pla.scala 98:74]
  wire [14:0] _decode_result_T_40 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_1_12,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_6,decode_result_andMatrixInput_7_1,decode_result_lo_5}
    ; // @[Cat.scala 33:92]
  wire  _decode_result_T_41 = &_decode_result_T_40; // @[pla.scala 98:74]
  wire [6:0] decode_result_lo_13 = {decode_result_andMatrixInput_6_3,decode_result_andMatrixInput_9,
    decode_result_andMatrixInput_10,decode_result_andMatrixInput_11,decode_result_andMatrixInput_12,
    decode_result_andMatrixInput_9_2,decode_result_andMatrixInput_13}; // @[Cat.scala 33:92]
  wire [14:0] _decode_result_T_42 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_1_12,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_6,decode_result_andMatrixInput_7_1,decode_result_lo_13
    }; // @[Cat.scala 33:92]
  wire  _decode_result_T_43 = &_decode_result_T_42; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_2_18 = io_in_instr[5]; // @[pla.scala 90:45]
  wire [3:0] _decode_result_T_44 = {decode_result_andMatrixInput_0,decode_result_andMatrixInput_1_1,
    decode_result_andMatrixInput_2_18,decode_result_andMatrixInput_1_2}; // @[Cat.scala 33:92]
  wire  _decode_result_T_45 = &_decode_result_T_44; // @[pla.scala 98:74]
  wire [4:0] _decode_result_T_46 = {decode_result_andMatrixInput_0_9,decode_result_andMatrixInput_1_12,
    decode_result_andMatrixInput_2_18,decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_11}; // @[Cat.scala 33:92]
  wire  _decode_result_T_47 = &_decode_result_T_46; // @[pla.scala 98:74]
  wire [8:0] _decode_result_T_48 = {decode_result_andMatrixInput_0_9,decode_result_andMatrixInput_1_12,
    decode_result_andMatrixInput_2_18,decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_10,
    decode_result_andMatrixInput_11,decode_result_andMatrixInput_12,decode_result_andMatrixInput_9_2,
    decode_result_andMatrixInput_13}; // @[Cat.scala 33:92]
  wire  _decode_result_T_49 = &_decode_result_T_48; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_3_17 = io_in_instr[6]; // @[pla.scala 90:45]
  wire [4:0] _decode_result_T_50 = {decode_result_andMatrixInput_0,decode_result_andMatrixInput_3,
    decode_result_andMatrixInput_1_1,decode_result_andMatrixInput_3_17,decode_result_andMatrixInput_6_3}; // @[Cat.scala 33:92]
  wire  _decode_result_T_51 = &_decode_result_T_50; // @[pla.scala 98:74]
  wire [2:0] _decode_result_T_52 = {decode_result_andMatrixInput_0_9,decode_result_andMatrixInput_1_12,
    decode_result_andMatrixInput_3_17}; // @[Cat.scala 33:92]
  wire  _decode_result_T_53 = &_decode_result_T_52; // @[pla.scala 98:74]
  wire [1:0] _decode_result_T_54 = {decode_result_andMatrixInput_3_7,decode_result_andMatrixInput_3_17}; // @[Cat.scala 33:92]
  wire  _decode_result_T_55 = &_decode_result_T_54; // @[pla.scala 98:74]
  wire [7:0] _decode_result_T_56 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3,decode_result_andMatrixInput_1_1,
    decode_result_andMatrixInput_2_18,decode_result_andMatrixInput_3_17,decode_result_andMatrixInput_7_1}; // @[Cat.scala 33:92]
  wire  _decode_result_T_57 = &_decode_result_T_56; // @[pla.scala 98:74]
  wire [8:0] _decode_result_T_58 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_3,decode_result_andMatrixInput_1_1,decode_result_andMatrixInput_2_18,
    decode_result_andMatrixInput_3_17,decode_result_andMatrixInput_6,decode_result_andMatrixInput_7_1,
    decode_result_andMatrixInput_6_3}; // @[Cat.scala 33:92]
  wire  _decode_result_T_59 = &_decode_result_T_58; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_5_17 = decode_result_invInputs[7]; // @[pla.scala 91:29]
  wire  decode_result_andMatrixInput_6_16 = decode_result_invInputs[8]; // @[pla.scala 91:29]
  wire  decode_result_andMatrixInput_7_14 = decode_result_invInputs[9]; // @[pla.scala 91:29]
  wire  decode_result_andMatrixInput_8_10 = decode_result_invInputs[10]; // @[pla.scala 91:29]
  wire  decode_result_andMatrixInput_9_6 = decode_result_invInputs[11]; // @[pla.scala 91:29]
  wire  decode_result_andMatrixInput_13_4 = decode_result_invInputs[15]; // @[pla.scala 91:29]
  wire  decode_result_andMatrixInput_14_2 = decode_result_invInputs[16]; // @[pla.scala 91:29]
  wire  decode_result_andMatrixInput_15 = decode_result_invInputs[17]; // @[pla.scala 91:29]
  wire  decode_result_andMatrixInput_16 = decode_result_invInputs[18]; // @[pla.scala 91:29]
  wire  decode_result_andMatrixInput_17 = decode_result_invInputs[19]; // @[pla.scala 91:29]
  wire  decode_result_andMatrixInput_18 = decode_result_invInputs[20]; // @[pla.scala 91:29]
  wire  decode_result_andMatrixInput_19 = decode_result_invInputs[21]; // @[pla.scala 91:29]
  wire  decode_result_andMatrixInput_20 = decode_result_invInputs[22]; // @[pla.scala 91:29]
  wire  decode_result_andMatrixInput_21 = decode_result_invInputs[23]; // @[pla.scala 91:29]
  wire  decode_result_andMatrixInput_22 = decode_result_invInputs[24]; // @[pla.scala 91:29]
  wire [6:0] decode_result_lo_lo_14 = {decode_result_andMatrixInput_8,decode_result_andMatrixInput_9,
    decode_result_andMatrixInput_10,decode_result_andMatrixInput_11,decode_result_andMatrixInput_12,
    decode_result_andMatrixInput_9_2,decode_result_andMatrixInput_13}; // @[Cat.scala 33:92]
  wire [14:0] decode_result_lo_20 = {decode_result_andMatrixInput_15,decode_result_andMatrixInput_16,
    decode_result_andMatrixInput_17,decode_result_andMatrixInput_18,decode_result_andMatrixInput_19,
    decode_result_andMatrixInput_20,decode_result_andMatrixInput_21,decode_result_andMatrixInput_22,
    decode_result_lo_lo_14}; // @[Cat.scala 33:92]
  wire [6:0] decode_result_hi_lo_16 = {decode_result_andMatrixInput_8_10,decode_result_andMatrixInput_9_6,
    decode_result_andMatrixInput_6,decode_result_andMatrixInput_7_1,decode_result_andMatrixInput_6_3,
    decode_result_andMatrixInput_13_4,decode_result_andMatrixInput_14_2}; // @[Cat.scala 33:92]
  wire [29:0] _decode_result_T_60 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_1_1,decode_result_andMatrixInput_2_18,decode_result_andMatrixInput_3_17,
    decode_result_andMatrixInput_5_17,decode_result_andMatrixInput_6_16,decode_result_andMatrixInput_7_14,
    decode_result_hi_lo_16,decode_result_lo_20}; // @[Cat.scala 33:92]
  wire  _decode_result_T_61 = &_decode_result_T_60; // @[pla.scala 98:74]
  wire [8:0] _decode_result_T_62 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0_9,decode_result_andMatrixInput_1_1,decode_result_andMatrixInput_2_18,
    decode_result_andMatrixInput_3_17,decode_result_andMatrixInput_6,decode_result_andMatrixInput_7_1,
    decode_result_andMatrixInput_6_3}; // @[Cat.scala 33:92]
  wire  _decode_result_T_63 = &_decode_result_T_62; // @[pla.scala 98:74]
  wire [6:0] _decode_result_T_64 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0_9,decode_result_andMatrixInput_1_12,decode_result_andMatrixInput_1_1,
    decode_result_andMatrixInput_2_18,decode_result_andMatrixInput_3_17}; // @[Cat.scala 33:92]
  wire  _decode_result_T_65 = &_decode_result_T_64; // @[pla.scala 98:74]
  wire [14:0] decode_result_lo_23 = {decode_result_andMatrixInput_14_2,decode_result_andMatrixInput_15,
    decode_result_andMatrixInput_16,decode_result_andMatrixInput_17,decode_result_andMatrixInput_19,
    decode_result_andMatrixInput_20,decode_result_andMatrixInput_21,decode_result_andMatrixInput_22,
    decode_result_lo_lo_14}; // @[Cat.scala 33:92]
  wire [7:0] decode_result_hi_lo_19 = {decode_result_andMatrixInput_6_16,decode_result_andMatrixInput_7_14,
    decode_result_andMatrixInput_8_10,decode_result_andMatrixInput_9_6,decode_result_andMatrixInput_6,
    decode_result_andMatrixInput_7_1,decode_result_andMatrixInput_6_3,decode_result_andMatrixInput_13_4}; // @[Cat.scala 33:92]
  wire [30:0] _decode_result_T_66 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_2_18,decode_result_andMatrixInput_3_17,decode_result_andMatrixInput_5_17,
    decode_result_hi_lo_19,decode_result_lo_23}; // @[Cat.scala 33:92]
  wire  _decode_result_T_67 = &_decode_result_T_66; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_0_34 = io_in_instr[12]; // @[pla.scala 90:45]
  wire  _decode_result_T_68 = &decode_result_andMatrixInput_0_34; // @[pla.scala 98:74]
  wire [3:0] _decode_result_T_69 = {decode_result_andMatrixInput_0_9,decode_result_andMatrixInput_1_12,
    decode_result_andMatrixInput_1,decode_result_andMatrixInput_0_34}; // @[Cat.scala 33:92]
  wire  _decode_result_T_70 = &_decode_result_T_69; // @[pla.scala 98:74]
  wire [3:0] _decode_result_T_71 = {decode_result_andMatrixInput_0,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_0_34,decode_result_andMatrixInput_7_1}; // @[Cat.scala 33:92]
  wire  _decode_result_T_72 = &_decode_result_T_71; // @[pla.scala 98:74]
  wire [13:0] _decode_result_T_73 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3_7,decode_result_andMatrixInput_1_2,
    decode_result_andMatrixInput_0_34,decode_result_andMatrixInput_7_1,decode_result_lo_lo_14}; // @[Cat.scala 33:92]
  wire  _decode_result_T_74 = &_decode_result_T_73; // @[pla.scala 98:74]
  wire [14:0] _decode_result_T_75 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_1_12,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_0_34,decode_result_andMatrixInput_7_1,
    decode_result_lo_lo_14}; // @[Cat.scala 33:92]
  wire  _decode_result_T_76 = &_decode_result_T_75; // @[pla.scala 98:74]
  wire [2:0] _decode_result_T_77 = {decode_result_andMatrixInput_0,decode_result_andMatrixInput_3_17,
    decode_result_andMatrixInput_0_34}; // @[Cat.scala 33:92]
  wire  _decode_result_T_78 = &_decode_result_T_77; // @[pla.scala 98:74]
  wire [2:0] _decode_result_T_79 = {decode_result_andMatrixInput_3_7,decode_result_andMatrixInput_3_17,
    decode_result_andMatrixInput_0_34}; // @[Cat.scala 33:92]
  wire  _decode_result_T_80 = &_decode_result_T_79; // @[pla.scala 98:74]
  wire [7:0] _decode_result_T_81 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3,decode_result_andMatrixInput_2_18,
    decode_result_andMatrixInput_3_17,decode_result_andMatrixInput_0_34,decode_result_andMatrixInput_7_1}; // @[Cat.scala 33:92]
  wire  _decode_result_T_82 = &_decode_result_T_81; // @[pla.scala 98:74]
  wire [7:0] _decode_result_T_83 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_2_18,decode_result_andMatrixInput_3_17,decode_result_andMatrixInput_0_34}; // @[Cat.scala 33:92]
  wire  _decode_result_T_84 = &_decode_result_T_83; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_1_42 = io_in_instr[13]; // @[pla.scala 90:45]
  wire [1:0] _decode_result_T_85 = {decode_result_andMatrixInput_0,decode_result_andMatrixInput_1_42}; // @[Cat.scala 33:92]
  wire  _decode_result_T_86 = &_decode_result_T_85; // @[pla.scala 98:74]
  wire [3:0] _decode_result_T_87 = {decode_result_andMatrixInput_0,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_1_42,decode_result_andMatrixInput_6_3}; // @[Cat.scala 33:92]
  wire  _decode_result_T_88 = &_decode_result_T_87; // @[pla.scala 98:74]
  wire [6:0] _decode_result_T_89 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_3,decode_result_andMatrixInput_3_7,decode_result_andMatrixInput_1,
    decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_1_42}; // @[Cat.scala 33:92]
  wire  _decode_result_T_90 = &_decode_result_T_89; // @[pla.scala 98:74]
  wire [9:0] _decode_result_T_91 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0_9,decode_result_andMatrixInput_1_12,decode_result_andMatrixInput_1_1,
    decode_result_andMatrixInput_2_18,decode_result_andMatrixInput_1_42,decode_result_andMatrixInput_6_3,
    decode_result_andMatrixInput_10,decode_result_andMatrixInput_11}; // @[Cat.scala 33:92]
  wire  _decode_result_T_92 = &_decode_result_T_91; // @[pla.scala 98:74]
  wire [4:0] decode_result_lo_33 = {decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_1_42,
    decode_result_andMatrixInput_6_3,decode_result_andMatrixInput_10,decode_result_andMatrixInput_11}; // @[Cat.scala 33:92]
  wire [10:0] _decode_result_T_93 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0_9,decode_result_andMatrixInput_1_12,decode_result_andMatrixInput_1_1,
    decode_result_andMatrixInput_2_18,decode_result_lo_33}; // @[Cat.scala 33:92]
  wire  _decode_result_T_94 = &_decode_result_T_93; // @[pla.scala 98:74]
  wire [7:0] decode_result_lo_34 = {decode_result_andMatrixInput_18,decode_result_andMatrixInput_19,
    decode_result_andMatrixInput_20,decode_result_andMatrixInput_21,decode_result_andMatrixInput_22,
    decode_result_andMatrixInput_12,decode_result_andMatrixInput_9_2,decode_result_andMatrixInput_13}; // @[Cat.scala 33:92]
  wire [15:0] _decode_result_T_95 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0_9,decode_result_andMatrixInput_1_12,decode_result_andMatrixInput_1_1,
    decode_result_andMatrixInput_2_18,decode_result_andMatrixInput_1_42,decode_result_andMatrixInput_6_3,
    decode_result_lo_34}; // @[Cat.scala 33:92]
  wire  _decode_result_T_96 = &_decode_result_T_95; // @[pla.scala 98:74]
  wire [16:0] _decode_result_T_97 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0_9,decode_result_andMatrixInput_1_12,decode_result_andMatrixInput_1_1,
    decode_result_andMatrixInput_2_18,decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_1_42,
    decode_result_andMatrixInput_6_3,decode_result_lo_34}; // @[Cat.scala 33:92]
  wire  _decode_result_T_98 = &_decode_result_T_97; // @[pla.scala 98:74]
  wire [2:0] _decode_result_T_99 = {decode_result_andMatrixInput_3_7,decode_result_andMatrixInput_3_17,
    decode_result_andMatrixInput_1_42}; // @[Cat.scala 33:92]
  wire  _decode_result_T_100 = &_decode_result_T_99; // @[pla.scala 98:74]
  wire [7:0] _decode_result_T_101 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_2_18,decode_result_andMatrixInput_3_17,decode_result_andMatrixInput_1_42}; // @[Cat.scala 33:92]
  wire  _decode_result_T_102 = &_decode_result_T_101; // @[pla.scala 98:74]
  wire [3:0] _decode_result_T_103 = {decode_result_andMatrixInput_0,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_0_34,decode_result_andMatrixInput_1_42}; // @[Cat.scala 33:92]
  wire  _decode_result_T_104 = &_decode_result_T_103; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_2_46 = io_in_instr[14]; // @[pla.scala 90:45]
  wire [2:0] _decode_result_T_105 = {decode_result_andMatrixInput_1_1,decode_result_andMatrixInput_1,
    decode_result_andMatrixInput_2_46}; // @[Cat.scala 33:92]
  wire  _decode_result_T_106 = &_decode_result_T_105; // @[pla.scala 98:74]
  wire [3:0] _decode_result_T_107 = {decode_result_andMatrixInput_0,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_6,decode_result_andMatrixInput_2_46}; // @[Cat.scala 33:92]
  wire  _decode_result_T_108 = &_decode_result_T_107; // @[pla.scala 98:74]
  wire [3:0] _decode_result_T_109 = {decode_result_andMatrixInput_0,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_2_46,decode_result_andMatrixInput_9_2}; // @[Cat.scala 33:92]
  wire  _decode_result_T_110 = &_decode_result_T_109; // @[pla.scala 98:74]
  wire [5:0] decode_result_lo_40 = {decode_result_andMatrixInput_2_46,decode_result_andMatrixInput_9,
    decode_result_andMatrixInput_10,decode_result_andMatrixInput_11,decode_result_andMatrixInput_12,
    decode_result_andMatrixInput_13}; // @[Cat.scala 33:92]
  wire [11:0] _decode_result_T_111 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_3,decode_result_andMatrixInput_3_7,decode_result_andMatrixInput_1,
    decode_result_andMatrixInput_1_2,decode_result_lo_40}; // @[Cat.scala 33:92]
  wire  _decode_result_T_112 = &_decode_result_T_111; // @[pla.scala 98:74]
  wire [3:0] _decode_result_T_113 = {decode_result_andMatrixInput_0,decode_result_andMatrixInput_1_1,
    decode_result_andMatrixInput_2_18,decode_result_andMatrixInput_2_46}; // @[Cat.scala 33:92]
  wire  _decode_result_T_114 = &_decode_result_T_113; // @[pla.scala 98:74]
  wire [2:0] _decode_result_T_115 = {decode_result_andMatrixInput_3_7,decode_result_andMatrixInput_3_17,
    decode_result_andMatrixInput_2_46}; // @[Cat.scala 33:92]
  wire  _decode_result_T_116 = &_decode_result_T_115; // @[pla.scala 98:74]
  wire [7:0] _decode_result_T_117 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3,decode_result_andMatrixInput_1_1,
    decode_result_andMatrixInput_2_18,decode_result_andMatrixInput_3_17,decode_result_andMatrixInput_2_46}; // @[Cat.scala 33:92]
  wire  _decode_result_T_118 = &_decode_result_T_117; // @[pla.scala 98:74]
  wire [3:0] _decode_result_T_119 = {decode_result_andMatrixInput_0,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_0_34,decode_result_andMatrixInput_2_46}; // @[Cat.scala 33:92]
  wire  _decode_result_T_120 = &_decode_result_T_119; // @[pla.scala 98:74]
  wire [6:0] decode_result_lo_44 = {decode_result_andMatrixInput_2_46,decode_result_andMatrixInput_8,
    decode_result_andMatrixInput_9,decode_result_andMatrixInput_10,decode_result_andMatrixInput_11,
    decode_result_andMatrixInput_12,decode_result_andMatrixInput_13}; // @[Cat.scala 33:92]
  wire [13:0] _decode_result_T_121 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3_7,decode_result_andMatrixInput_1_2,
    decode_result_andMatrixInput_0_34,decode_result_andMatrixInput_7_1,decode_result_lo_44}; // @[Cat.scala 33:92]
  wire  _decode_result_T_122 = &_decode_result_T_121; // @[pla.scala 98:74]
  wire [14:0] _decode_result_T_123 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_1_12,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_0_34,decode_result_andMatrixInput_7_1,
    decode_result_lo_44}; // @[Cat.scala 33:92]
  wire  _decode_result_T_124 = &_decode_result_T_123; // @[pla.scala 98:74]
  wire [3:0] _decode_result_T_125 = {decode_result_andMatrixInput_0,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_1_42,decode_result_andMatrixInput_2_46}; // @[Cat.scala 33:92]
  wire  _decode_result_T_126 = &_decode_result_T_125; // @[pla.scala 98:74]
  wire [3:0] _decode_result_T_127 = {decode_result_andMatrixInput_0,decode_result_andMatrixInput_2_18,
    decode_result_andMatrixInput_1_42,decode_result_andMatrixInput_2_46}; // @[Cat.scala 33:92]
  wire  _decode_result_T_128 = &_decode_result_T_127; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_20_2 = io_in_instr[20]; // @[pla.scala 90:45]
  wire [7:0] decode_result_lo_lo_30 = {decode_result_andMatrixInput_22,decode_result_andMatrixInput_8,
    decode_result_andMatrixInput_9,decode_result_andMatrixInput_10,decode_result_andMatrixInput_11,
    decode_result_andMatrixInput_12,decode_result_andMatrixInput_9_2,decode_result_andMatrixInput_13}; // @[Cat.scala 33:92]
  wire [15:0] decode_result_lo_48 = {decode_result_andMatrixInput_14_2,decode_result_andMatrixInput_15,
    decode_result_andMatrixInput_16,decode_result_andMatrixInput_17,decode_result_andMatrixInput_20_2,
    decode_result_andMatrixInput_19,decode_result_andMatrixInput_20,decode_result_andMatrixInput_21,
    decode_result_lo_lo_30}; // @[Cat.scala 33:92]
  wire [31:0] _decode_result_T_129 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_2_18,decode_result_andMatrixInput_3_17,decode_result_andMatrixInput_5_17,
    decode_result_hi_lo_19,decode_result_lo_48}; // @[Cat.scala 33:92]
  wire  _decode_result_T_130 = &_decode_result_T_129; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_4_38 = io_in_instr[21]; // @[pla.scala 90:45]
  wire [5:0] _decode_result_T_131 = {decode_result_andMatrixInput_3_7,decode_result_andMatrixInput_3_17,
    decode_result_andMatrixInput_6,decode_result_andMatrixInput_7_1,decode_result_andMatrixInput_4_38,
    decode_result_andMatrixInput_12}; // @[Cat.scala 33:92]
  wire  _decode_result_T_132 = &_decode_result_T_131; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_7_31 = io_in_instr[25]; // @[pla.scala 90:45]
  wire [6:0] decode_result_lo_50 = {decode_result_andMatrixInput_7_31,decode_result_andMatrixInput_9,
    decode_result_andMatrixInput_10,decode_result_andMatrixInput_11,decode_result_andMatrixInput_12,
    decode_result_andMatrixInput_9_2,decode_result_andMatrixInput_13}; // @[Cat.scala 33:92]
  wire [13:0] _decode_result_T_133 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_2_18,decode_result_andMatrixInput_1_2,decode_result_lo_50}; // @[Cat.scala 33:92]
  wire  _decode_result_T_134 = &_decode_result_T_133; // @[pla.scala 98:74]
  wire [14:0] _decode_result_T_135 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3_7,decode_result_andMatrixInput_2_18,
    decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_6,decode_result_andMatrixInput_7_1,decode_result_lo_50
    }; // @[Cat.scala 33:92]
  wire  _decode_result_T_136 = &_decode_result_T_135; // @[pla.scala 98:74]
  wire [4:0] _decode_result_T_137 = {decode_result_andMatrixInput_3_7,decode_result_andMatrixInput_3_17,
    decode_result_andMatrixInput_6,decode_result_andMatrixInput_7_1,decode_result_andMatrixInput_7_31}; // @[Cat.scala 33:92]
  wire  _decode_result_T_138 = &_decode_result_T_137; // @[pla.scala 98:74]
  wire [13:0] _decode_result_T_139 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3_7,decode_result_andMatrixInput_2_18,
    decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_2_46,decode_result_lo_50}; // @[Cat.scala 33:92]
  wire  _decode_result_T_140 = &_decode_result_T_139; // @[pla.scala 98:74]
  wire [14:0] _decode_result_T_141 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_1_12,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_2_18,decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_2_46,
    decode_result_lo_50}; // @[Cat.scala 33:92]
  wire  _decode_result_T_142 = &_decode_result_T_141; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_3_55 = io_in_instr[27]; // @[pla.scala 90:45]
  wire [3:0] _decode_result_T_143 = {decode_result_andMatrixInput_1_12,decode_result_andMatrixInput_2_18,
    decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_3_55}; // @[Cat.scala 33:92]
  wire  _decode_result_T_144 = &_decode_result_T_143; // @[pla.scala 98:74]
  wire [4:0] _decode_result_T_145 = {decode_result_andMatrixInput_1_12,decode_result_andMatrixInput_2_18,
    decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_3_55,decode_result_andMatrixInput_11}; // @[Cat.scala 33:92]
  wire  _decode_result_T_146 = &_decode_result_T_145; // @[pla.scala 98:74]
  wire [5:0] decode_result_lo_57 = {decode_result_andMatrixInput_1_42,decode_result_andMatrixInput_6_3,
    decode_result_andMatrixInput_3_55,decode_result_andMatrixInput_12,decode_result_andMatrixInput_9_2,
    decode_result_andMatrixInput_13}; // @[Cat.scala 33:92]
  wire [11:0] _decode_result_T_147 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0_9,decode_result_andMatrixInput_1_12,decode_result_andMatrixInput_1_1,
    decode_result_andMatrixInput_2_18,decode_result_lo_57}; // @[Cat.scala 33:92]
  wire  _decode_result_T_148 = &_decode_result_T_147; // @[pla.scala 98:74]
  wire [12:0] _decode_result_T_149 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0_9,decode_result_andMatrixInput_1_12,decode_result_andMatrixInput_1_1,
    decode_result_andMatrixInput_2_18,decode_result_andMatrixInput_1_2,decode_result_lo_57}; // @[Cat.scala 33:92]
  wire  _decode_result_T_150 = &_decode_result_T_149; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_4_47 = io_in_instr[28]; // @[pla.scala 90:45]
  wire [4:0] _decode_result_T_151 = {decode_result_andMatrixInput_1_12,decode_result_andMatrixInput_2_18,
    decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_10,decode_result_andMatrixInput_4_47}; // @[Cat.scala 33:92]
  wire  _decode_result_T_152 = &_decode_result_T_151; // @[pla.scala 98:74]
  wire [6:0] decode_result_lo_lo_37 = {decode_result_andMatrixInput_22,decode_result_andMatrixInput_8,
    decode_result_andMatrixInput_9,decode_result_andMatrixInput_10,decode_result_andMatrixInput_4_47,
    decode_result_andMatrixInput_9_2,decode_result_andMatrixInput_13}; // @[Cat.scala 33:92]
  wire [13:0] decode_result_lo_60 = {decode_result_andMatrixInput_15,decode_result_andMatrixInput_16,
    decode_result_andMatrixInput_17,decode_result_andMatrixInput_18,decode_result_andMatrixInput_4_38,
    decode_result_andMatrixInput_20,decode_result_andMatrixInput_21,decode_result_lo_lo_37}; // @[Cat.scala 33:92]
  wire [6:0] decode_result_hi_lo_41 = {decode_result_andMatrixInput_6_16,decode_result_andMatrixInput_7_14,
    decode_result_andMatrixInput_8_10,decode_result_andMatrixInput_9_6,decode_result_andMatrixInput_6_3,
    decode_result_andMatrixInput_13_4,decode_result_andMatrixInput_14_2}; // @[Cat.scala 33:92]
  wire [28:0] _decode_result_T_153 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_2_18,decode_result_andMatrixInput_3_17,decode_result_andMatrixInput_5_17,
    decode_result_hi_lo_41,decode_result_lo_60}; // @[Cat.scala 33:92]
  wire  _decode_result_T_154 = &_decode_result_T_153; // @[pla.scala 98:74]
  wire [14:0] decode_result_lo_61 = {decode_result_andMatrixInput_14_2,decode_result_andMatrixInput_15,
    decode_result_andMatrixInput_16,decode_result_andMatrixInput_17,decode_result_andMatrixInput_18,
    decode_result_andMatrixInput_4_38,decode_result_andMatrixInput_20,decode_result_andMatrixInput_21,
    decode_result_lo_lo_37}; // @[Cat.scala 33:92]
  wire [30:0] _decode_result_T_155 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_2_18,decode_result_andMatrixInput_3_17,decode_result_andMatrixInput_5_17,
    decode_result_hi_lo_19,decode_result_lo_61}; // @[Cat.scala 33:92]
  wire  _decode_result_T_156 = &_decode_result_T_155; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_20_5 = io_in_instr[22]; // @[pla.scala 90:45]
  wire [6:0] decode_result_lo_lo_39 = {decode_result_andMatrixInput_22,decode_result_andMatrixInput_9,
    decode_result_andMatrixInput_10,decode_result_andMatrixInput_4_47,decode_result_andMatrixInput_12,
    decode_result_andMatrixInput_9_2,decode_result_andMatrixInput_13}; // @[Cat.scala 33:92]
  wire [13:0] decode_result_lo_62 = {decode_result_andMatrixInput_15,decode_result_andMatrixInput_16,
    decode_result_andMatrixInput_17,decode_result_andMatrixInput_20_2,decode_result_andMatrixInput_19,
    decode_result_andMatrixInput_20_5,decode_result_andMatrixInput_21,decode_result_lo_lo_39}; // @[Cat.scala 33:92]
  wire [28:0] _decode_result_T_157 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_2_18,decode_result_andMatrixInput_3_17,decode_result_andMatrixInput_5_17,
    decode_result_hi_lo_41,decode_result_lo_62}; // @[Cat.scala 33:92]
  wire  _decode_result_T_158 = &_decode_result_T_157; // @[pla.scala 98:74]
  wire [4:0] decode_result_lo_lo_40 = {decode_result_andMatrixInput_10,decode_result_andMatrixInput_4_47,
    decode_result_andMatrixInput_12,decode_result_andMatrixInput_9_2,decode_result_andMatrixInput_13}; // @[Cat.scala 33:92]
  wire [9:0] decode_result_lo_63 = {decode_result_andMatrixInput_8_10,decode_result_andMatrixInput_9_6,
    decode_result_andMatrixInput_6_3,decode_result_andMatrixInput_7_31,decode_result_andMatrixInput_9,
    decode_result_andMatrixInput_10,decode_result_andMatrixInput_4_47,decode_result_andMatrixInput_12,
    decode_result_andMatrixInput_9_2,decode_result_andMatrixInput_13}; // @[Cat.scala 33:92]
  wire [9:0] decode_result_hi_73 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_2_18,decode_result_andMatrixInput_3_17,decode_result_andMatrixInput_5_17,
    decode_result_andMatrixInput_6_16,decode_result_andMatrixInput_7_14}; // @[Cat.scala 33:92]
  wire [19:0] _decode_result_T_159 = {decode_result_hi_73,decode_result_lo_63}; // @[Cat.scala 33:92]
  wire  _decode_result_T_160 = &_decode_result_T_159; // @[pla.scala 98:74]
  wire [10:0] decode_result_lo_64 = {decode_result_andMatrixInput_9_6,decode_result_andMatrixInput_6,
    decode_result_andMatrixInput_7_1,decode_result_andMatrixInput_6_3,decode_result_andMatrixInput_7_31,
    decode_result_andMatrixInput_9,decode_result_lo_lo_40}; // @[Cat.scala 33:92]
  wire [4:0] decode_result_hi_lo_45 = {decode_result_andMatrixInput_3_17,decode_result_andMatrixInput_5_17,
    decode_result_andMatrixInput_6_16,decode_result_andMatrixInput_7_14,decode_result_andMatrixInput_8_10}; // @[Cat.scala 33:92]
  wire [21:0] _decode_result_T_161 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_2_18,decode_result_hi_lo_45,decode_result_lo_64}; // @[Cat.scala 33:92]
  wire  _decode_result_T_162 = &_decode_result_T_161; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_3_65 = io_in_instr[29]; // @[pla.scala 90:45]
  wire [4:0] _decode_result_T_163 = {decode_result_andMatrixInput_1_12,decode_result_andMatrixInput_2_18,
    decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_3_65,decode_result_andMatrixInput_13}; // @[Cat.scala 33:92]
  wire  _decode_result_T_164 = &_decode_result_T_163; // @[pla.scala 98:74]
  wire [4:0] _decode_result_T_165 = {decode_result_andMatrixInput_3_7,decode_result_andMatrixInput_3_17,
    decode_result_andMatrixInput_6,decode_result_andMatrixInput_7_1,decode_result_andMatrixInput_3_65}; // @[Cat.scala 33:92]
  wire  _decode_result_T_166 = &_decode_result_T_165; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_3_67 = io_in_instr[30]; // @[pla.scala 90:45]
  wire [3:0] _decode_result_T_167 = {decode_result_andMatrixInput_0,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_2_18,decode_result_andMatrixInput_3_67}; // @[Cat.scala 33:92]
  wire  _decode_result_T_168 = &_decode_result_T_167; // @[pla.scala 98:74]
  wire [4:0] _decode_result_T_169 = {decode_result_andMatrixInput_0,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_0_34,decode_result_andMatrixInput_7_1,decode_result_andMatrixInput_3_67}; // @[Cat.scala 33:92]
  wire  _decode_result_T_170 = &_decode_result_T_169; // @[pla.scala 98:74]
  wire [5:0] _decode_result_T_171 = {decode_result_andMatrixInput_1_12,decode_result_andMatrixInput_1_2,
    decode_result_andMatrixInput_1_42,decode_result_andMatrixInput_12,decode_result_andMatrixInput_3_67,
    decode_result_andMatrixInput_13}; // @[Cat.scala 33:92]
  wire  _decode_result_T_172 = &_decode_result_T_171; // @[pla.scala 98:74]
  wire [4:0] _decode_result_T_173 = {decode_result_andMatrixInput_1_12,decode_result_andMatrixInput_2_18,
    decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_3_65,decode_result_andMatrixInput_3_67}; // @[Cat.scala 33:92]
  wire  _decode_result_T_174 = &_decode_result_T_173; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_4_58 = io_in_instr[31]; // @[pla.scala 90:45]
  wire [4:0] _decode_result_T_175 = {decode_result_andMatrixInput_1_12,decode_result_andMatrixInput_2_18,
    decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_3_65,decode_result_andMatrixInput_4_58}; // @[Cat.scala 33:92]
  wire  _decode_result_T_176 = &_decode_result_T_175; // @[pla.scala 98:74]
  wire [4:0] _decode_result_T_177 = {decode_result_andMatrixInput_1_12,decode_result_andMatrixInput_2_18,
    decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_3_67,decode_result_andMatrixInput_4_58}; // @[Cat.scala 33:92]
  wire  _decode_result_T_178 = &_decode_result_T_177; // @[pla.scala 98:74]
  wire [5:0] _decode_result_orMatrixOutputs_T = {_decode_result_T_39,_decode_result_T_41,_decode_result_T_43,
    _decode_result_T_76,_decode_result_T_124,_decode_result_T_142}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_1 = |_decode_result_orMatrixOutputs_T; // @[pla.scala 114:39]
  wire [2:0] _decode_result_orMatrixOutputs_T_2 = {_decode_result_T_35,_decode_result_T_45,_decode_result_T_55}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_3 = |_decode_result_orMatrixOutputs_T_2; // @[pla.scala 114:39]
  wire [2:0] _decode_result_orMatrixOutputs_T_4 = {_decode_result_T_35,_decode_result_T_51,_decode_result_T_114}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_5 = |_decode_result_orMatrixOutputs_T_4; // @[pla.scala 114:39]
  wire [1:0] _decode_result_orMatrixOutputs_T_6 = {_decode_result_T_53,_decode_result_T_55}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_7 = |_decode_result_orMatrixOutputs_T_6; // @[pla.scala 114:39]
  wire [9:0] decode_result_orMatrixOutputs_lo_1 = {_decode_result_T_84,_decode_result_T_90,_decode_result_T_94,
    _decode_result_T_98,_decode_result_T_102,_decode_result_T_112,_decode_result_T_122,_decode_result_T_136,
    _decode_result_T_140,_decode_result_T_150}; // @[Cat.scala 33:92]
  wire [9:0] decode_result_orMatrixOutputs_hi_3 = {_decode_result_T_7,_decode_result_T_11,_decode_result_T_15,
    _decode_result_T_29,_decode_result_T_31,_decode_result_T_33,_decode_result_T_37,_decode_result_T_63,
    _decode_result_T_65,_decode_result_T_74}; // @[Cat.scala 33:92]
  wire [19:0] _decode_result_orMatrixOutputs_T_8 = {decode_result_orMatrixOutputs_hi_3,
    decode_result_orMatrixOutputs_lo_1}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_9 = |_decode_result_orMatrixOutputs_T_8; // @[pla.scala 114:39]
  wire [4:0] _decode_result_orMatrixOutputs_T_10 = {_decode_result_T_1,_decode_result_T_19,_decode_result_T_35,
    _decode_result_T_45,_decode_result_T_53}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_11 = |_decode_result_orMatrixOutputs_T_10; // @[pla.scala 114:39]
  wire [6:0] _decode_result_orMatrixOutputs_T_12 = {_decode_result_T_5,_decode_result_T_19,_decode_result_T_25,
    _decode_result_T_35,_decode_result_T_51,_decode_result_T_53,_decode_result_T_114}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_13 = |_decode_result_orMatrixOutputs_T_12; // @[pla.scala 114:39]
  wire [2:0] _decode_result_orMatrixOutputs_T_14 = {_decode_result_T_21,_decode_result_T_53,_decode_result_T_116}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_15 = |_decode_result_orMatrixOutputs_T_14; // @[pla.scala 114:39]
  wire [9:0] _decode_result_orMatrixOutputs_T_16 = {_decode_result_T_5,_decode_result_T_19,_decode_result_T_25,
    _decode_result_T_47,_decode_result_T_51,_decode_result_T_72,_decode_result_T_86,_decode_result_T_114,
    _decode_result_T_144,_decode_result_T_152}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_17 = |_decode_result_orMatrixOutputs_T_16; // @[pla.scala 114:39]
  wire [1:0] _decode_result_orMatrixOutputs_T_18 = {_decode_result_T_70,_decode_result_T_166}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_19 = |_decode_result_orMatrixOutputs_T_18; // @[pla.scala 114:39]
  wire [1:0] _decode_result_orMatrixOutputs_T_20 = {_decode_result_T_132,_decode_result_T_138}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_21 = |_decode_result_orMatrixOutputs_T_20; // @[pla.scala 114:39]
  wire [1:0] _decode_result_orMatrixOutputs_T_22 = {_decode_result_T_23,_decode_result_T_138}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_23 = |_decode_result_orMatrixOutputs_T_22; // @[pla.scala 114:39]
  wire  _decode_result_orMatrixOutputs_T_24 = |_decode_result_T_80; // @[pla.scala 114:39]
  wire  _decode_result_orMatrixOutputs_T_25 = |_decode_result_T_100; // @[pla.scala 114:39]
  wire  _decode_result_orMatrixOutputs_T_26 = |_decode_result_T_68; // @[pla.scala 114:39]
  wire [3:0] _decode_result_orMatrixOutputs_T_27 = {_decode_result_T_47,_decode_result_T_86,_decode_result_T_144,
    _decode_result_T_152}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_28 = |_decode_result_orMatrixOutputs_T_27; // @[pla.scala 114:39]
  wire [3:0] _decode_result_orMatrixOutputs_T_29 = {_decode_result_T_45,_decode_result_T_144,_decode_result_T_172,
    _decode_result_T_176}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_30 = |_decode_result_orMatrixOutputs_T_29; // @[pla.scala 114:39]
  wire [4:0] _decode_result_orMatrixOutputs_T_31 = {_decode_result_T_3,_decode_result_T_146,_decode_result_T_152,
    _decode_result_T_174,_decode_result_T_178}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_32 = |_decode_result_orMatrixOutputs_T_31; // @[pla.scala 114:39]
  wire [1:0] _decode_result_orMatrixOutputs_T_33 = {_decode_result_T_49,_decode_result_T_106}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_34 = |_decode_result_orMatrixOutputs_T_33; // @[pla.scala 114:39]
  wire [3:0] _decode_result_orMatrixOutputs_T_35 = {_decode_result_T_144,_decode_result_T_152,_decode_result_T_164,
    _decode_result_T_172}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_36 = |_decode_result_orMatrixOutputs_T_35; // @[pla.scala 114:39]
  wire  _decode_result_orMatrixOutputs_T_37 = |_decode_result_T_47; // @[pla.scala 114:39]
  wire [1:0] _decode_result_orMatrixOutputs_T_38 = {_decode_result_T_72,_decode_result_T_104}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_39 = |_decode_result_orMatrixOutputs_T_38; // @[pla.scala 114:39]
  wire  _decode_result_orMatrixOutputs_T_40 = |_decode_result_T_86; // @[pla.scala 114:39]
  wire  _decode_result_orMatrixOutputs_T_41 = |_decode_result_T_110; // @[pla.scala 114:39]
  wire [2:0] _decode_result_orMatrixOutputs_T_42 = {_decode_result_T_19,_decode_result_T_51,_decode_result_T_114}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_43 = |_decode_result_orMatrixOutputs_T_42; // @[pla.scala 114:39]
  wire [1:0] _decode_result_orMatrixOutputs_T_44 = {_decode_result_T_19,_decode_result_T_53}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_45 = |_decode_result_orMatrixOutputs_T_44; // @[pla.scala 114:39]
  wire [2:0] _decode_result_orMatrixOutputs_T_46 = {_decode_result_T_72,_decode_result_T_78,_decode_result_T_120}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_47 = |_decode_result_orMatrixOutputs_T_46; // @[pla.scala 114:39]
  wire [5:0] _decode_result_orMatrixOutputs_T_48 = {_decode_result_T_51,_decode_result_T_104,_decode_result_T_126,
    _decode_result_T_128,_decode_result_T_168,_decode_result_T_170}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_49 = |_decode_result_orMatrixOutputs_T_48; // @[pla.scala 114:39]
  wire [4:0] _decode_result_orMatrixOutputs_T_50 = {_decode_result_T_88,_decode_result_T_108,_decode_result_T_110,
    _decode_result_T_114,_decode_result_T_126}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_51 = |_decode_result_orMatrixOutputs_T_50; // @[pla.scala 114:39]
  wire [3:0] _decode_result_orMatrixOutputs_T_52 = {_decode_result_T_88,_decode_result_T_114,_decode_result_T_168,
    _decode_result_T_170}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_53 = |_decode_result_orMatrixOutputs_T_52; // @[pla.scala 114:39]
  wire [6:0] decode_result_orMatrixOutputs_lo_12 = {_decode_result_T_67,_decode_result_T_94,_decode_result_T_98,
    _decode_result_T_118,_decode_result_T_150,_decode_result_T_156,_decode_result_T_162}; // @[Cat.scala 33:92]
  wire [13:0] _decode_result_orMatrixOutputs_T_54 = {_decode_result_T_9,_decode_result_T_11,_decode_result_T_13,
    _decode_result_T_27,_decode_result_T_57,_decode_result_T_63,_decode_result_T_65,decode_result_orMatrixOutputs_lo_12}
    ; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_55 = |_decode_result_orMatrixOutputs_T_54; // @[pla.scala 114:39]
  wire [8:0] _decode_result_orMatrixOutputs_T_56 = {_decode_result_T_9,_decode_result_T_11,_decode_result_T_13,
    _decode_result_T_94,_decode_result_T_98,_decode_result_T_134,_decode_result_T_136,_decode_result_T_140,
    _decode_result_T_150}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_57 = |_decode_result_orMatrixOutputs_T_56; // @[pla.scala 114:39]
  wire [5:0] _decode_result_orMatrixOutputs_T_58 = {_decode_result_T_27,_decode_result_T_67,_decode_result_T_84,
    _decode_result_T_102,_decode_result_T_156,_decode_result_T_162}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_59 = |_decode_result_orMatrixOutputs_T_58; // @[pla.scala 114:39]
  wire  _decode_result_orMatrixOutputs_T_60 = |_decode_result_T_67; // @[pla.scala 114:39]
  wire  _decode_result_orMatrixOutputs_T_61 = |_decode_result_T_130; // @[pla.scala 114:39]
  wire [5:0] decode_result_orMatrixOutputs_lo_lo_4 = {_decode_result_T_122,_decode_result_T_142,_decode_result_T_148,
    _decode_result_T_154,_decode_result_T_158,_decode_result_T_160}; // @[Cat.scala 33:92]
  wire [12:0] decode_result_orMatrixOutputs_lo_15 = {_decode_result_T_82,_decode_result_T_90,_decode_result_T_92,
    _decode_result_T_96,_decode_result_T_102,_decode_result_T_112,_decode_result_T_118,
    decode_result_orMatrixOutputs_lo_lo_4}; // @[Cat.scala 33:92]
  wire [6:0] decode_result_orMatrixOutputs_hi_lo_5 = {_decode_result_T_39,_decode_result_T_41,_decode_result_T_43,
    _decode_result_T_59,_decode_result_T_61,_decode_result_T_65,_decode_result_T_76}; // @[Cat.scala 33:92]
  wire [26:0] _decode_result_orMatrixOutputs_T_62 = {_decode_result_T_7,_decode_result_T_11,_decode_result_T_13,
    _decode_result_T_17,_decode_result_T_27,_decode_result_T_33,_decode_result_T_37,
    decode_result_orMatrixOutputs_hi_lo_5,decode_result_orMatrixOutputs_lo_15}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_63 = |_decode_result_orMatrixOutputs_T_62; // @[pla.scala 114:39]
  wire [6:0] decode_result_orMatrixOutputs_lo_lo_5 = {_decode_result_T_122,_decode_result_T_136,_decode_result_T_140,
    _decode_result_T_150,_decode_result_T_156,_decode_result_T_158,_decode_result_T_162}; // @[Cat.scala 33:92]
  wire [13:0] decode_result_orMatrixOutputs_lo_16 = {_decode_result_T_84,_decode_result_T_90,_decode_result_T_94,
    _decode_result_T_98,_decode_result_T_102,_decode_result_T_112,_decode_result_T_118,
    decode_result_orMatrixOutputs_lo_lo_5}; // @[Cat.scala 33:92]
  wire [6:0] decode_result_orMatrixOutputs_hi_lo_6 = {_decode_result_T_37,_decode_result_T_57,_decode_result_T_61,
    _decode_result_T_63,_decode_result_T_65,_decode_result_T_67,_decode_result_T_74}; // @[Cat.scala 33:92]
  wire [27:0] _decode_result_orMatrixOutputs_T_64 = {_decode_result_T_7,_decode_result_T_11,_decode_result_T_13,
    _decode_result_T_27,_decode_result_T_29,_decode_result_T_31,_decode_result_T_33,
    decode_result_orMatrixOutputs_hi_lo_6,decode_result_orMatrixOutputs_lo_16}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_65 = |_decode_result_orMatrixOutputs_T_64; // @[pla.scala 114:39]
  wire [9:0] decode_result_orMatrixOutputs_lo_hi_10 = {_decode_result_orMatrixOutputs_T_34,
    _decode_result_orMatrixOutputs_T_32,_decode_result_orMatrixOutputs_T_30,_decode_result_orMatrixOutputs_T_28,
    _decode_result_orMatrixOutputs_T_26,_decode_result_orMatrixOutputs_T_25,_decode_result_orMatrixOutputs_T_24,
    _decode_result_orMatrixOutputs_T_23,_decode_result_orMatrixOutputs_T_21,_decode_result_orMatrixOutputs_T_19}; // @[Cat.scala 33:92]
  wire [18:0] decode_result_orMatrixOutputs_lo_17 = {decode_result_orMatrixOutputs_lo_hi_10,
    _decode_result_orMatrixOutputs_T_17,_decode_result_orMatrixOutputs_T_15,_decode_result_orMatrixOutputs_T_13,
    _decode_result_orMatrixOutputs_T_11,_decode_result_orMatrixOutputs_T_9,_decode_result_orMatrixOutputs_T_7,
    _decode_result_orMatrixOutputs_T_5,_decode_result_orMatrixOutputs_T_3,_decode_result_orMatrixOutputs_T_1}; // @[Cat.scala 33:92]
  wire [9:0] decode_result_orMatrixOutputs_hi_hi_13 = {_decode_result_orMatrixOutputs_T_65,
    _decode_result_orMatrixOutputs_T_63,_decode_result_orMatrixOutputs_T_61,_decode_result_orMatrixOutputs_T_60,
    _decode_result_orMatrixOutputs_T_59,_decode_result_orMatrixOutputs_T_57,_decode_result_orMatrixOutputs_T_55,
    _decode_result_orMatrixOutputs_T_53,_decode_result_orMatrixOutputs_T_51,_decode_result_orMatrixOutputs_T_49}; // @[Cat.scala 33:92]
  wire [18:0] decode_result_orMatrixOutputs_hi_22 = {decode_result_orMatrixOutputs_hi_hi_13,
    _decode_result_orMatrixOutputs_T_47,_decode_result_orMatrixOutputs_T_45,_decode_result_orMatrixOutputs_T_43,1'h0,
    _decode_result_orMatrixOutputs_T_41,_decode_result_orMatrixOutputs_T_40,_decode_result_orMatrixOutputs_T_39,
    _decode_result_orMatrixOutputs_T_37,_decode_result_orMatrixOutputs_T_36}; // @[Cat.scala 33:92]
  wire [37:0] decode_result_orMatrixOutputs = {decode_result_orMatrixOutputs_hi_22,decode_result_orMatrixOutputs_lo_17}; // @[Cat.scala 33:92]
  wire  _decode_result_invMatrixOutputs_T_1 = ~decode_result_orMatrixOutputs[0]; // @[pla.scala 123:40]
  wire  _decode_result_invMatrixOutputs_T_38 = ~decode_result_orMatrixOutputs[36]; // @[pla.scala 123:40]
  wire [9:0] decode_result_invMatrixOutputs_lo_hi = {decode_result_orMatrixOutputs[18],decode_result_orMatrixOutputs[17]
    ,decode_result_orMatrixOutputs[16],decode_result_orMatrixOutputs[15],decode_result_orMatrixOutputs[14],
    decode_result_orMatrixOutputs[13],decode_result_orMatrixOutputs[12],decode_result_orMatrixOutputs[11],
    decode_result_orMatrixOutputs[10],decode_result_orMatrixOutputs[9]}; // @[Cat.scala 33:92]
  wire [18:0] decode_result_invMatrixOutputs_lo = {decode_result_invMatrixOutputs_lo_hi,decode_result_orMatrixOutputs[8]
    ,decode_result_orMatrixOutputs[7],decode_result_orMatrixOutputs[6],decode_result_orMatrixOutputs[5],
    decode_result_orMatrixOutputs[4],decode_result_orMatrixOutputs[3],decode_result_orMatrixOutputs[2],
    decode_result_orMatrixOutputs[1],_decode_result_invMatrixOutputs_T_1}; // @[Cat.scala 33:92]
  wire [9:0] decode_result_invMatrixOutputs_hi_hi = {decode_result_orMatrixOutputs[37],
    _decode_result_invMatrixOutputs_T_38,decode_result_orMatrixOutputs[35],decode_result_orMatrixOutputs[34],
    decode_result_orMatrixOutputs[33],decode_result_orMatrixOutputs[32],decode_result_orMatrixOutputs[31],
    decode_result_orMatrixOutputs[30],decode_result_orMatrixOutputs[29],decode_result_orMatrixOutputs[28]}; // @[Cat.scala 33:92]
  wire [18:0] decode_result_invMatrixOutputs_hi = {decode_result_invMatrixOutputs_hi_hi,decode_result_orMatrixOutputs[27
    ],decode_result_orMatrixOutputs[26],decode_result_orMatrixOutputs[25],decode_result_orMatrixOutputs[24],
    decode_result_orMatrixOutputs[23],decode_result_orMatrixOutputs[22],decode_result_orMatrixOutputs[21],
    decode_result_orMatrixOutputs[20],decode_result_orMatrixOutputs[19]}; // @[Cat.scala 33:92]
  wire [37:0] decode_result_invMatrixOutputs = {decode_result_invMatrixOutputs_hi,decode_result_invMatrixOutputs_lo}; // @[Cat.scala 33:92]
  wire  uop_dw = decode_result_invMatrixOutputs[0]; // @[MicroOp.scala 56:20]
  wire [2:0] imm_type = decode_result_invMatrixOutputs[3:1]; // @[MicroOp.scala 58:20]
  wire  uop_rd_wen = decode_result_invMatrixOutputs[4]; // @[MicroOp.scala 56:20]
  wire [1:0] uop_rs2_src = decode_result_invMatrixOutputs[6:5]; // @[MicroOp.scala 58:20]
  wire [1:0] uop_rs1_src = decode_result_invMatrixOutputs[8:7]; // @[MicroOp.scala 58:20]
  wire [2:0] uop_sys_op = decode_result_invMatrixOutputs[11:9]; // @[MicroOp.scala 58:20]
  wire [1:0] uop_csr_op = decode_result_invMatrixOutputs[13:12]; // @[MicroOp.scala 58:20]
  wire [1:0] uop_mem_len = decode_result_invMatrixOutputs[15:14]; // @[MicroOp.scala 58:20]
  wire [4:0] uop_lsu_op = decode_result_invMatrixOutputs[20:16]; // @[MicroOp.scala 58:20]
  wire [3:0] uop_mdu_op = decode_result_invMatrixOutputs[24:21]; // @[MicroOp.scala 58:20]
  wire [1:0] uop_jmp_op = decode_result_invMatrixOutputs[26:25]; // @[MicroOp.scala 58:20]
  wire [3:0] uop_alu_op = decode_result_invMatrixOutputs[30:27]; // @[MicroOp.scala 58:20]
  wire [2:0] uop_fu = decode_result_invMatrixOutputs[33:31]; // @[MicroOp.scala 58:20]
  wire [20:0] _imm_i_T_2 = decode_result_andMatrixInput_4_58 ? 21'h1fffff : 21'h0; // @[Bitwise.scala 77:12]
  wire [31:0] imm_i = {_imm_i_T_2,io_in_instr[30:20]}; // @[Cat.scala 33:92]
  wire [31:0] imm_s = {_imm_i_T_2,io_in_instr[30:25],uop_rd_index}; // @[Cat.scala 33:92]
  wire [19:0] _imm_b_T_2 = decode_result_andMatrixInput_4_58 ? 20'hfffff : 20'h0; // @[Bitwise.scala 77:12]
  wire [31:0] imm_b = {_imm_b_T_2,io_in_instr[7],io_in_instr[30:25],io_in_instr[11:8],1'h0}; // @[Cat.scala 33:92]
  wire [31:0] imm_u = {io_in_instr[31:12],12'h0}; // @[Cat.scala 33:92]
  wire [11:0] _imm_j_T_2 = decode_result_andMatrixInput_4_58 ? 12'hfff : 12'h0; // @[Bitwise.scala 77:12]
  wire [31:0] imm_j = {_imm_j_T_2,io_in_instr[19:12],decode_result_andMatrixInput_20_2,io_in_instr[30:21],1'h0}; // @[Cat.scala 33:92]
  wire [31:0] imm_csr = {27'h0,uop_rs1_index}; // @[Cat.scala 33:92]
  wire [31:0] _uop_imm_T_1 = 3'h0 == imm_type ? imm_i : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] _uop_imm_T_3 = 3'h1 == imm_type ? imm_s : _uop_imm_T_1; // @[Mux.scala 81:58]
  wire [31:0] _uop_imm_T_5 = 3'h2 == imm_type ? imm_b : _uop_imm_T_3; // @[Mux.scala 81:58]
  wire [31:0] _uop_imm_T_7 = 3'h3 == imm_type ? imm_u : _uop_imm_T_5; // @[Mux.scala 81:58]
  wire [31:0] _uop_imm_T_9 = 3'h4 == imm_type ? imm_j : _uop_imm_T_7; // @[Mux.scala 81:58]
  wire [31:0] uop_imm = 3'h5 == imm_type ? imm_csr : _uop_imm_T_9; // @[Mux.scala 81:58]
  wire [2:0] _GEN_0 = io_in_access_fault ? 3'h2 : decode_result_invMatrixOutputs[36:34]; // @[Decode.scala 30:36 31:17 MicroOp.scala 58:15]
  wire  _GEN_1 = io_in_access_fault ? 1'h0 : decode_result_invMatrixOutputs[37]; // @[Decode.scala 30:36 32:17 MicroOp.scala 56:15]
  wire [2:0] _GEN_2 = io_in_page_fault ? 3'h3 : _GEN_0; // @[Decode.scala 27:28 28:17]
  wire  _GEN_3 = io_in_page_fault ? 1'h0 : _GEN_1; // @[Decode.scala 27:28 29:17]
  wire [2:0] uop_exc = io_in_valid ? _GEN_2 : decode_result_invMatrixOutputs[36:34]; // @[Decode.scala 26:21 MicroOp.scala 58:15]
  wire  uop_valid = io_in_valid ? _GEN_3 : decode_result_invMatrixOutputs[37]; // @[Decode.scala 26:21 MicroOp.scala 56:15]
  assign io_out_valid = io_in_valid & uop_valid; // @[Decode.scala 36:16]
  assign io_out_exc = io_in_valid ? uop_exc : 3'h0; // @[Decode.scala 36:16]
  assign io_out_pc = io_in_valid ? io_in_pc : 64'h0; // @[Decode.scala 36:16]
  assign io_out_npc = io_in_valid ? uop_npc : 64'h0; // @[Decode.scala 36:16]
  assign io_out_instr = io_in_valid ? io_in_instr : 32'h0; // @[Decode.scala 36:16]
  assign io_out_fu = io_in_valid ? uop_fu : 3'h0; // @[Decode.scala 36:16]
  assign io_out_alu_op = io_in_valid ? uop_alu_op : 4'h0; // @[Decode.scala 36:16]
  assign io_out_jmp_op = io_in_valid ? uop_jmp_op : 2'h0; // @[Decode.scala 36:16]
  assign io_out_mdu_op = io_in_valid ? uop_mdu_op : 4'h0; // @[Decode.scala 36:16]
  assign io_out_lsu_op = io_in_valid ? uop_lsu_op : 5'h0; // @[Decode.scala 36:16]
  assign io_out_mem_len = io_in_valid ? uop_mem_len : 2'h0; // @[Decode.scala 36:16]
  assign io_out_csr_op = io_in_valid ? uop_csr_op : 2'h0; // @[Decode.scala 36:16]
  assign io_out_sys_op = io_in_valid ? uop_sys_op : 3'h0; // @[Decode.scala 36:16]
  assign io_out_rs1_src = io_in_valid ? uop_rs1_src : 2'h0; // @[Decode.scala 36:16]
  assign io_out_rs2_src = io_in_valid ? uop_rs2_src : 2'h0; // @[Decode.scala 36:16]
  assign io_out_rs1_index = io_in_valid ? uop_rs1_index : 5'h0; // @[Decode.scala 36:16]
  assign io_out_rs2_index = io_in_valid ? uop_rs2_index : 5'h0; // @[Decode.scala 36:16]
  assign io_out_rd_index = io_in_valid ? uop_rd_index : 5'h0; // @[Decode.scala 36:16]
  assign io_out_rd_wen = io_in_valid & uop_rd_wen; // @[Decode.scala 36:16]
  assign io_out_imm = io_in_valid ? uop_imm : 32'h0; // @[Decode.scala 36:16]
  assign io_out_dw = io_in_valid & uop_dw; // @[Decode.scala 36:16]
endmodule
module RegFile(
  input         clock,
  input         reset,
  input  [4:0]  io_rs1_index,
  input  [4:0]  io_rs2_index,
  output [63:0] io_rs1_data,
  output [63:0] io_rs2_data,
  input  [4:0]  io_rd_index,
  input  [63:0] io_rd_data,
  input         io_rd_wen
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] rf_0; // @[RegFile.scala 21:19]
  reg [63:0] rf_1; // @[RegFile.scala 21:19]
  reg [63:0] rf_2; // @[RegFile.scala 21:19]
  reg [63:0] rf_3; // @[RegFile.scala 21:19]
  reg [63:0] rf_4; // @[RegFile.scala 21:19]
  reg [63:0] rf_5; // @[RegFile.scala 21:19]
  reg [63:0] rf_6; // @[RegFile.scala 21:19]
  reg [63:0] rf_7; // @[RegFile.scala 21:19]
  reg [63:0] rf_8; // @[RegFile.scala 21:19]
  reg [63:0] rf_9; // @[RegFile.scala 21:19]
  reg [63:0] rf_10; // @[RegFile.scala 21:19]
  reg [63:0] rf_11; // @[RegFile.scala 21:19]
  reg [63:0] rf_12; // @[RegFile.scala 21:19]
  reg [63:0] rf_13; // @[RegFile.scala 21:19]
  reg [63:0] rf_14; // @[RegFile.scala 21:19]
  reg [63:0] rf_15; // @[RegFile.scala 21:19]
  reg [63:0] rf_16; // @[RegFile.scala 21:19]
  reg [63:0] rf_17; // @[RegFile.scala 21:19]
  reg [63:0] rf_18; // @[RegFile.scala 21:19]
  reg [63:0] rf_19; // @[RegFile.scala 21:19]
  reg [63:0] rf_20; // @[RegFile.scala 21:19]
  reg [63:0] rf_21; // @[RegFile.scala 21:19]
  reg [63:0] rf_22; // @[RegFile.scala 21:19]
  reg [63:0] rf_23; // @[RegFile.scala 21:19]
  reg [63:0] rf_24; // @[RegFile.scala 21:19]
  reg [63:0] rf_25; // @[RegFile.scala 21:19]
  reg [63:0] rf_26; // @[RegFile.scala 21:19]
  reg [63:0] rf_27; // @[RegFile.scala 21:19]
  reg [63:0] rf_28; // @[RegFile.scala 21:19]
  reg [63:0] rf_29; // @[RegFile.scala 21:19]
  reg [63:0] rf_30; // @[RegFile.scala 21:19]
  wire  _T_1 = io_rd_wen & io_rd_index != 5'h0; // @[RegFile.scala 23:18]
  wire [4:0] _T_2 = ~io_rd_index; // @[RegFile.scala 18:28]
  wire [4:0] _io_rs1_data_T_1 = ~io_rs1_index; // @[RegFile.scala 18:28]
  wire [63:0] _GEN_63 = 5'h1 == _io_rs1_data_T_1 ? rf_1 : rf_0; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_64 = 5'h2 == _io_rs1_data_T_1 ? rf_2 : _GEN_63; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_65 = 5'h3 == _io_rs1_data_T_1 ? rf_3 : _GEN_64; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_66 = 5'h4 == _io_rs1_data_T_1 ? rf_4 : _GEN_65; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_67 = 5'h5 == _io_rs1_data_T_1 ? rf_5 : _GEN_66; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_68 = 5'h6 == _io_rs1_data_T_1 ? rf_6 : _GEN_67; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_69 = 5'h7 == _io_rs1_data_T_1 ? rf_7 : _GEN_68; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_70 = 5'h8 == _io_rs1_data_T_1 ? rf_8 : _GEN_69; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_71 = 5'h9 == _io_rs1_data_T_1 ? rf_9 : _GEN_70; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_72 = 5'ha == _io_rs1_data_T_1 ? rf_10 : _GEN_71; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_73 = 5'hb == _io_rs1_data_T_1 ? rf_11 : _GEN_72; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_74 = 5'hc == _io_rs1_data_T_1 ? rf_12 : _GEN_73; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_75 = 5'hd == _io_rs1_data_T_1 ? rf_13 : _GEN_74; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_76 = 5'he == _io_rs1_data_T_1 ? rf_14 : _GEN_75; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_77 = 5'hf == _io_rs1_data_T_1 ? rf_15 : _GEN_76; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_78 = 5'h10 == _io_rs1_data_T_1 ? rf_16 : _GEN_77; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_79 = 5'h11 == _io_rs1_data_T_1 ? rf_17 : _GEN_78; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_80 = 5'h12 == _io_rs1_data_T_1 ? rf_18 : _GEN_79; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_81 = 5'h13 == _io_rs1_data_T_1 ? rf_19 : _GEN_80; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_82 = 5'h14 == _io_rs1_data_T_1 ? rf_20 : _GEN_81; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_83 = 5'h15 == _io_rs1_data_T_1 ? rf_21 : _GEN_82; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_84 = 5'h16 == _io_rs1_data_T_1 ? rf_22 : _GEN_83; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_85 = 5'h17 == _io_rs1_data_T_1 ? rf_23 : _GEN_84; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_86 = 5'h18 == _io_rs1_data_T_1 ? rf_24 : _GEN_85; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_87 = 5'h19 == _io_rs1_data_T_1 ? rf_25 : _GEN_86; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_88 = 5'h1a == _io_rs1_data_T_1 ? rf_26 : _GEN_87; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_89 = 5'h1b == _io_rs1_data_T_1 ? rf_27 : _GEN_88; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_90 = 5'h1c == _io_rs1_data_T_1 ? rf_28 : _GEN_89; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_91 = 5'h1d == _io_rs1_data_T_1 ? rf_29 : _GEN_90; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_92 = 5'h1e == _io_rs1_data_T_1 ? rf_30 : _GEN_91; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _io_rs1_data_T_2 = io_rs1_index != 5'h0 ? _GEN_92 : 64'h0; // @[RegFile.scala 27:21]
  wire [4:0] _io_rs2_data_T_1 = ~io_rs2_index; // @[RegFile.scala 18:28]
  wire [63:0] _GEN_94 = 5'h1 == _io_rs2_data_T_1 ? rf_1 : rf_0; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_95 = 5'h2 == _io_rs2_data_T_1 ? rf_2 : _GEN_94; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_96 = 5'h3 == _io_rs2_data_T_1 ? rf_3 : _GEN_95; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_97 = 5'h4 == _io_rs2_data_T_1 ? rf_4 : _GEN_96; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_98 = 5'h5 == _io_rs2_data_T_1 ? rf_5 : _GEN_97; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_99 = 5'h6 == _io_rs2_data_T_1 ? rf_6 : _GEN_98; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_100 = 5'h7 == _io_rs2_data_T_1 ? rf_7 : _GEN_99; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_101 = 5'h8 == _io_rs2_data_T_1 ? rf_8 : _GEN_100; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_102 = 5'h9 == _io_rs2_data_T_1 ? rf_9 : _GEN_101; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_103 = 5'ha == _io_rs2_data_T_1 ? rf_10 : _GEN_102; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_104 = 5'hb == _io_rs2_data_T_1 ? rf_11 : _GEN_103; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_105 = 5'hc == _io_rs2_data_T_1 ? rf_12 : _GEN_104; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_106 = 5'hd == _io_rs2_data_T_1 ? rf_13 : _GEN_105; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_107 = 5'he == _io_rs2_data_T_1 ? rf_14 : _GEN_106; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_108 = 5'hf == _io_rs2_data_T_1 ? rf_15 : _GEN_107; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_109 = 5'h10 == _io_rs2_data_T_1 ? rf_16 : _GEN_108; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_110 = 5'h11 == _io_rs2_data_T_1 ? rf_17 : _GEN_109; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_111 = 5'h12 == _io_rs2_data_T_1 ? rf_18 : _GEN_110; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_112 = 5'h13 == _io_rs2_data_T_1 ? rf_19 : _GEN_111; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_113 = 5'h14 == _io_rs2_data_T_1 ? rf_20 : _GEN_112; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_114 = 5'h15 == _io_rs2_data_T_1 ? rf_21 : _GEN_113; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_115 = 5'h16 == _io_rs2_data_T_1 ? rf_22 : _GEN_114; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_116 = 5'h17 == _io_rs2_data_T_1 ? rf_23 : _GEN_115; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_117 = 5'h18 == _io_rs2_data_T_1 ? rf_24 : _GEN_116; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_118 = 5'h19 == _io_rs2_data_T_1 ? rf_25 : _GEN_117; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_119 = 5'h1a == _io_rs2_data_T_1 ? rf_26 : _GEN_118; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_120 = 5'h1b == _io_rs2_data_T_1 ? rf_27 : _GEN_119; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_121 = 5'h1c == _io_rs2_data_T_1 ? rf_28 : _GEN_120; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_122 = 5'h1d == _io_rs2_data_T_1 ? rf_29 : _GEN_121; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_123 = 5'h1e == _io_rs2_data_T_1 ? rf_30 : _GEN_122; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _io_rs2_data_T_2 = io_rs2_index != 5'h0 ? _GEN_123 : 64'h0; // @[RegFile.scala 28:21]
  wire [63:0] _GEN_124 = io_rd_index == io_rs1_index ? io_rd_data : _io_rs1_data_T_2; // @[RegFile.scala 27:15 32:40 33:19]
  wire [63:0] _GEN_125 = io_rd_index == io_rs2_index ? io_rd_data : _io_rs2_data_T_2; // @[RegFile.scala 28:15 35:40 36:19]
  assign io_rs1_data = _T_1 ? _GEN_124 : _io_rs1_data_T_2; // @[RegFile.scala 27:15 31:44]
  assign io_rs2_data = _T_1 ? _GEN_125 : _io_rs2_data_T_2; // @[RegFile.scala 28:15 31:44]
  always @(posedge clock) begin
    if (reset) begin // @[RegFile.scala 21:19]
      rf_0 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h0 == _T_2) begin // @[RegFile.scala 24:25]
        rf_0 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_1 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h1 == _T_2) begin // @[RegFile.scala 24:25]
        rf_1 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_2 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h2 == _T_2) begin // @[RegFile.scala 24:25]
        rf_2 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_3 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h3 == _T_2) begin // @[RegFile.scala 24:25]
        rf_3 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_4 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h4 == _T_2) begin // @[RegFile.scala 24:25]
        rf_4 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_5 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h5 == _T_2) begin // @[RegFile.scala 24:25]
        rf_5 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_6 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h6 == _T_2) begin // @[RegFile.scala 24:25]
        rf_6 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_7 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h7 == _T_2) begin // @[RegFile.scala 24:25]
        rf_7 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_8 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h8 == _T_2) begin // @[RegFile.scala 24:25]
        rf_8 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_9 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h9 == _T_2) begin // @[RegFile.scala 24:25]
        rf_9 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_10 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'ha == _T_2) begin // @[RegFile.scala 24:25]
        rf_10 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_11 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'hb == _T_2) begin // @[RegFile.scala 24:25]
        rf_11 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_12 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'hc == _T_2) begin // @[RegFile.scala 24:25]
        rf_12 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_13 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'hd == _T_2) begin // @[RegFile.scala 24:25]
        rf_13 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_14 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'he == _T_2) begin // @[RegFile.scala 24:25]
        rf_14 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_15 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'hf == _T_2) begin // @[RegFile.scala 24:25]
        rf_15 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_16 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h10 == _T_2) begin // @[RegFile.scala 24:25]
        rf_16 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_17 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h11 == _T_2) begin // @[RegFile.scala 24:25]
        rf_17 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_18 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h12 == _T_2) begin // @[RegFile.scala 24:25]
        rf_18 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_19 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h13 == _T_2) begin // @[RegFile.scala 24:25]
        rf_19 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_20 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h14 == _T_2) begin // @[RegFile.scala 24:25]
        rf_20 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_21 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h15 == _T_2) begin // @[RegFile.scala 24:25]
        rf_21 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_22 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h16 == _T_2) begin // @[RegFile.scala 24:25]
        rf_22 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_23 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h17 == _T_2) begin // @[RegFile.scala 24:25]
        rf_23 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_24 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h18 == _T_2) begin // @[RegFile.scala 24:25]
        rf_24 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_25 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h19 == _T_2) begin // @[RegFile.scala 24:25]
        rf_25 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_26 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h1a == _T_2) begin // @[RegFile.scala 24:25]
        rf_26 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_27 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h1b == _T_2) begin // @[RegFile.scala 24:25]
        rf_27 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_28 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h1c == _T_2) begin // @[RegFile.scala 24:25]
        rf_28 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_29 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h1d == _T_2) begin // @[RegFile.scala 24:25]
        rf_29 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_30 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h1e == _T_2) begin // @[RegFile.scala 24:25]
        rf_30 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  rf_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  rf_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  rf_2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  rf_3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  rf_4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  rf_5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  rf_6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  rf_7 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  rf_8 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  rf_9 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  rf_10 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  rf_11 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  rf_12 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  rf_13 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  rf_14 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  rf_15 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  rf_16 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  rf_17 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  rf_18 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  rf_19 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  rf_20 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  rf_21 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  rf_22 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  rf_23 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  rf_24 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  rf_25 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  rf_26 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  rf_27 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  rf_28 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  rf_29 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  rf_30 = _RAND_30[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PipelineReg(
  input         clock,
  input         reset,
  input         io_in_uop_valid,
  input  [2:0]  io_in_uop_exc,
  input  [63:0] io_in_uop_pc,
  input  [63:0] io_in_uop_npc,
  input  [31:0] io_in_uop_instr,
  input  [2:0]  io_in_uop_fu,
  input  [3:0]  io_in_uop_alu_op,
  input  [1:0]  io_in_uop_jmp_op,
  input  [3:0]  io_in_uop_mdu_op,
  input  [4:0]  io_in_uop_lsu_op,
  input  [1:0]  io_in_uop_mem_len,
  input  [1:0]  io_in_uop_csr_op,
  input  [2:0]  io_in_uop_sys_op,
  input  [4:0]  io_in_uop_rd_index,
  input         io_in_uop_rd_wen,
  input  [31:0] io_in_uop_imm,
  input         io_in_uop_dw,
  input  [63:0] io_in_rs1_data,
  input  [63:0] io_in_rs2_data,
  input  [63:0] io_in_rs2_data_from_rf,
  input  [63:0] io_in_bp_npc,
  output        io_out_uop_valid,
  output [2:0]  io_out_uop_exc,
  output [63:0] io_out_uop_pc,
  output [63:0] io_out_uop_npc,
  output [31:0] io_out_uop_instr,
  output [2:0]  io_out_uop_fu,
  output [3:0]  io_out_uop_alu_op,
  output [1:0]  io_out_uop_jmp_op,
  output [3:0]  io_out_uop_mdu_op,
  output [4:0]  io_out_uop_lsu_op,
  output [1:0]  io_out_uop_mem_len,
  output [1:0]  io_out_uop_csr_op,
  output [2:0]  io_out_uop_sys_op,
  output [4:0]  io_out_uop_rd_index,
  output        io_out_uop_rd_wen,
  output [31:0] io_out_uop_imm,
  output        io_out_uop_dw,
  output [63:0] io_out_rs1_data,
  output [63:0] io_out_rs2_data,
  output [63:0] io_out_rs2_data_from_rf,
  output [63:0] io_out_bp_npc,
  input         io_en,
  input         io_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
`endif // RANDOMIZE_REG_INIT
  reg  reg_uop_valid; // @[Reg.scala 35:20]
  reg [2:0] reg_uop_exc; // @[Reg.scala 35:20]
  reg [63:0] reg_uop_pc; // @[Reg.scala 35:20]
  reg [63:0] reg_uop_npc; // @[Reg.scala 35:20]
  reg [31:0] reg_uop_instr; // @[Reg.scala 35:20]
  reg [2:0] reg_uop_fu; // @[Reg.scala 35:20]
  reg [3:0] reg_uop_alu_op; // @[Reg.scala 35:20]
  reg [1:0] reg_uop_jmp_op; // @[Reg.scala 35:20]
  reg [3:0] reg_uop_mdu_op; // @[Reg.scala 35:20]
  reg [4:0] reg_uop_lsu_op; // @[Reg.scala 35:20]
  reg [1:0] reg_uop_mem_len; // @[Reg.scala 35:20]
  reg [1:0] reg_uop_csr_op; // @[Reg.scala 35:20]
  reg [2:0] reg_uop_sys_op; // @[Reg.scala 35:20]
  reg [4:0] reg_uop_rd_index; // @[Reg.scala 35:20]
  reg  reg_uop_rd_wen; // @[Reg.scala 35:20]
  reg [31:0] reg_uop_imm; // @[Reg.scala 35:20]
  reg  reg_uop_dw; // @[Reg.scala 35:20]
  reg [63:0] reg_rs1_data; // @[Reg.scala 35:20]
  reg [63:0] reg_rs2_data; // @[Reg.scala 35:20]
  reg [63:0] reg_rs2_data_from_rf; // @[Reg.scala 35:20]
  reg [63:0] reg_bp_npc; // @[Reg.scala 35:20]
  assign io_out_uop_valid = reg_uop_valid; // @[DataType.scala 41:10]
  assign io_out_uop_exc = reg_uop_exc; // @[DataType.scala 41:10]
  assign io_out_uop_pc = reg_uop_pc; // @[DataType.scala 41:10]
  assign io_out_uop_npc = reg_uop_npc; // @[DataType.scala 41:10]
  assign io_out_uop_instr = reg_uop_instr; // @[DataType.scala 41:10]
  assign io_out_uop_fu = reg_uop_fu; // @[DataType.scala 41:10]
  assign io_out_uop_alu_op = reg_uop_alu_op; // @[DataType.scala 41:10]
  assign io_out_uop_jmp_op = reg_uop_jmp_op; // @[DataType.scala 41:10]
  assign io_out_uop_mdu_op = reg_uop_mdu_op; // @[DataType.scala 41:10]
  assign io_out_uop_lsu_op = reg_uop_lsu_op; // @[DataType.scala 41:10]
  assign io_out_uop_mem_len = reg_uop_mem_len; // @[DataType.scala 41:10]
  assign io_out_uop_csr_op = reg_uop_csr_op; // @[DataType.scala 41:10]
  assign io_out_uop_sys_op = reg_uop_sys_op; // @[DataType.scala 41:10]
  assign io_out_uop_rd_index = reg_uop_rd_index; // @[DataType.scala 41:10]
  assign io_out_uop_rd_wen = reg_uop_rd_wen; // @[DataType.scala 41:10]
  assign io_out_uop_imm = reg_uop_imm; // @[DataType.scala 41:10]
  assign io_out_uop_dw = reg_uop_dw; // @[DataType.scala 41:10]
  assign io_out_rs1_data = reg_rs1_data; // @[DataType.scala 41:10]
  assign io_out_rs2_data = reg_rs2_data; // @[DataType.scala 41:10]
  assign io_out_rs2_data_from_rf = reg_rs2_data_from_rf; // @[DataType.scala 41:10]
  assign io_out_bp_npc = reg_bp_npc; // @[DataType.scala 41:10]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 35:20]
      reg_uop_valid <= 1'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_flush) begin // @[DataType.scala 40:26]
        reg_uop_valid <= 1'h0;
      end else begin
        reg_uop_valid <= io_in_uop_valid;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      reg_uop_exc <= 3'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_flush) begin // @[DataType.scala 40:26]
        reg_uop_exc <= 3'h0;
      end else begin
        reg_uop_exc <= io_in_uop_exc;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      reg_uop_pc <= 64'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_flush) begin // @[DataType.scala 40:26]
        reg_uop_pc <= 64'h0;
      end else begin
        reg_uop_pc <= io_in_uop_pc;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      reg_uop_npc <= 64'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_flush) begin // @[DataType.scala 40:26]
        reg_uop_npc <= 64'h0;
      end else begin
        reg_uop_npc <= io_in_uop_npc;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      reg_uop_instr <= 32'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_flush) begin // @[DataType.scala 40:26]
        reg_uop_instr <= 32'h0;
      end else begin
        reg_uop_instr <= io_in_uop_instr;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      reg_uop_fu <= 3'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_flush) begin // @[DataType.scala 40:26]
        reg_uop_fu <= 3'h0;
      end else begin
        reg_uop_fu <= io_in_uop_fu;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      reg_uop_alu_op <= 4'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_flush) begin // @[DataType.scala 40:26]
        reg_uop_alu_op <= 4'h0;
      end else begin
        reg_uop_alu_op <= io_in_uop_alu_op;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      reg_uop_jmp_op <= 2'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_flush) begin // @[DataType.scala 40:26]
        reg_uop_jmp_op <= 2'h0;
      end else begin
        reg_uop_jmp_op <= io_in_uop_jmp_op;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      reg_uop_mdu_op <= 4'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_flush) begin // @[DataType.scala 40:26]
        reg_uop_mdu_op <= 4'h0;
      end else begin
        reg_uop_mdu_op <= io_in_uop_mdu_op;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      reg_uop_lsu_op <= 5'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_flush) begin // @[DataType.scala 40:26]
        reg_uop_lsu_op <= 5'h0;
      end else begin
        reg_uop_lsu_op <= io_in_uop_lsu_op;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      reg_uop_mem_len <= 2'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_flush) begin // @[DataType.scala 40:26]
        reg_uop_mem_len <= 2'h0;
      end else begin
        reg_uop_mem_len <= io_in_uop_mem_len;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      reg_uop_csr_op <= 2'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_flush) begin // @[DataType.scala 40:26]
        reg_uop_csr_op <= 2'h0;
      end else begin
        reg_uop_csr_op <= io_in_uop_csr_op;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      reg_uop_sys_op <= 3'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_flush) begin // @[DataType.scala 40:26]
        reg_uop_sys_op <= 3'h0;
      end else begin
        reg_uop_sys_op <= io_in_uop_sys_op;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      reg_uop_rd_index <= 5'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_flush) begin // @[DataType.scala 40:26]
        reg_uop_rd_index <= 5'h0;
      end else begin
        reg_uop_rd_index <= io_in_uop_rd_index;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      reg_uop_rd_wen <= 1'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_flush) begin // @[DataType.scala 40:26]
        reg_uop_rd_wen <= 1'h0;
      end else begin
        reg_uop_rd_wen <= io_in_uop_rd_wen;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      reg_uop_imm <= 32'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_flush) begin // @[DataType.scala 40:26]
        reg_uop_imm <= 32'h0;
      end else begin
        reg_uop_imm <= io_in_uop_imm;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      reg_uop_dw <= 1'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_flush) begin // @[DataType.scala 40:26]
        reg_uop_dw <= 1'h0;
      end else begin
        reg_uop_dw <= io_in_uop_dw;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      reg_rs1_data <= 64'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_flush) begin // @[DataType.scala 40:26]
        reg_rs1_data <= 64'h0;
      end else begin
        reg_rs1_data <= io_in_rs1_data;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      reg_rs2_data <= 64'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_flush) begin // @[DataType.scala 40:26]
        reg_rs2_data <= 64'h0;
      end else begin
        reg_rs2_data <= io_in_rs2_data;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      reg_rs2_data_from_rf <= 64'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_flush) begin // @[DataType.scala 40:26]
        reg_rs2_data_from_rf <= 64'h0;
      end else begin
        reg_rs2_data_from_rf <= io_in_rs2_data_from_rf;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      reg_bp_npc <= 64'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_flush) begin // @[DataType.scala 40:26]
        reg_bp_npc <= 64'h0;
      end else begin
        reg_bp_npc <= io_in_bp_npc;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_uop_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  reg_uop_exc = _RAND_1[2:0];
  _RAND_2 = {2{`RANDOM}};
  reg_uop_pc = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  reg_uop_npc = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  reg_uop_instr = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  reg_uop_fu = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  reg_uop_alu_op = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  reg_uop_jmp_op = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  reg_uop_mdu_op = _RAND_8[3:0];
  _RAND_9 = {1{`RANDOM}};
  reg_uop_lsu_op = _RAND_9[4:0];
  _RAND_10 = {1{`RANDOM}};
  reg_uop_mem_len = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  reg_uop_csr_op = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  reg_uop_sys_op = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  reg_uop_rd_index = _RAND_13[4:0];
  _RAND_14 = {1{`RANDOM}};
  reg_uop_rd_wen = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  reg_uop_imm = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  reg_uop_dw = _RAND_16[0:0];
  _RAND_17 = {2{`RANDOM}};
  reg_rs1_data = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  reg_rs2_data = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  reg_rs2_data_from_rf = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  reg_bp_npc = _RAND_20[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ALU(
  input  [3:0]  io_uop_alu_op,
  input  [1:0]  io_uop_jmp_op,
  input         io_uop_dw,
  input  [63:0] io_in1,
  input  [63:0] io_in2,
  output [63:0] io_out,
  output [63:0] io_adder_out,
  output        io_cmp_out
);
  wire  is_sub = io_uop_alu_op[3]; // @[ALU.scala 19:24]
  wire  is_cmp = io_uop_alu_op >= 4'hc; // @[ALU.scala 20:25]
  wire  cmp_unsigned = io_uop_alu_op[1]; // @[ALU.scala 21:24]
  wire  cmp_inverted = io_uop_alu_op[0]; // @[ALU.scala 22:24]
  wire  cmp_eq = ~is_sub; // @[ALU.scala 23:22]
  wire [63:0] _in2_inv_T = ~io_in2; // @[ALU.scala 26:34]
  wire [63:0] in2_inv = is_sub ? _in2_inv_T : io_in2; // @[ALU.scala 26:24]
  wire [63:0] in1_xor_in2 = io_in1 ^ in2_inv; // @[ALU.scala 27:28]
  wire [63:0] _io_adder_out_T_1 = io_in1 + in2_inv; // @[ALU.scala 28:26]
  wire [63:0] _GEN_1 = {{63'd0}, is_sub}; // @[ALU.scala 28:36]
  wire  _slt_T_2 = io_in1[63] == io_in2[63]; // @[ALU.scala 32:22]
  wire  _slt_T_6 = cmp_unsigned ? io_in2[63] : io_in1[63]; // @[ALU.scala 34:8]
  wire  slt = _slt_T_2 ? io_adder_out[63] : _slt_T_6; // @[ALU.scala 31:16]
  wire  _io_cmp_out_T_1 = cmp_eq ? in1_xor_in2 == 64'h0 : slt; // @[ALU.scala 36:35]
  wire  _T_1 = is_sub & io_in1[31]; // @[ALU.scala 43:40]
  wire [31:0] _T_3 = _T_1 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [31:0] _T_5 = io_uop_dw ? io_in1[63:32] : _T_3; // @[ALU.scala 44:27]
  wire  _T_7 = io_in2[5] & io_uop_dw; // @[ALU.scala 45:38]
  wire [5:0] shamt = {_T_7,io_in2[4:0]}; // @[Cat.scala 33:92]
  wire [63:0] shin_r = {_T_5,io_in1[31:0]}; // @[Cat.scala 33:92]
  wire  _shin_T_2 = io_uop_alu_op == 4'h5 | io_uop_alu_op == 4'hb; // @[ALU.scala 48:43]
  wire [63:0] _GEN_2 = {{32'd0}, shin_r[63:32]}; // @[Bitwise.scala 108:31]
  wire [63:0] _shin_T_6 = _GEN_2 & 64'hffffffff; // @[Bitwise.scala 108:31]
  wire [63:0] _shin_T_8 = {shin_r[31:0], 32'h0}; // @[Bitwise.scala 108:70]
  wire [63:0] _shin_T_10 = _shin_T_8 & 64'hffffffff00000000; // @[Bitwise.scala 108:80]
  wire [63:0] _shin_T_11 = _shin_T_6 | _shin_T_10; // @[Bitwise.scala 108:39]
  wire [63:0] _GEN_3 = {{16'd0}, _shin_T_11[63:16]}; // @[Bitwise.scala 108:31]
  wire [63:0] _shin_T_16 = _GEN_3 & 64'hffff0000ffff; // @[Bitwise.scala 108:31]
  wire [63:0] _shin_T_18 = {_shin_T_11[47:0], 16'h0}; // @[Bitwise.scala 108:70]
  wire [63:0] _shin_T_20 = _shin_T_18 & 64'hffff0000ffff0000; // @[Bitwise.scala 108:80]
  wire [63:0] _shin_T_21 = _shin_T_16 | _shin_T_20; // @[Bitwise.scala 108:39]
  wire [63:0] _GEN_4 = {{8'd0}, _shin_T_21[63:8]}; // @[Bitwise.scala 108:31]
  wire [63:0] _shin_T_26 = _GEN_4 & 64'hff00ff00ff00ff; // @[Bitwise.scala 108:31]
  wire [63:0] _shin_T_28 = {_shin_T_21[55:0], 8'h0}; // @[Bitwise.scala 108:70]
  wire [63:0] _shin_T_30 = _shin_T_28 & 64'hff00ff00ff00ff00; // @[Bitwise.scala 108:80]
  wire [63:0] _shin_T_31 = _shin_T_26 | _shin_T_30; // @[Bitwise.scala 108:39]
  wire [63:0] _GEN_5 = {{4'd0}, _shin_T_31[63:4]}; // @[Bitwise.scala 108:31]
  wire [63:0] _shin_T_36 = _GEN_5 & 64'hf0f0f0f0f0f0f0f; // @[Bitwise.scala 108:31]
  wire [63:0] _shin_T_38 = {_shin_T_31[59:0], 4'h0}; // @[Bitwise.scala 108:70]
  wire [63:0] _shin_T_40 = _shin_T_38 & 64'hf0f0f0f0f0f0f0f0; // @[Bitwise.scala 108:80]
  wire [63:0] _shin_T_41 = _shin_T_36 | _shin_T_40; // @[Bitwise.scala 108:39]
  wire [63:0] _GEN_6 = {{2'd0}, _shin_T_41[63:2]}; // @[Bitwise.scala 108:31]
  wire [63:0] _shin_T_46 = _GEN_6 & 64'h3333333333333333; // @[Bitwise.scala 108:31]
  wire [63:0] _shin_T_48 = {_shin_T_41[61:0], 2'h0}; // @[Bitwise.scala 108:70]
  wire [63:0] _shin_T_50 = _shin_T_48 & 64'hcccccccccccccccc; // @[Bitwise.scala 108:80]
  wire [63:0] _shin_T_51 = _shin_T_46 | _shin_T_50; // @[Bitwise.scala 108:39]
  wire [63:0] _GEN_7 = {{1'd0}, _shin_T_51[63:1]}; // @[Bitwise.scala 108:31]
  wire [63:0] _shin_T_56 = _GEN_7 & 64'h5555555555555555; // @[Bitwise.scala 108:31]
  wire [63:0] _shin_T_58 = {_shin_T_51[62:0], 1'h0}; // @[Bitwise.scala 108:70]
  wire [63:0] _shin_T_60 = _shin_T_58 & 64'haaaaaaaaaaaaaaaa; // @[Bitwise.scala 108:80]
  wire [63:0] _shin_T_61 = _shin_T_56 | _shin_T_60; // @[Bitwise.scala 108:39]
  wire [63:0] shin = io_uop_alu_op == 4'h5 | io_uop_alu_op == 4'hb ? shin_r : _shin_T_61; // @[ALU.scala 48:20]
  wire  _shout_r_T_1 = is_sub & shin[63]; // @[ALU.scala 49:29]
  wire [64:0] _shout_r_T_3 = {_shout_r_T_1,shin}; // @[ALU.scala 49:53]
  wire [64:0] _shout_r_T_4 = $signed(_shout_r_T_3) >>> shamt; // @[ALU.scala 49:60]
  wire [63:0] shout_r = _shout_r_T_4[63:0]; // @[ALU.scala 49:69]
  wire [63:0] _GEN_8 = {{32'd0}, shout_r[63:32]}; // @[Bitwise.scala 108:31]
  wire [63:0] _shout_l_T_3 = _GEN_8 & 64'hffffffff; // @[Bitwise.scala 108:31]
  wire [63:0] _shout_l_T_5 = {shout_r[31:0], 32'h0}; // @[Bitwise.scala 108:70]
  wire [63:0] _shout_l_T_7 = _shout_l_T_5 & 64'hffffffff00000000; // @[Bitwise.scala 108:80]
  wire [63:0] _shout_l_T_8 = _shout_l_T_3 | _shout_l_T_7; // @[Bitwise.scala 108:39]
  wire [63:0] _GEN_9 = {{16'd0}, _shout_l_T_8[63:16]}; // @[Bitwise.scala 108:31]
  wire [63:0] _shout_l_T_13 = _GEN_9 & 64'hffff0000ffff; // @[Bitwise.scala 108:31]
  wire [63:0] _shout_l_T_15 = {_shout_l_T_8[47:0], 16'h0}; // @[Bitwise.scala 108:70]
  wire [63:0] _shout_l_T_17 = _shout_l_T_15 & 64'hffff0000ffff0000; // @[Bitwise.scala 108:80]
  wire [63:0] _shout_l_T_18 = _shout_l_T_13 | _shout_l_T_17; // @[Bitwise.scala 108:39]
  wire [63:0] _GEN_10 = {{8'd0}, _shout_l_T_18[63:8]}; // @[Bitwise.scala 108:31]
  wire [63:0] _shout_l_T_23 = _GEN_10 & 64'hff00ff00ff00ff; // @[Bitwise.scala 108:31]
  wire [63:0] _shout_l_T_25 = {_shout_l_T_18[55:0], 8'h0}; // @[Bitwise.scala 108:70]
  wire [63:0] _shout_l_T_27 = _shout_l_T_25 & 64'hff00ff00ff00ff00; // @[Bitwise.scala 108:80]
  wire [63:0] _shout_l_T_28 = _shout_l_T_23 | _shout_l_T_27; // @[Bitwise.scala 108:39]
  wire [63:0] _GEN_11 = {{4'd0}, _shout_l_T_28[63:4]}; // @[Bitwise.scala 108:31]
  wire [63:0] _shout_l_T_33 = _GEN_11 & 64'hf0f0f0f0f0f0f0f; // @[Bitwise.scala 108:31]
  wire [63:0] _shout_l_T_35 = {_shout_l_T_28[59:0], 4'h0}; // @[Bitwise.scala 108:70]
  wire [63:0] _shout_l_T_37 = _shout_l_T_35 & 64'hf0f0f0f0f0f0f0f0; // @[Bitwise.scala 108:80]
  wire [63:0] _shout_l_T_38 = _shout_l_T_33 | _shout_l_T_37; // @[Bitwise.scala 108:39]
  wire [63:0] _GEN_12 = {{2'd0}, _shout_l_T_38[63:2]}; // @[Bitwise.scala 108:31]
  wire [63:0] _shout_l_T_43 = _GEN_12 & 64'h3333333333333333; // @[Bitwise.scala 108:31]
  wire [63:0] _shout_l_T_45 = {_shout_l_T_38[61:0], 2'h0}; // @[Bitwise.scala 108:70]
  wire [63:0] _shout_l_T_47 = _shout_l_T_45 & 64'hcccccccccccccccc; // @[Bitwise.scala 108:80]
  wire [63:0] _shout_l_T_48 = _shout_l_T_43 | _shout_l_T_47; // @[Bitwise.scala 108:39]
  wire [63:0] _GEN_13 = {{1'd0}, _shout_l_T_48[63:1]}; // @[Bitwise.scala 108:31]
  wire [63:0] _shout_l_T_53 = _GEN_13 & 64'h5555555555555555; // @[Bitwise.scala 108:31]
  wire [63:0] _shout_l_T_55 = {_shout_l_T_48[62:0], 1'h0}; // @[Bitwise.scala 108:70]
  wire [63:0] _shout_l_T_57 = _shout_l_T_55 & 64'haaaaaaaaaaaaaaaa; // @[Bitwise.scala 108:80]
  wire [63:0] shout_l = _shout_l_T_53 | _shout_l_T_57; // @[Bitwise.scala 108:39]
  wire [63:0] _shout_T_3 = _shin_T_2 ? shout_r : 64'h0; // @[ALU.scala 51:18]
  wire [63:0] _shout_T_5 = io_uop_alu_op == 4'h1 ? shout_l : 64'h0; // @[ALU.scala 52:8]
  wire [63:0] shout = _shout_T_3 | _shout_T_5; // @[ALU.scala 51:81]
  wire  _logic_T_1 = io_uop_alu_op == 4'h6; // @[ALU.scala 55:47]
  wire [63:0] _logic_T_3 = io_uop_alu_op == 4'h4 | io_uop_alu_op == 4'h6 ? in1_xor_in2 : 64'h0; // @[ALU.scala 55:18]
  wire [63:0] _logic_T_7 = io_in1 & io_in2; // @[ALU.scala 56:63]
  wire [63:0] _logic_T_8 = _logic_T_1 | io_uop_alu_op == 4'h7 ? _logic_T_7 : 64'h0; // @[ALU.scala 56:8]
  wire [63:0] logic_ = _logic_T_3 | _logic_T_8; // @[ALU.scala 55:84]
  wire  _shift_logic_T = is_cmp & slt; // @[ALU.scala 57:29]
  wire [63:0] _GEN_14 = {{63'd0}, _shift_logic_T}; // @[ALU.scala 57:37]
  wire [63:0] _shift_logic_T_1 = _GEN_14 | logic_; // @[ALU.scala 57:37]
  wire [63:0] shift_logic = _shift_logic_T_1 | shout; // @[ALU.scala 57:45]
  wire [63:0] out = io_uop_alu_op == 4'h0 | io_uop_alu_op == 4'ha ? io_adder_out : shift_logic; // @[ALU.scala 58:24]
  wire [31:0] _io_out_T_2 = out[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _io_out_T_4 = {_io_out_T_2,out[31:0]}; // @[Cat.scala 33:92]
  assign io_out = ~io_uop_dw ? _io_out_T_4 : out; // @[ALU.scala 60:10 63:{22,31}]
  assign io_adder_out = _io_adder_out_T_1 + _GEN_1; // @[ALU.scala 28:36]
  assign io_cmp_out = cmp_inverted ^ _io_cmp_out_T_1; // @[ALU.scala 36:30]
endmodule
module LSU(
  input         clock,
  input         reset,
  input  [4:0]  io_uop_lsu_op,
  input  [1:0]  io_uop_mem_len,
  input         io_is_mem,
  input         io_is_store,
  input         io_is_amo,
  input  [63:0] io_addr,
  input  [63:0] io_wdata,
  output [63:0] io_rdata,
  output        io_valid,
  output [3:0]  io_exc_code,
  input         io_dmem_req_ready,
  output        io_dmem_req_valid,
  output [38:0] io_dmem_req_bits_addr,
  output [63:0] io_dmem_req_bits_wdata,
  output [7:0]  io_dmem_req_bits_wmask,
  output        io_dmem_req_bits_wen,
  output [1:0]  io_dmem_req_bits_len,
  output        io_dmem_req_bits_lrsc,
  output [4:0]  io_dmem_req_bits_amo,
  output        io_dmem_resp_ready,
  input         io_dmem_resp_valid,
  input  [63:0] io_dmem_resp_bits_rdata,
  input         io_dmem_resp_bits_page_fault,
  input         io_dmem_resp_bits_access_fault,
  output        io_ready
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[LSU.scala 31:58]
  wire [2:0] addr_offset = io_addr[2:0]; // @[LSU.scala 33:28]
  wire [5:0] _wdata_T = {addr_offset, 3'h0}; // @[LSU.scala 35:41]
  wire [126:0] _GEN_7 = {{63'd0}, io_wdata}; // @[LSU.scala 35:25]
  wire [126:0] _wdata_T_1 = _GEN_7 << _wdata_T; // @[LSU.scala 35:25]
  wire [7:0] _wmask_T_1 = 2'h1 == io_uop_mem_len ? 8'h3 : 8'h1; // @[Mux.scala 81:58]
  wire [7:0] _wmask_T_3 = 2'h2 == io_uop_mem_len ? 8'hf : _wmask_T_1; // @[Mux.scala 81:58]
  wire [7:0] _wmask_T_5 = 2'h3 == io_uop_mem_len ? 8'hff : _wmask_T_3; // @[Mux.scala 81:58]
  wire [14:0] _GEN_8 = {{7'd0}, _wmask_T_5}; // @[LSU.scala 45:5]
  wire [14:0] _wmask_T_6 = _GEN_8 << addr_offset; // @[LSU.scala 45:5]
  wire  _io_dmem_req_bits_wen_T = io_is_store | io_is_amo; // @[LSU.scala 51:33]
  wire  _io_dmem_req_bits_lrsc_T_2 = ~io_uop_lsu_op[4]; // @[Constant.scala 85:32]
  wire  _io_dmem_resp_ready_T = state == 2'h2; // @[LSU.scala 55:28]
  wire  _misaligned_T_3 = io_addr[1:0] != 2'h0; // @[LSU.scala 63:42]
  wire  _misaligned_T_5 = addr_offset != 3'h0; // @[LSU.scala 64:42]
  wire  _misaligned_T_9 = 2'h2 == io_uop_mem_len ? _misaligned_T_3 : 2'h1 == io_uop_mem_len & io_addr[0]; // @[Mux.scala 81:58]
  wire  misaligned = 2'h3 == io_uop_mem_len ? _misaligned_T_5 : _misaligned_T_9; // @[Mux.scala 81:58]
  wire  _T_2 = io_dmem_req_ready & io_dmem_req_valid; // @[Decoupled.scala 51:35]
  wire  _T_4 = io_dmem_resp_ready & io_dmem_resp_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _state_T_2 = io_dmem_resp_bits_page_fault | io_dmem_resp_bits_access_fault ? 2'h3 : 2'h0; // @[LSU.scala 81:21]
  wire [1:0] _GEN_2 = _T_4 ? _state_T_2 : state; // @[LSU.scala 80:23 81:15 31:58]
  wire [1:0] _GEN_3 = 2'h3 == state ? 2'h0 : state; // @[LSU.scala 68:17 85:13 31:58]
  wire [63:0] resp_data = io_dmem_resp_bits_rdata >> _wdata_T; // @[LSU.scala 89:35]
  wire  _sign_T_5 = _io_dmem_req_bits_lrsc_T_2 & io_uop_lsu_op[1]; // @[Constant.scala 83:45]
  wire  _sign_T_8 = _sign_T_5 & io_uop_lsu_op[2]; // @[Constant.scala 84:42]
  wire  _sign_T_16 = 2'h1 == io_uop_mem_len ? resp_data[15] : 2'h0 == io_uop_mem_len & resp_data[7]; // @[Mux.scala 81:58]
  wire  _sign_T_18 = 2'h2 == io_uop_mem_len ? resp_data[31] : _sign_T_16; // @[Mux.scala 81:58]
  wire  sign = ~_sign_T_8 & _sign_T_18; // @[LSU.scala 90:37]
  wire [55:0] _rdata_T_1 = sign ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _rdata_T_3 = {_rdata_T_1,resp_data[7:0]}; // @[Cat.scala 33:92]
  wire [47:0] _rdata_T_5 = sign ? 48'hffffffffffff : 48'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _rdata_T_7 = {_rdata_T_5,resp_data[15:0]}; // @[Cat.scala 33:92]
  wire [31:0] _rdata_T_9 = sign ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _rdata_T_11 = {_rdata_T_9,resp_data[31:0]}; // @[Cat.scala 33:92]
  wire [63:0] _rdata_T_13 = 2'h1 == io_uop_mem_len ? _rdata_T_7 : _rdata_T_3; // @[Mux.scala 81:58]
  wire [63:0] _rdata_T_15 = 2'h2 == io_uop_mem_len ? _rdata_T_11 : _rdata_T_13; // @[Mux.scala 81:58]
  wire  _io_valid_T_7 = state == 2'h3; // @[LSU.scala 111:115]
  reg  exc_code_REG; // @[LSU.scala 131:20]
  wire [3:0] _exc_code_T_1 = exc_code_REG ? 4'h7 : 4'hf; // @[LSU.scala 131:12]
  wire [3:0] _exc_code_T_2 = misaligned ? 4'h6 : _exc_code_T_1; // @[LSU.scala 128:10]
  reg  exc_code_REG_1; // @[LSU.scala 136:20]
  wire [3:0] _exc_code_T_3 = exc_code_REG_1 ? 4'h5 : 4'hd; // @[LSU.scala 136:12]
  wire [3:0] _exc_code_T_4 = misaligned ? 4'h4 : _exc_code_T_3; // @[LSU.scala 133:10]
  wire [3:0] exc_code = _io_dmem_req_bits_wen_T ? _exc_code_T_2 : _exc_code_T_4; // @[LSU.scala 126:8]
  assign io_rdata = 2'h3 == io_uop_mem_len ? resp_data : _rdata_T_15; // @[Mux.scala 81:58]
  assign io_valid = _io_dmem_resp_ready_T & (_T_4 & ~io_dmem_resp_bits_page_fault & ~io_dmem_resp_bits_access_fault) |
    state == 2'h3; // @[LSU.scala 111:105]
  assign io_exc_code = _io_valid_T_7 ? exc_code : 4'h0; // @[LSU.scala 139:21]
  assign io_dmem_req_valid = state == 2'h1; // @[LSU.scala 54:28]
  assign io_dmem_req_bits_addr = io_addr[38:0]; // @[LSU.scala 47:18]
  assign io_dmem_req_bits_wdata = _wdata_T_1[63:0]; // @[LSU.scala 35:47]
  assign io_dmem_req_bits_wmask = _wmask_T_6[7:0]; // @[LSU.scala 45:20]
  assign io_dmem_req_bits_wen = io_is_store | io_is_amo; // @[LSU.scala 51:33]
  assign io_dmem_req_bits_len = io_uop_mem_len; // @[LSU.scala 50:18]
  assign io_dmem_req_bits_lrsc = ~io_uop_lsu_op[4] & io_uop_lsu_op[3]; // @[Constant.scala 85:45]
  assign io_dmem_req_bits_amo = io_uop_lsu_op; // @[LSU.scala 53:18]
  assign io_dmem_resp_ready = state == 2'h2; // @[LSU.scala 55:28]
  assign io_ready = state == 2'h0 & ~io_is_mem | io_valid; // @[LSU.scala 113:52]
  always @(posedge clock) begin
    if (reset) begin // @[LSU.scala 31:58]
      state <= 2'h0; // @[LSU.scala 31:58]
    end else if (2'h0 == state) begin // @[LSU.scala 68:17]
      if (io_is_mem) begin // @[LSU.scala 70:23]
        if (misaligned) begin // @[LSU.scala 71:21]
          state <= 2'h3;
        end else begin
          state <= 2'h1;
        end
      end
    end else if (2'h1 == state) begin // @[LSU.scala 68:17]
      if (_T_2) begin // @[LSU.scala 75:22]
        state <= 2'h2; // @[LSU.scala 76:15]
      end
    end else if (2'h2 == state) begin // @[LSU.scala 68:17]
      state <= _GEN_2;
    end else begin
      state <= _GEN_3;
    end
    exc_code_REG <= io_dmem_resp_bits_access_fault; // @[LSU.scala 131:20]
    exc_code_REG_1 <= io_dmem_resp_bits_access_fault; // @[LSU.scala 136:20]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  exc_code_REG = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  exc_code_REG_1 = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MulDiv(
  input         clock,
  input         reset,
  output        io_req_ready,
  input         io_req_valid,
  input  [3:0]  io_req_bits_fn,
  input         io_req_bits_dw,
  input  [63:0] io_req_bits_in1,
  input  [63:0] io_req_bits_in2,
  input         io_resp_ready,
  output        io_resp_valid,
  output [63:0] io_resp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [95:0] _RAND_6;
  reg [159:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] state; // @[Multiplier.scala 48:22]
  reg  req_dw; // @[Multiplier.scala 50:16]
  reg [6:0] count; // @[Multiplier.scala 51:18]
  reg  neg_out; // @[Multiplier.scala 54:20]
  reg  isHi; // @[Multiplier.scala 55:17]
  reg  resHi; // @[Multiplier.scala 56:18]
  reg [64:0] divisor; // @[Multiplier.scala 57:20]
  reg [129:0] remainder; // @[Multiplier.scala 58:22]
  wire [2:0] decoded_plaInput = io_req_bits_fn[2:0]; // @[decoder.scala 40:16 pla.scala 77:22]
  wire [2:0] decoded_invInputs = ~decoded_plaInput; // @[pla.scala 78:21]
  wire  decoded_andMatrixInput_0 = decoded_invInputs[0]; // @[pla.scala 91:29]
  wire  _decoded_T = &decoded_andMatrixInput_0; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_0_1 = decoded_invInputs[2]; // @[pla.scala 91:29]
  wire  _decoded_T_1 = &decoded_andMatrixInput_0_1; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_0_2 = decoded_invInputs[1]; // @[pla.scala 91:29]
  wire [1:0] _decoded_T_2 = {decoded_andMatrixInput_0_2,decoded_andMatrixInput_0_1}; // @[Cat.scala 33:92]
  wire  _decoded_T_3 = &_decoded_T_2; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_0_3 = decoded_plaInput[0]; // @[pla.scala 90:45]
  wire [1:0] _decoded_T_4 = {decoded_andMatrixInput_0_3,decoded_andMatrixInput_0_1}; // @[Cat.scala 33:92]
  wire  _decoded_T_5 = &_decoded_T_4; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_0_4 = decoded_plaInput[1]; // @[pla.scala 90:45]
  wire  _decoded_T_6 = &decoded_andMatrixInput_0_4; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_1_2 = decoded_plaInput[2]; // @[pla.scala 90:45]
  wire [1:0] _decoded_T_7 = {decoded_andMatrixInput_0,decoded_andMatrixInput_1_2}; // @[Cat.scala 33:92]
  wire  _decoded_T_8 = &_decoded_T_7; // @[pla.scala 98:74]
  wire [1:0] _decoded_orMatrixOutputs_T = {_decoded_T_3,_decoded_T_8}; // @[Cat.scala 33:92]
  wire  _decoded_orMatrixOutputs_T_1 = |_decoded_orMatrixOutputs_T; // @[pla.scala 114:39]
  wire [1:0] _decoded_orMatrixOutputs_T_2 = {_decoded_T,_decoded_T_3}; // @[Cat.scala 33:92]
  wire  _decoded_orMatrixOutputs_T_3 = |_decoded_orMatrixOutputs_T_2; // @[pla.scala 114:39]
  wire [1:0] _decoded_orMatrixOutputs_T_4 = {_decoded_T_5,_decoded_T_6}; // @[Cat.scala 33:92]
  wire  _decoded_orMatrixOutputs_T_5 = |_decoded_orMatrixOutputs_T_4; // @[pla.scala 114:39]
  wire  _decoded_orMatrixOutputs_T_6 = |_decoded_T_1; // @[pla.scala 114:39]
  wire [3:0] decoded_orMatrixOutputs = {_decoded_orMatrixOutputs_T_6,_decoded_orMatrixOutputs_T_5,
    _decoded_orMatrixOutputs_T_3,_decoded_orMatrixOutputs_T_1}; // @[Cat.scala 33:92]
  wire [3:0] decoded_invMatrixOutputs = {decoded_orMatrixOutputs[3],decoded_orMatrixOutputs[2],decoded_orMatrixOutputs[1
    ],decoded_orMatrixOutputs[0]}; // @[Cat.scala 33:92]
  wire  cmdMul = decoded_invMatrixOutputs[3]; // @[Decode.scala 50:77]
  wire  cmdHi = decoded_invMatrixOutputs[2]; // @[Decode.scala 50:77]
  wire  lhsSigned = decoded_invMatrixOutputs[1]; // @[Decode.scala 50:77]
  wire  rhsSigned = decoded_invMatrixOutputs[0]; // @[Decode.scala 50:77]
  wire  _T_4 = ~io_req_bits_dw; // @[Multiplier.scala 75:60]
  wire  _sign_T_2 = _T_4 ? io_req_bits_in1[31] : io_req_bits_in1[63]; // @[Multiplier.scala 78:29]
  wire  lhs_sign = lhsSigned & _sign_T_2; // @[Multiplier.scala 78:23]
  wire [31:0] _hi_T_1 = lhs_sign ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [31:0] hi = _T_4 ? _hi_T_1 : io_req_bits_in1[63:32]; // @[Multiplier.scala 79:17]
  wire [63:0] lhs_in = {hi,io_req_bits_in1[31:0]}; // @[Cat.scala 33:92]
  wire  _sign_T_5 = _T_4 ? io_req_bits_in2[31] : io_req_bits_in2[63]; // @[Multiplier.scala 78:29]
  wire  rhs_sign = rhsSigned & _sign_T_5; // @[Multiplier.scala 78:23]
  wire [31:0] _hi_T_4 = rhs_sign ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [31:0] hi_1 = _T_4 ? _hi_T_4 : io_req_bits_in2[63:32]; // @[Multiplier.scala 79:17]
  wire [64:0] subtractor = remainder[128:64] - divisor; // @[Multiplier.scala 85:37]
  wire [63:0] result = resHi ? remainder[128:65] : remainder[63:0]; // @[Multiplier.scala 86:19]
  wire [63:0] negated_remainder = 64'h0 - result; // @[Multiplier.scala 87:27]
  wire [129:0] _GEN_0 = remainder[63] ? {{66'd0}, negated_remainder} : remainder; // @[Multiplier.scala 90:27 91:17 58:22]
  wire [129:0] _GEN_2 = state == 3'h1 ? _GEN_0 : remainder; // @[Multiplier.scala 58:22 89:57]
  wire [2:0] _GEN_4 = state == 3'h1 ? 3'h3 : state; // @[Multiplier.scala 89:57 96:11 48:22]
  wire [2:0] _GEN_6 = state == 3'h5 ? 3'h7 : _GEN_4; // @[Multiplier.scala 100:11 98:57]
  wire  _GEN_7 = state == 3'h5 ? 1'h0 : resHi; // @[Multiplier.scala 101:11 56:18 98:57]
  wire [128:0] mulReg = {remainder[129:65],remainder[63:0]}; // @[Cat.scala 33:92]
  wire  mplierSign = remainder[64]; // @[Multiplier.scala 105:31]
  wire [63:0] mplier = mulReg[63:0]; // @[Multiplier.scala 106:24]
  wire [64:0] accum = mulReg[128:64]; // @[Multiplier.scala 107:37]
  wire [1:0] _prod_T_2 = {mplierSign,mplier[0]}; // @[Multiplier.scala 109:60]
  wire [66:0] _prod_T_3 = $signed(_prod_T_2) * $signed(divisor); // @[Multiplier.scala 109:67]
  wire [66:0] _GEN_35 = {{2{accum[64]}},accum}; // @[Multiplier.scala 109:76]
  wire [66:0] nextMulReg_hi = $signed(_prod_T_3) + $signed(_GEN_35); // @[Cat.scala 33:92]
  wire [129:0] nextMulReg = {nextMulReg_hi,mplier[63:1]}; // @[Cat.scala 33:92]
  wire  nextMplierSign = count == 7'h3e & neg_out; // @[Multiplier.scala 111:61]
  wire  _eOut_T_4 = ~isHi; // @[Multiplier.scala 115:7]
  wire [128:0] nextMulReg1 = {nextMulReg[128:64],nextMulReg[63:0]}; // @[Cat.scala 33:92]
  wire [129:0] _remainder_T_2 = {nextMulReg1[128:64],nextMplierSign,nextMulReg1[63:0]}; // @[Cat.scala 33:92]
  wire [6:0] _count_T_1 = count + 7'h1; // @[Multiplier.scala 120:20]
  wire [2:0] _GEN_8 = count == 7'h3f ? 3'h6 : _GEN_6; // @[Multiplier.scala 121:55 122:13]
  wire  _GEN_9 = count == 7'h3f ? isHi : _GEN_7; // @[Multiplier.scala 121:55 123:13]
  wire [2:0] _GEN_12 = state == 3'h2 ? _GEN_8 : _GEN_6; // @[Multiplier.scala 103:50]
  wire  _GEN_13 = state == 3'h2 ? _GEN_9 : _GEN_7; // @[Multiplier.scala 103:50]
  wire  unrolls_less = subtractor[64]; // @[Multiplier.scala 130:28]
  wire [63:0] _unrolls_T_2 = unrolls_less ? remainder[127:64] : subtractor[63:0]; // @[Multiplier.scala 131:14]
  wire  _unrolls_T_4 = ~unrolls_less; // @[Multiplier.scala 131:67]
  wire [128:0] unrolls_0 = {_unrolls_T_2,remainder[63:0],_unrolls_T_4}; // @[Cat.scala 33:92]
  wire [2:0] _state_T = neg_out ? 3'h5 : 3'h7; // @[Multiplier.scala 136:19]
  wire [2:0] _GEN_14 = count == 7'h40 ? _state_T : _GEN_12; // @[Multiplier.scala 135:42 136:13]
  wire  divby0 = count == 7'h0 & _unrolls_T_4; // @[Multiplier.scala 143:32]
  wire  _T_23 = io_req_ready & io_req_valid; // @[Decoupled.scala 51:35]
  wire [5:0] _count_T_7 = cmdMul & _T_4 ? 6'h20 : 6'h0; // @[Multiplier.scala 165:38]
  wire [64:0] _divisor_T = {rhs_sign,hi_1,io_req_bits_in2[31:0]}; // @[Cat.scala 33:92]
  wire [2:0] _outMul_T_1 = state & 3'h1; // @[Multiplier.scala 172:23]
  wire  outMul = _outMul_T_1 == 3'h0; // @[Multiplier.scala 172:52]
  wire  _loOut_T = ~req_dw; // @[Multiplier.scala 75:60]
  wire [31:0] loOut = _loOut_T & outMul ? result[63:32] : result[31:0]; // @[Multiplier.scala 173:18]
  wire [31:0] _hiOut_T_4 = loOut[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [31:0] hiOut = _loOut_T ? _hiOut_T_4 : result[63:32]; // @[Multiplier.scala 174:18]
  assign io_req_ready = state == 3'h0; // @[Multiplier.scala 179:25]
  assign io_resp_valid = state == 3'h6 | state == 3'h7; // @[Multiplier.scala 178:42]
  assign io_resp_bits_data = {hiOut,loOut}; // @[Cat.scala 33:92]
  always @(posedge clock) begin
    if (reset) begin // @[Multiplier.scala 48:22]
      state <= 3'h0; // @[Multiplier.scala 48:22]
    end else if (_T_23) begin // @[Multiplier.scala 161:24]
      if (cmdMul) begin // @[Multiplier.scala 162:17]
        state <= 3'h2;
      end else if (lhs_sign | rhs_sign) begin // @[Multiplier.scala 162:36]
        state <= 3'h1;
      end else begin
        state <= 3'h3;
      end
    end else if (io_resp_valid) begin // @[Multiplier.scala 158:36]
      state <= 3'h0; // @[Multiplier.scala 159:11]
    end else if (state == 3'h3) begin // @[Multiplier.scala 126:50]
      state <= _GEN_14;
    end else begin
      state <= _GEN_12;
    end
    if (_T_23) begin // @[Multiplier.scala 161:24]
      req_dw <= io_req_bits_dw; // @[Multiplier.scala 169:9]
    end
    if (_T_23) begin // @[Multiplier.scala 161:24]
      count <= {{1'd0}, _count_T_7}; // @[Multiplier.scala 165:11]
    end else if (state == 3'h3) begin // @[Multiplier.scala 126:50]
      count <= _count_T_1; // @[Multiplier.scala 141:11]
    end else if (state == 3'h2) begin // @[Multiplier.scala 103:50]
      count <= _count_T_1; // @[Multiplier.scala 120:11]
    end
    if (_T_23) begin // @[Multiplier.scala 161:24]
      if (cmdHi) begin // @[Multiplier.scala 166:19]
        neg_out <= lhs_sign;
      end else begin
        neg_out <= lhs_sign != rhs_sign;
      end
    end else if (state == 3'h3) begin // @[Multiplier.scala 126:50]
      if (divby0 & _eOut_T_4) begin // @[Multiplier.scala 156:28]
        neg_out <= 1'h0; // @[Multiplier.scala 156:38]
      end
    end
    if (_T_23) begin // @[Multiplier.scala 161:24]
      isHi <= cmdHi; // @[Multiplier.scala 163:10]
    end
    if (_T_23) begin // @[Multiplier.scala 161:24]
      resHi <= 1'h0; // @[Multiplier.scala 164:11]
    end else if (state == 3'h3) begin // @[Multiplier.scala 126:50]
      if (count == 7'h40) begin // @[Multiplier.scala 135:42]
        resHi <= isHi; // @[Multiplier.scala 137:13]
      end else begin
        resHi <= _GEN_13;
      end
    end else begin
      resHi <= _GEN_13;
    end
    if (_T_23) begin // @[Multiplier.scala 161:24]
      divisor <= _divisor_T; // @[Multiplier.scala 167:13]
    end else if (state == 3'h1) begin // @[Multiplier.scala 89:57]
      if (divisor[63]) begin // @[Multiplier.scala 93:25]
        divisor <= subtractor; // @[Multiplier.scala 94:15]
      end
    end
    if (_T_23) begin // @[Multiplier.scala 161:24]
      remainder <= {{66'd0}, lhs_in}; // @[Multiplier.scala 168:15]
    end else if (state == 3'h3) begin // @[Multiplier.scala 126:50]
      remainder <= {{1'd0}, unrolls_0}; // @[Multiplier.scala 134:15]
    end else if (state == 3'h2) begin // @[Multiplier.scala 103:50]
      remainder <= _remainder_T_2; // @[Multiplier.scala 118:15]
    end else if (state == 3'h5) begin // @[Multiplier.scala 98:57]
      remainder <= {{66'd0}, negated_remainder}; // @[Multiplier.scala 99:15]
    end else begin
      remainder <= _GEN_2;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  req_dw = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  count = _RAND_2[6:0];
  _RAND_3 = {1{`RANDOM}};
  neg_out = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  isHi = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  resHi = _RAND_5[0:0];
  _RAND_6 = {3{`RANDOM}};
  divisor = _RAND_6[64:0];
  _RAND_7 = {5{`RANDOM}};
  remainder = _RAND_7[129:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MDU(
  input         clock,
  input         reset,
  input         io_uop_valid,
  input  [3:0]  io_uop_mdu_op,
  input         io_uop_dw,
  input         io_is_mdu,
  input  [63:0] io_in1,
  input  [63:0] io_in2,
  output [63:0] io_out,
  output        io_valid,
  output        io_ready
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  rocket_mdu_clock; // @[MDU.scala 26:26]
  wire  rocket_mdu_reset; // @[MDU.scala 26:26]
  wire  rocket_mdu_io_req_ready; // @[MDU.scala 26:26]
  wire  rocket_mdu_io_req_valid; // @[MDU.scala 26:26]
  wire [3:0] rocket_mdu_io_req_bits_fn; // @[MDU.scala 26:26]
  wire  rocket_mdu_io_req_bits_dw; // @[MDU.scala 26:26]
  wire [63:0] rocket_mdu_io_req_bits_in1; // @[MDU.scala 26:26]
  wire [63:0] rocket_mdu_io_req_bits_in2; // @[MDU.scala 26:26]
  wire  rocket_mdu_io_resp_ready; // @[MDU.scala 26:26]
  wire  rocket_mdu_io_resp_valid; // @[MDU.scala 26:26]
  wire [63:0] rocket_mdu_io_resp_bits_data; // @[MDU.scala 26:26]
  reg [1:0] state; // @[MDU.scala 24:49]
  wire  _T_2 = rocket_mdu_io_req_ready & rocket_mdu_io_req_valid; // @[Decoupled.scala 51:35]
  wire  _T_4 = rocket_mdu_io_resp_ready & rocket_mdu_io_resp_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _GEN_2 = _T_4 ? 2'h0 : state; // @[MDU.scala 48:37 49:15 24:49]
  MulDiv rocket_mdu ( // @[MDU.scala 26:26]
    .clock(rocket_mdu_clock),
    .reset(rocket_mdu_reset),
    .io_req_ready(rocket_mdu_io_req_ready),
    .io_req_valid(rocket_mdu_io_req_valid),
    .io_req_bits_fn(rocket_mdu_io_req_bits_fn),
    .io_req_bits_dw(rocket_mdu_io_req_bits_dw),
    .io_req_bits_in1(rocket_mdu_io_req_bits_in1),
    .io_req_bits_in2(rocket_mdu_io_req_bits_in2),
    .io_resp_ready(rocket_mdu_io_resp_ready),
    .io_resp_valid(rocket_mdu_io_resp_valid),
    .io_resp_bits_data(rocket_mdu_io_resp_bits_data)
  );
  assign io_out = rocket_mdu_io_resp_bits_data; // @[MDU.scala 54:12]
  assign io_valid = state == 2'h2 & _T_4; // @[MDU.scala 55:34]
  assign io_ready = state == 2'h0 & ~io_is_mdu | io_valid; // @[MDU.scala 56:47]
  assign rocket_mdu_clock = clock;
  assign rocket_mdu_reset = reset;
  assign rocket_mdu_io_req_valid = state == 2'h1 & io_uop_valid & io_is_mdu; // @[MDU.scala 27:64]
  assign rocket_mdu_io_req_bits_fn = io_uop_mdu_op; // @[MDU.scala 28:30]
  assign rocket_mdu_io_req_bits_dw = io_uop_dw; // @[MDU.scala 29:30]
  assign rocket_mdu_io_req_bits_in1 = io_in1; // @[MDU.scala 30:30]
  assign rocket_mdu_io_req_bits_in2 = io_in2; // @[MDU.scala 31:30]
  assign rocket_mdu_io_resp_ready = 1'h1; // @[MDU.scala 34:30]
  always @(posedge clock) begin
    if (reset) begin // @[MDU.scala 24:49]
      state <= 2'h0; // @[MDU.scala 24:49]
    end else if (2'h0 == state) begin // @[MDU.scala 36:17]
      if (io_is_mdu) begin // @[MDU.scala 38:20]
        state <= 2'h1; // @[MDU.scala 39:15]
      end
    end else if (2'h1 == state) begin // @[MDU.scala 36:17]
      if (_T_2) begin // @[MDU.scala 43:36]
        state <= 2'h2; // @[MDU.scala 44:15]
      end
    end else if (2'h2 == state) begin // @[MDU.scala 36:17]
      state <= _GEN_2;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CSR(
  input         clock,
  input         reset,
  input         io_uop_valid,
  input  [2:0]  io_uop_exc,
  input  [63:0] io_uop_pc,
  input  [63:0] io_uop_npc,
  input  [2:0]  io_uop_fu,
  input  [2:0]  io_uop_sys_op,
  input  [11:0] io_rw_addr,
  input  [1:0]  io_rw_cmd,
  input  [63:0] io_rw_wdata,
  output [63:0] io_rw_rdata,
  output        io_rw_valid,
  output [1:0]  io_prv,
  output        io_mprv,
  output [1:0]  io_mpp,
  output        io_sv39_en,
  output [15:0] io_satp_asid,
  output [43:0] io_satp_ppn,
  output        io_sfence_vma,
  output        io_fence_i,
  output        io_jmp_packet_valid,
  output [63:0] io_jmp_packet_target,
  input  [63:0] io_lsu_addr,
  input  [3:0]  io_lsu_exc_code,
  input         io_interrupt_mtip,
  input         io_interrupt_msip,
  input         io_interrupt_meip,
  input         io_interrupt_seip,
  output        io_is_int,
  input         io_commit
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] prv; // @[CSR.scala 49:26]
  wire  mret_legal = prv == 2'h3; // @[CSR.scala 50:24]
  wire  prv_is_s = prv == 2'h1; // @[CSR.scala 51:24]
  wire  prv_is_ms = mret_legal | prv_is_s; // @[CSR.scala 52:28]
  wire  prv_is_u = prv == 2'h0; // @[CSR.scala 53:24]
  wire  _wen_T = io_rw_cmd != 2'h0; // @[CSR.scala 58:30]
  reg [63:0] mcounteren; // @[CSR.scala 477:27]
  reg [63:0] scounteren; // @[CSR.scala 208:27]
  reg  mstatus_tvm; // @[CSR.scala 117:29]
  wire  tvm_en = prv_is_s & mstatus_tvm; // @[CSR.scala 285:31]
  wire  _csr_legal_T_1 = prv_is_ms & ~tvm_en; // @[CSR.scala 300:28]
  wire  _GEN_13 = io_rw_addr == 12'h100 & prv_is_ms; // @[CSR.scala 151:39 162:15 55:30]
  wire  _GEN_41 = io_rw_addr == 12'h300 ? mret_legal : _GEN_13; // @[CSR.scala 164:39 182:15]
  wire  _GEN_45 = io_rw_addr == 12'h105 ? prv_is_ms : _GEN_41; // @[CSR.scala 194:37 199:15]
  wire  _GEN_49 = io_rw_addr == 12'h106 ? prv_is_ms : _GEN_45; // @[CSR.scala 209:42 214:15]
  wire  _GEN_53 = io_rw_addr == 12'h140 ? prv_is_ms : _GEN_49; // @[CSR.scala 224:40 229:15]
  wire  _GEN_57 = io_rw_addr == 12'h141 ? prv_is_ms : _GEN_53; // @[CSR.scala 239:36 244:15]
  wire  _GEN_61 = io_rw_addr == 12'h142 ? prv_is_ms : _GEN_57; // @[CSR.scala 254:38 259:15]
  wire  _GEN_65 = io_rw_addr == 12'h143 ? prv_is_ms : _GEN_61; // @[CSR.scala 269:37 274:15]
  wire  _GEN_77 = io_rw_addr == 12'h180 ? prv_is_ms & ~tvm_en : _GEN_65; // @[CSR.scala 291:36 300:15]
  wire  _GEN_79 = io_rw_addr == 12'hf11 ? mret_legal : _GEN_77; // @[CSR.scala 309:41 311:15]
  wire  _GEN_81 = io_rw_addr == 12'hf12 ? mret_legal : _GEN_79; // @[CSR.scala 320:39 322:15]
  wire  _GEN_83 = io_rw_addr == 12'hf13 ? mret_legal : _GEN_81; // @[CSR.scala 331:38 333:15]
  wire  _GEN_89 = io_rw_addr == 12'hf14 ? mret_legal : _GEN_83; // @[CSR.scala 344:39 350:15]
  wire  _GEN_91 = io_rw_addr == 12'h301 ? mret_legal : _GEN_89; // @[CSR.scala 361:36 363:15]
  wire  _GEN_95 = io_rw_addr == 12'h302 ? mret_legal : _GEN_91; // @[CSR.scala 373:39 378:15]
  wire  _GEN_99 = io_rw_addr == 12'h303 ? mret_legal : _GEN_95; // @[CSR.scala 388:39 393:15]
  wire  _GEN_113 = io_rw_addr == 12'h304 ? mret_legal : _GEN_99; // @[CSR.scala 434:35 444:15]
  wire  _GEN_121 = io_rw_addr == 12'h104 ? prv_is_ms : _GEN_113; // @[CSR.scala 446:35 453:15]
  wire  _GEN_125 = io_rw_addr == 12'h305 ? mret_legal : _GEN_121; // @[CSR.scala 463:37 468:15]
  wire  _GEN_129 = io_rw_addr == 12'h306 ? mret_legal : _GEN_125; // @[CSR.scala 478:42 483:15]
  wire  _GEN_133 = io_rw_addr == 12'h340 ? mret_legal : _GEN_129; // @[CSR.scala 493:40 498:15]
  wire  _GEN_137 = io_rw_addr == 12'h341 ? mret_legal : _GEN_133; // @[CSR.scala 508:36 513:15]
  wire  _GEN_141 = io_rw_addr == 12'h342 ? mret_legal : _GEN_137; // @[CSR.scala 523:38 528:15]
  wire  _GEN_145 = io_rw_addr == 12'h343 ? mret_legal : _GEN_141; // @[CSR.scala 538:37 543:15]
  wire  _GEN_153 = io_rw_addr == 12'h344 ? mret_legal : _GEN_145; // @[CSR.scala 585:35 592:15]
  wire  _GEN_157 = io_rw_addr == 12'h144 ? prv_is_ms : _GEN_153; // @[CSR.scala 594:35 599:15]
  wire  _GEN_161 = io_rw_addr == 12'hb00 ? mret_legal : _GEN_157; // @[CSR.scala 610:38 615:15]
  wire  _GEN_163 = io_rw_addr == 12'hc00 ? mret_legal | prv_is_s & mcounteren[0] | prv_is_u & mcounteren[0] & scounteren
    [0] : _GEN_161; // @[CSR.scala 617:37 619:15]
  wire  _GEN_167 = io_rw_addr == 12'hb02 ? mret_legal : _GEN_163; // @[CSR.scala 632:40 637:15]
  wire  csr_legal = io_rw_addr == 12'hc02 ? mret_legal | prv_is_s & mcounteren[2] | prv_is_u & mcounteren[2] &
    scounteren[2] : _GEN_167; // @[CSR.scala 639:39 641:15]
  wire  wen = io_rw_cmd != 2'h0 & io_uop_exc == 3'h0 & csr_legal; // @[CSR.scala 58:81]
  reg [63:0] instret; // @[CSR.scala 630:24]
  reg [63:0] cycle; // @[CSR.scala 608:22]
  reg  ip_seip_r; // @[CSR.scala 558:26]
  wire  ip_seip = io_interrupt_seip | ip_seip_r; // @[CSR.scala 559:38]
  reg  ip_stip; // @[CSR.scala 556:26]
  reg  ip_ssip; // @[CSR.scala 554:26]
  wire [63:0] sip = {54'h0,ip_seip,3'h0,ip_stip,3'h0,ip_ssip,1'h0}; // @[Cat.scala 33:92]
  wire [5:0] mip_lo = {ip_stip,1'h0,io_interrupt_msip,1'h0,ip_ssip,1'h0}; // @[Cat.scala 33:92]
  wire [63:0] mip = {52'h0,io_interrupt_meip,1'h0,ip_seip,1'h0,io_interrupt_mtip,1'h0,mip_lo}; // @[Cat.scala 33:92]
  reg [63:0] mtval; // @[CSR.scala 537:22]
  reg [63:0] mcause; // @[CSR.scala 522:23]
  reg [63:0] mepc; // @[CSR.scala 507:21]
  reg [63:0] mscratch; // @[CSR.scala 492:25]
  reg [63:0] mtvec; // @[CSR.scala 462:22]
  reg  ie_seie; // @[CSR.scala 408:24]
  reg  ie_stie; // @[CSR.scala 406:24]
  reg  ie_ssie; // @[CSR.scala 404:24]
  wire [63:0] sie = {54'h0,ie_seie,3'h0,ie_stie,3'h0,ie_ssie,1'h0}; // @[Cat.scala 33:92]
  reg  ie_meie; // @[CSR.scala 409:24]
  reg  ie_mtie; // @[CSR.scala 407:24]
  reg  ie_msie; // @[CSR.scala 405:24]
  wire [5:0] mie_lo = {ie_stie,1'h0,ie_msie,1'h0,ie_ssie,1'h0}; // @[Cat.scala 33:92]
  wire [63:0] mie = {52'h0,ie_meie,1'h0,ie_seie,1'h0,ie_mtie,1'h0,mie_lo}; // @[Cat.scala 33:92]
  reg [63:0] mideleg; // @[CSR.scala 387:24]
  reg [63:0] medeleg; // @[CSR.scala 372:24]
  reg [63:0] mhartid; // @[CSR.scala 342:33]
  reg [63:0] satp; // @[CSR.scala 283:29]
  reg [63:0] stval; // @[CSR.scala 268:22]
  reg [63:0] scause; // @[CSR.scala 253:23]
  reg [63:0] sepc; // @[CSR.scala 238:21]
  reg [63:0] sscratch; // @[CSR.scala 223:25]
  reg [63:0] stvec; // @[CSR.scala 193:22]
  reg [1:0] status_fs; // @[CSR.scala 86:28]
  wire  status_sd = |status_fs; // @[CSR.scala 91:31]
  reg  mstatus_tsr; // @[CSR.scala 119:29]
  reg  mstatus_tw; // @[CSR.scala 118:29]
  reg  status_mxr; // @[CSR.scala 89:28]
  reg  status_sum; // @[CSR.scala 88:28]
  reg  mstatus_mprv; // @[CSR.scala 116:29]
  wire [46:0] mstatus_hi = {status_sd,25'h0,2'h0,13'h1400,mstatus_tsr,mstatus_tw,mstatus_tvm,status_mxr,status_sum,
    mstatus_mprv}; // @[Cat.scala 33:92]
  reg [1:0] mstatus_mpp; // @[CSR.scala 115:29]
  reg  status_spp; // @[CSR.scala 84:28]
  reg  mstatus_mpie; // @[CSR.scala 114:29]
  reg  status_spie; // @[CSR.scala 82:28]
  reg  mstatus_mie; // @[CSR.scala 113:29]
  reg  status_sie; // @[CSR.scala 81:28]
  wire [5:0] mstatus_lo_lo = {status_spie,1'h0,mstatus_mie,1'h0,status_sie,1'h0}; // @[Cat.scala 33:92]
  wire [63:0] mstatus = {mstatus_hi,2'h0,status_fs,mstatus_mpp,2'h0,status_spp,mstatus_mpie,1'h0,mstatus_lo_lo}; // @[Cat.scala 33:92]
  wire [12:0] sstatus_lo = {4'h0,status_spp,2'h0,status_spie,3'h0,status_sie,1'h0}; // @[Cat.scala 33:92]
  wire [63:0] sstatus = {status_sd,29'h0,2'h2,12'h0,status_mxr,status_sum,1'h0,2'h0,status_fs,sstatus_lo}; // @[Cat.scala 33:92]
  wire [63:0] _GEN_6 = io_rw_addr == 12'h100 ? sstatus : 64'h0; // @[CSR.scala 151:39 152:11 56:30]
  wire [63:0] _GEN_27 = io_rw_addr == 12'h300 ? mstatus : _GEN_6; // @[CSR.scala 164:39 165:11]
  wire [63:0] _GEN_43 = io_rw_addr == 12'h105 ? stvec : _GEN_27; // @[CSR.scala 194:37 195:11]
  wire [63:0] _GEN_47 = io_rw_addr == 12'h106 ? scounteren : _GEN_43; // @[CSR.scala 209:42 210:11]
  wire [63:0] _GEN_51 = io_rw_addr == 12'h140 ? sscratch : _GEN_47; // @[CSR.scala 224:40 225:11]
  wire [63:0] _GEN_55 = io_rw_addr == 12'h141 ? sepc : _GEN_51; // @[CSR.scala 239:36 240:11]
  wire [63:0] _GEN_59 = io_rw_addr == 12'h142 ? scause : _GEN_55; // @[CSR.scala 254:38 255:11]
  wire [63:0] _GEN_63 = io_rw_addr == 12'h143 ? stval : _GEN_59; // @[CSR.scala 269:37 270:11]
  wire [63:0] _GEN_71 = io_rw_addr == 12'h180 ? satp : _GEN_63; // @[CSR.scala 291:36 292:11]
  wire [63:0] _GEN_78 = io_rw_addr == 12'hf11 ? 64'h0 : _GEN_71; // @[CSR.scala 309:41 310:15]
  wire [63:0] _GEN_80 = io_rw_addr == 12'hf12 ? 64'h0 : _GEN_78; // @[CSR.scala 320:39 321:15]
  wire [63:0] _GEN_82 = io_rw_addr == 12'hf13 ? 64'h0 : _GEN_80; // @[CSR.scala 331:38 332:15]
  wire [63:0] _GEN_86 = io_rw_addr == 12'hf14 ? mhartid : _GEN_82; // @[CSR.scala 344:39 345:11]
  wire [63:0] _GEN_90 = io_rw_addr == 12'h301 ? 64'h8000000000141101 : _GEN_86; // @[CSR.scala 361:36 362:15]
  wire [63:0] _GEN_93 = io_rw_addr == 12'h302 ? medeleg : _GEN_90; // @[CSR.scala 373:39 374:11]
  wire [63:0] _GEN_97 = io_rw_addr == 12'h303 ? mideleg : _GEN_93; // @[CSR.scala 388:39 389:11]
  wire [63:0] _GEN_106 = io_rw_addr == 12'h304 ? mie : _GEN_97; // @[CSR.scala 434:35 435:11]
  wire [63:0] _GEN_117 = io_rw_addr == 12'h104 ? sie : _GEN_106; // @[CSR.scala 446:35 447:11]
  wire [63:0] _GEN_123 = io_rw_addr == 12'h305 ? mtvec : _GEN_117; // @[CSR.scala 463:37 464:11]
  wire [63:0] _GEN_127 = io_rw_addr == 12'h306 ? mcounteren : _GEN_123; // @[CSR.scala 478:42 479:11]
  wire [63:0] _GEN_131 = io_rw_addr == 12'h340 ? mscratch : _GEN_127; // @[CSR.scala 493:40 494:11]
  wire [63:0] _GEN_135 = io_rw_addr == 12'h341 ? mepc : _GEN_131; // @[CSR.scala 508:36 509:11]
  wire [63:0] _GEN_139 = io_rw_addr == 12'h342 ? mcause : _GEN_135; // @[CSR.scala 523:38 524:11]
  wire [63:0] _GEN_143 = io_rw_addr == 12'h343 ? mtval : _GEN_139; // @[CSR.scala 538:37 539:11]
  wire [63:0] _GEN_149 = io_rw_addr == 12'h344 ? mip : _GEN_143; // @[CSR.scala 585:35 586:11]
  wire [63:0] _GEN_155 = io_rw_addr == 12'h144 ? sip : _GEN_149; // @[CSR.scala 594:35 595:11]
  wire [63:0] _GEN_159 = io_rw_addr == 12'hb00 ? cycle : _GEN_155; // @[CSR.scala 610:38 611:11]
  wire [63:0] _GEN_162 = io_rw_addr == 12'hc00 ? cycle : _GEN_159; // @[CSR.scala 617:37 618:15]
  wire [63:0] _GEN_165 = io_rw_addr == 12'hb02 ? instret : _GEN_162; // @[CSR.scala 632:40 633:11]
  wire [63:0] rdata = io_rw_addr == 12'hc02 ? instret : _GEN_165; // @[CSR.scala 639:39 640:15]
  wire [63:0] _wdata_T = rdata | io_rw_wdata; // @[CSR.scala 64:31]
  wire [63:0] _wdata_T_1 = ~io_rw_wdata; // @[CSR.scala 65:33]
  wire [63:0] _wdata_T_2 = rdata & _wdata_T_1; // @[CSR.scala 65:31]
  wire [63:0] _wdata_T_4 = 2'h1 == io_rw_cmd ? io_rw_wdata : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _wdata_T_6 = 2'h2 == io_rw_cmd ? _wdata_T : _wdata_T_4; // @[Mux.scala 81:58]
  wire [63:0] wdata = 2'h3 == io_rw_cmd ? _wdata_T_2 : _wdata_T_6; // @[Mux.scala 81:58]
  wire  _GEN_0 = wen ? wdata[1] : status_sie; // @[CSR.scala 153:15 154:19 81:28]
  wire  _GEN_1 = wen ? wdata[5] : status_spie; // @[CSR.scala 153:15 155:19 82:28]
  wire  _GEN_2 = wen ? wdata[8] : status_spp; // @[CSR.scala 153:15 156:19 84:28]
  wire [1:0] _GEN_3 = wen ? wdata[14:13] : status_fs; // @[CSR.scala 153:15 157:19 86:28]
  wire  _GEN_4 = wen ? wdata[18] : status_sum; // @[CSR.scala 153:15 159:18 88:28]
  wire  _GEN_5 = wen ? wdata[19] : status_mxr; // @[CSR.scala 153:15 160:18 89:28]
  wire  _GEN_7 = io_rw_addr == 12'h100 ? _GEN_0 : status_sie; // @[CSR.scala 151:39 81:28]
  wire  _GEN_8 = io_rw_addr == 12'h100 ? _GEN_1 : status_spie; // @[CSR.scala 151:39 82:28]
  wire  _GEN_9 = io_rw_addr == 12'h100 ? _GEN_2 : status_spp; // @[CSR.scala 151:39 84:28]
  wire [1:0] _GEN_10 = io_rw_addr == 12'h100 ? _GEN_3 : status_fs; // @[CSR.scala 151:39 86:28]
  wire  _GEN_11 = io_rw_addr == 12'h100 ? _GEN_4 : status_sum; // @[CSR.scala 151:39 88:28]
  wire  _GEN_12 = io_rw_addr == 12'h100 ? _GEN_5 : status_mxr; // @[CSR.scala 151:39 89:28]
  wire  _GEN_14 = wen ? wdata[1] : _GEN_7; // @[CSR.scala 166:15 167:19]
  wire  _GEN_15 = wen ? wdata[5] : _GEN_8; // @[CSR.scala 166:15 168:19]
  wire  _GEN_16 = wen ? wdata[8] : _GEN_9; // @[CSR.scala 166:15 169:19]
  wire  _GEN_20 = wen ? wdata[3] : mstatus_mie; // @[CSR.scala 166:15 174:20 113:29]
  wire  _GEN_21 = wen ? wdata[7] : mstatus_mpie; // @[CSR.scala 166:15 175:20 114:29]
  wire [1:0] _GEN_22 = wen ? wdata[12:11] : mstatus_mpp; // @[CSR.scala 166:15 176:20 115:29]
  wire  _GEN_23 = wen ? wdata[17] : mstatus_mprv; // @[CSR.scala 166:15 177:20 116:29]
  wire  _GEN_29 = io_rw_addr == 12'h300 ? _GEN_15 : _GEN_8; // @[CSR.scala 164:39]
  wire  _GEN_30 = io_rw_addr == 12'h300 ? _GEN_16 : _GEN_9; // @[CSR.scala 164:39]
  wire  _GEN_35 = io_rw_addr == 12'h300 ? _GEN_21 : mstatus_mpie; // @[CSR.scala 114:29 164:39]
  wire  _GEN_37 = io_rw_addr == 12'h300 ? _GEN_23 : mstatus_mprv; // @[CSR.scala 116:29 164:39]
  wire  satp_wen = wdata[62:60] == 3'h0; // @[CSR.scala 287:33]
  wire  _GEN_67 = wen & satp_wen ? wdata[63] : satp[63]; // @[CSR.scala 288:16 293:27 295:20]
  wire [15:0] _GEN_68 = wen & satp_wen ? wdata[59:44] : satp[59:44]; // @[CSR.scala 289:16 293:27 296:20]
  wire [43:0] _GEN_69 = wen & satp_wen ? wdata[43:0] : satp[43:0]; // @[CSR.scala 290:16 293:27 297:20]
  wire  _GEN_70 = wen & satp_wen & prv_is_s; // @[CSR.scala 293:27 298:20 284:33]
  wire  satp_updated = io_rw_addr == 12'h180 & _GEN_70; // @[CSR.scala 284:33 291:36]
  reg  mhartid_writable; // @[CSR.scala 343:33]
  wire  _GEN_85 = wen & mhartid_writable ? 1'h0 : mhartid_writable; // @[CSR.scala 346:35 348:24 343:33]
  wire  _GEN_88 = io_rw_addr == 12'hf14 ? _GEN_85 : mhartid_writable; // @[CSR.scala 343:33 344:39]
  wire [63:0] _medeleg_T = wdata & 64'hf7ff; // @[CSR.scala 376:24]
  wire [63:0] _mideleg_T = wdata & 64'h222; // @[CSR.scala 391:24]
  wire  _GEN_100 = wen ? wdata[1] : ie_ssie; // @[CSR.scala 436:15 437:15 404:24]
  wire  _GEN_102 = wen ? wdata[5] : ie_stie; // @[CSR.scala 436:15 439:15 406:24]
  wire  _GEN_104 = wen ? wdata[9] : ie_seie; // @[CSR.scala 436:15 441:15 408:24]
  wire  _GEN_107 = io_rw_addr == 12'h304 ? _GEN_100 : ie_ssie; // @[CSR.scala 404:24 434:35]
  wire  _GEN_109 = io_rw_addr == 12'h304 ? _GEN_102 : ie_stie; // @[CSR.scala 406:24 434:35]
  wire  _GEN_111 = io_rw_addr == 12'h304 ? _GEN_104 : ie_seie; // @[CSR.scala 408:24 434:35]
  wire  _GEN_146 = wen ? wdata[1] : ip_ssip; // @[CSR.scala 587:15 588:17 554:26]
  wire  _GEN_150 = io_rw_addr == 12'h344 ? _GEN_146 : ip_ssip; // @[CSR.scala 554:26 585:35]
  wire [63:0] _cycle_T_1 = cycle + 64'h1; // @[CSR.scala 609:18]
  wire [63:0] _GEN_218 = {{63'd0}, io_commit}; // @[CSR.scala 631:22]
  wire [63:0] _instret_T_1 = instret + _GEN_218; // @[CSR.scala 631:22]
  wire  is_mret = io_uop_sys_op == 3'h1; // @[CSR.scala 656:34]
  wire  _T_32 = is_mret & mret_legal; // @[CSR.scala 658:16]
  wire  _GEN_170 = mstatus_mpp != 2'h3 ? 1'h0 : _GEN_37; // @[CSR.scala 664:35 665:20]
  wire [1:0] _GEN_171 = is_mret & mret_legal ? mstatus_mpp : prv; // @[CSR.scala 658:31 659:18 49:26]
  wire  _GEN_173 = is_mret & mret_legal | _GEN_35; // @[CSR.scala 658:31 662:18]
  wire  _GEN_175 = is_mret & mret_legal ? _GEN_170 : _GEN_37; // @[CSR.scala 658:31]
  wire  is_sret = io_uop_sys_op == 3'h2; // @[CSR.scala 669:34]
  wire  sret_legal = prv_is_ms & ~mstatus_tsr; // @[CSR.scala 670:30]
  wire  _T_34 = is_sret & sret_legal; // @[CSR.scala 671:16]
  wire [1:0] _GEN_219 = {{1'd0}, status_spp}; // @[CSR.scala 677:21]
  wire [1:0] _GEN_177 = is_sret & sret_legal ? {{1'd0}, status_spp} : _GEN_171; // @[CSR.scala 671:31 672:17]
  wire  _GEN_179 = is_sret & sret_legal | _GEN_29; // @[CSR.scala 671:31 675:17]
  wire  _GEN_180 = is_sret & sret_legal ? 1'h0 : _GEN_30; // @[CSR.scala 671:31 676:17]
  wire  is_sfv = io_uop_sys_op == 3'h6 & io_uop_valid; // @[CSR.scala 685:55]
  wire  is_fence_i = io_uop_sys_op == 3'h5 & io_uop_valid; // @[CSR.scala 687:58]
  wire  is_sys = io_sfence_vma | is_fence_i; // @[CSR.scala 688:34]
  wire  is_exc_from_prev = io_uop_exc != 3'h0; // @[CSR.scala 695:38]
  wire  is_exc_from_lsu = io_lsu_exc_code != 4'h0; // @[CSR.scala 696:43]
  wire  is_exc_from_csr = ~csr_legal & _wen_T; // @[CSR.scala 697:37]
  wire  _is_exc_from_sys_T = ~mret_legal; // @[CSR.scala 698:38]
  wire  is_exc_from_sys = is_mret & ~mret_legal | is_sret & ~sret_legal | is_sfv & ~_csr_legal_T_1; // @[CSR.scala 698:79]
  wire  is_exc = is_exc_from_prev | is_exc_from_lsu | is_exc_from_csr; // @[CSR.scala 699:62]
  wire  int_attach = io_uop_valid & (io_uop_fu == 3'h0 | io_uop_fu == 3'h1); // @[CSR.scala 719:37]
  wire [63:0] int_bits = mip & mie; // @[CSR.scala 720:28]
  wire [63:0] _int_bits_mmode_T = ~mideleg; // @[CSR.scala 721:36]
  wire [63:0] int_bits_mmode = int_bits & _int_bits_mmode_T; // @[CSR.scala 721:33]
  wire [3:0] _GEN_182 = int_bits[5] ? 4'h5 : 4'h0; // @[CSR.scala 713:22 702:24 714:9]
  wire [3:0] _GEN_183 = int_bits[1] ? 4'h1 : _GEN_182; // @[CSR.scala 711:22 712:9]
  wire [3:0] _GEN_184 = int_bits[9] ? 4'h9 : _GEN_183; // @[CSR.scala 709:22 710:9]
  wire [3:0] _GEN_185 = int_bits[7] ? 4'h7 : _GEN_184; // @[CSR.scala 707:22 708:9]
  wire [3:0] _GEN_186 = int_bits[3] ? 4'h3 : _GEN_185; // @[CSR.scala 705:22 706:9]
  wire [3:0] int_index_tmp = int_bits[11] ? 4'hb : _GEN_186; // @[CSR.scala 703:17 704:9]
  wire [3:0] _GEN_188 = int_bits_mmode[5] ? 4'h5 : 4'h0; // @[CSR.scala 713:22 702:24 714:9]
  wire [3:0] _GEN_189 = int_bits_mmode[1] ? 4'h1 : _GEN_188; // @[CSR.scala 711:22 712:9]
  wire [3:0] _GEN_190 = int_bits_mmode[9] ? 4'h9 : _GEN_189; // @[CSR.scala 709:22 710:9]
  wire [3:0] _GEN_191 = int_bits_mmode[7] ? 4'h7 : _GEN_190; // @[CSR.scala 707:22 708:9]
  wire [3:0] _GEN_192 = int_bits_mmode[3] ? 4'h3 : _GEN_191; // @[CSR.scala 705:22 706:9]
  wire [3:0] int_index_y = int_bits_mmode[11] ? 4'hb : _GEN_192; // @[CSR.scala 703:17 704:9]
  wire [3:0] _GEN_194 = mstatus_mie ? int_index_y : 4'h0; // @[CSR.scala 726:30 727:17 723:34]
  wire [15:0] _T_38 = 16'h1 << int_index_tmp; // @[CSR.scala 730:16]
  wire [63:0] _GEN_220 = {{48'd0}, _T_38}; // @[CSR.scala 730:34]
  wire [63:0] _T_39 = _GEN_220 & mideleg; // @[CSR.scala 730:34]
  wire [3:0] _GEN_195 = status_sie | prv_is_u ? int_index_tmp : 4'h0; // @[CSR.scala 731:50 732:19 723:34]
  wire [3:0] _GEN_196 = mstatus_mie | prv_is_u | prv_is_s ? int_index_tmp : 4'h0; // @[CSR.scala 735:70 736:19 723:34]
  wire [3:0] _GEN_197 = _T_39 != 64'h0 ? _GEN_195 : _GEN_196; // @[CSR.scala 730:54]
  wire [3:0] int_index = mret_legal ? _GEN_194 : _GEN_197; // @[CSR.scala 725:25]
  wire  is_int = int_attach & int_index != 4'h0; // @[CSR.scala 740:27]
  wire [1:0] _cause_exc_T_2 = is_exc_from_csr | is_exc_from_sys ? 2'h2 : 2'h0; // @[CSR.scala 751:10]
  wire [3:0] _cause_exc_T_3 = is_exc_from_lsu ? io_lsu_exc_code : {{2'd0}, _cause_exc_T_2}; // @[CSR.scala 748:8]
  wire [3:0] _cause_exc_T_4 = {2'h2,prv}; // @[Cat.scala 33:92]
  wire [3:0] _cause_exc_T_6 = 3'h1 == io_uop_exc ? 4'h0 : _cause_exc_T_3; // @[Mux.scala 81:58]
  wire [3:0] _cause_exc_T_8 = 3'h2 == io_uop_exc ? 4'h1 : _cause_exc_T_6; // @[Mux.scala 81:58]
  wire [3:0] _cause_exc_T_10 = 3'h4 == io_uop_exc ? 4'h2 : _cause_exc_T_8; // @[Mux.scala 81:58]
  wire [3:0] _cause_exc_T_12 = 3'h7 == io_uop_exc ? 4'h3 : _cause_exc_T_10; // @[Mux.scala 81:58]
  wire [3:0] _cause_exc_T_14 = 3'h5 == io_uop_exc ? _cause_exc_T_4 : _cause_exc_T_12; // @[Mux.scala 81:58]
  wire [3:0] cause_exc = 3'h3 == io_uop_exc ? 4'hc : _cause_exc_T_14; // @[Mux.scala 81:58]
  wire [15:0] cause_exc_onehot = 16'h1 << cause_exc; // @[OneHot.scala 57:35]
  wire [15:0] cause_int_onehot = 16'h1 << int_index; // @[OneHot.scala 57:35]
  wire  trap = is_exc | is_int; // @[CSR.scala 796:26]
  wire [63:0] _GEN_221 = {{48'd0}, cause_exc_onehot}; // @[CSR.scala 801:37]
  wire [63:0] _trap_to_s_T = _GEN_221 & medeleg; // @[CSR.scala 801:37]
  wire [63:0] _GEN_222 = {{48'd0}, cause_int_onehot}; // @[CSR.scala 802:37]
  wire [63:0] _trap_to_s_T_3 = _GEN_222 & mideleg; // @[CSR.scala 802:37]
  wire  _trap_to_s_T_5 = is_int & _trap_to_s_T_3 != 64'h0; // @[CSR.scala 802:15]
  wire  _trap_to_s_T_6 = is_exc & _trap_to_s_T != 64'h0 | _trap_to_s_T_5; // @[CSR.scala 801:58]
  wire  trap_to_s = _is_exc_from_sys_T & _trap_to_s_T_6; // @[CSR.scala 799:19 800:15 797:30]
  wire [63:0] _scause_T = {60'h800000000000000,int_index}; // @[Cat.scala 33:92]
  wire [3:0] _trap_pc_T_4 = is_int & stvec[1:0] == 2'h1 ? int_index : 4'h0; // @[CSR.scala 813:48]
  wire [61:0] _GEN_223 = {{58'd0}, _trap_pc_T_4}; // @[CSR.scala 813:43]
  wire [61:0] _trap_pc_T_6 = stvec[63:2] + _GEN_223; // @[CSR.scala 813:43]
  wire [63:0] _trap_pc_T_7 = {_trap_pc_T_6,2'h0}; // @[Cat.scala 33:92]
  wire [1:0] _GEN_207 = trap_to_s & trap ? prv : {{1'd0}, _GEN_180}; // @[CSR.scala 804:27 810:17]
  wire [1:0] _GEN_208 = trap_to_s & trap ? 2'h1 : _GEN_177; // @[CSR.scala 804:27 811:17]
  wire [63:0] _GEN_209 = trap_to_s & trap ? _trap_pc_T_7 : 64'h0; // @[CSR.scala 804:27 813:17 798:30]
  wire [3:0] _trap_pc_T_12 = is_int & mtvec[1:0] == 2'h1 ? int_index : 4'h0; // @[CSR.scala 824:49]
  wire [61:0] _GEN_224 = {{58'd0}, _trap_pc_T_12}; // @[CSR.scala 824:44]
  wire [61:0] _trap_pc_T_14 = mtvec[63:2] + _GEN_224; // @[CSR.scala 824:44]
  wire [63:0] _trap_pc_T_15 = {_trap_pc_T_14,2'h0}; // @[Cat.scala 33:92]
  wire [63:0] trap_pc = ~trap_to_s & trap ? _trap_pc_T_15 : _GEN_209; // @[CSR.scala 815:28 824:18]
  wire [63:0] _io_jmp_packet_target_T_1 = is_mret ? mepc : sepc; // @[CSR.scala 830:89]
  wire [63:0] _io_jmp_packet_target_T_2 = is_sys | satp_updated ? io_uop_npc : _io_jmp_packet_target_T_1; // @[CSR.scala 830:49]
  wire [1:0] _GEN_225 = reset ? 2'h0 : _GEN_207; // @[CSR.scala 84:{28,28}]
  assign io_rw_rdata = io_rw_addr == 12'hc02 ? instret : _GEN_165; // @[CSR.scala 639:39 640:15]
  assign io_rw_valid = io_rw_addr == 12'hc02 ? mret_legal | prv_is_s & mcounteren[2] | prv_is_u & mcounteren[2] &
    scounteren[2] : _GEN_167; // @[CSR.scala 639:39 641:15]
  assign io_prv = ~trap_to_s & trap ? 2'h3 : _GEN_208; // @[CSR.scala 815:28 822:18]
  assign io_mprv = mstatus_mprv; // @[CSR.scala 184:11]
  assign io_mpp = mstatus_mpp; // @[CSR.scala 185:11]
  assign io_sv39_en = io_rw_addr == 12'h180 ? _GEN_67 : satp[63]; // @[CSR.scala 288:16 291:36]
  assign io_satp_asid = io_rw_addr == 12'h180 ? _GEN_68 : satp[59:44]; // @[CSR.scala 289:16 291:36]
  assign io_satp_ppn = io_rw_addr == 12'h180 ? _GEN_69 : satp[43:0]; // @[CSR.scala 290:16 291:36]
  assign io_sfence_vma = is_sfv & _csr_legal_T_1; // @[CSR.scala 689:27]
  assign io_fence_i = io_uop_sys_op == 3'h5 & io_uop_valid; // @[CSR.scala 687:58]
  assign io_jmp_packet_valid = trap | is_sys | satp_updated | _T_32 | _T_34; // @[CSR.scala 829:85]
  assign io_jmp_packet_target = trap ? trap_pc : _io_jmp_packet_target_T_2; // @[CSR.scala 830:30]
  assign io_is_int = int_attach & int_index != 4'h0; // @[CSR.scala 740:27]
  always @(posedge clock) begin
    if (reset) begin // @[CSR.scala 49:26]
      prv <= 2'h3; // @[CSR.scala 49:26]
    end else if (~trap_to_s & trap) begin // @[CSR.scala 815:28]
      prv <= 2'h3; // @[CSR.scala 822:18]
    end else if (trap_to_s & trap) begin // @[CSR.scala 804:27]
      prv <= 2'h1; // @[CSR.scala 811:17]
    end else if (is_sret & sret_legal) begin // @[CSR.scala 671:31]
      prv <= {{1'd0}, status_spp}; // @[CSR.scala 672:17]
    end else begin
      prv <= _GEN_171;
    end
    if (reset) begin // @[CSR.scala 477:27]
      mcounteren <= 64'h0; // @[CSR.scala 477:27]
    end else if (io_rw_addr == 12'h306) begin // @[CSR.scala 478:42]
      if (wen) begin // @[CSR.scala 480:15]
        if (2'h3 == io_rw_cmd) begin // @[Mux.scala 81:58]
          mcounteren <= _wdata_T_2;
        end else begin
          mcounteren <= _wdata_T_6;
        end
      end
    end
    if (reset) begin // @[CSR.scala 208:27]
      scounteren <= 64'h0; // @[CSR.scala 208:27]
    end else if (io_rw_addr == 12'h106) begin // @[CSR.scala 209:42]
      if (wen) begin // @[CSR.scala 211:15]
        if (2'h3 == io_rw_cmd) begin // @[Mux.scala 81:58]
          scounteren <= _wdata_T_2;
        end else begin
          scounteren <= _wdata_T_6;
        end
      end
    end
    if (reset) begin // @[CSR.scala 117:29]
      mstatus_tvm <= 1'h0; // @[CSR.scala 117:29]
    end else if (io_rw_addr == 12'h300) begin // @[CSR.scala 164:39]
      if (wen) begin // @[CSR.scala 166:15]
        mstatus_tvm <= wdata[20]; // @[CSR.scala 178:20]
      end
    end
    if (reset) begin // @[CSR.scala 630:24]
      instret <= 64'h0; // @[CSR.scala 630:24]
    end else if (io_rw_addr == 12'hb02) begin // @[CSR.scala 632:40]
      if (wen) begin // @[CSR.scala 634:15]
        if (2'h3 == io_rw_cmd) begin // @[Mux.scala 81:58]
          instret <= _wdata_T_2;
        end else begin
          instret <= _wdata_T_6;
        end
      end else begin
        instret <= _instret_T_1; // @[CSR.scala 631:11]
      end
    end else begin
      instret <= _instret_T_1; // @[CSR.scala 631:11]
    end
    if (reset) begin // @[CSR.scala 608:22]
      cycle <= 64'h0; // @[CSR.scala 608:22]
    end else if (io_rw_addr == 12'hb00) begin // @[CSR.scala 610:38]
      if (wen) begin // @[CSR.scala 612:15]
        if (2'h3 == io_rw_cmd) begin // @[Mux.scala 81:58]
          cycle <= _wdata_T_2;
        end else begin
          cycle <= _wdata_T_6;
        end
      end else begin
        cycle <= _cycle_T_1; // @[CSR.scala 609:9]
      end
    end else begin
      cycle <= _cycle_T_1; // @[CSR.scala 609:9]
    end
    if (reset) begin // @[CSR.scala 558:26]
      ip_seip_r <= 1'h0; // @[CSR.scala 558:26]
    end else if (io_rw_addr == 12'h344) begin // @[CSR.scala 585:35]
      if (wen) begin // @[CSR.scala 587:15]
        ip_seip_r <= wdata[9]; // @[CSR.scala 590:17]
      end
    end
    if (reset) begin // @[CSR.scala 556:26]
      ip_stip <= 1'h0; // @[CSR.scala 556:26]
    end else if (io_rw_addr == 12'h344) begin // @[CSR.scala 585:35]
      if (wen) begin // @[CSR.scala 587:15]
        ip_stip <= wdata[5]; // @[CSR.scala 589:17]
      end
    end
    if (reset) begin // @[CSR.scala 554:26]
      ip_ssip <= 1'h0; // @[CSR.scala 554:26]
    end else if (io_rw_addr == 12'h144) begin // @[CSR.scala 594:35]
      if (wen) begin // @[CSR.scala 596:15]
        ip_ssip <= wdata[1]; // @[CSR.scala 597:15]
      end else begin
        ip_ssip <= _GEN_150;
      end
    end else begin
      ip_ssip <= _GEN_150;
    end
    if (reset) begin // @[CSR.scala 537:22]
      mtval <= 64'h0; // @[CSR.scala 537:22]
    end else if (~trap_to_s & trap) begin // @[CSR.scala 815:28]
      if (io_uop_exc == 3'h3) begin // @[CSR.scala 792:39]
        mtval <= io_uop_pc; // @[CSR.scala 793:10]
      end else if (is_exc_from_lsu) begin // @[CSR.scala 789:25]
        mtval <= io_lsu_addr; // @[CSR.scala 790:10]
      end else begin
        mtval <= 64'h0; // @[CSR.scala 788:25]
      end
    end else if (io_rw_addr == 12'h343) begin // @[CSR.scala 538:37]
      if (wen) begin // @[CSR.scala 540:15]
        mtval <= wdata; // @[CSR.scala 541:13]
      end
    end
    if (reset) begin // @[CSR.scala 522:23]
      mcause <= 64'h0; // @[CSR.scala 522:23]
    end else if (~trap_to_s & trap) begin // @[CSR.scala 815:28]
      if (is_exc) begin // @[CSR.scala 806:23]
        mcause <= {{60'd0}, cause_exc};
      end else begin
        mcause <= _scause_T;
      end
    end else if (io_rw_addr == 12'h342) begin // @[CSR.scala 523:38]
      if (wen) begin // @[CSR.scala 525:15]
        mcause <= wdata; // @[CSR.scala 526:14]
      end
    end
    if (reset) begin // @[CSR.scala 507:21]
      mepc <= 64'h0; // @[CSR.scala 507:21]
    end else if (~trap_to_s & trap) begin // @[CSR.scala 815:28]
      mepc <= io_uop_pc; // @[CSR.scala 818:18]
    end else if (io_rw_addr == 12'h341) begin // @[CSR.scala 508:36]
      if (wen) begin // @[CSR.scala 510:15]
        mepc <= wdata; // @[CSR.scala 511:12]
      end
    end
    if (reset) begin // @[CSR.scala 492:25]
      mscratch <= 64'h0; // @[CSR.scala 492:25]
    end else if (io_rw_addr == 12'h340) begin // @[CSR.scala 493:40]
      if (wen) begin // @[CSR.scala 495:15]
        if (2'h3 == io_rw_cmd) begin // @[Mux.scala 81:58]
          mscratch <= _wdata_T_2;
        end else begin
          mscratch <= _wdata_T_6;
        end
      end
    end
    if (reset) begin // @[CSR.scala 462:22]
      mtvec <= 64'h0; // @[CSR.scala 462:22]
    end else if (io_rw_addr == 12'h305) begin // @[CSR.scala 463:37]
      if (wen) begin // @[CSR.scala 465:15]
        if (2'h3 == io_rw_cmd) begin // @[Mux.scala 81:58]
          mtvec <= _wdata_T_2;
        end else begin
          mtvec <= _wdata_T_6;
        end
      end
    end
    if (reset) begin // @[CSR.scala 408:24]
      ie_seie <= 1'h0; // @[CSR.scala 408:24]
    end else if (io_rw_addr == 12'h104) begin // @[CSR.scala 446:35]
      if (wen) begin // @[CSR.scala 448:15]
        ie_seie <= wdata[9]; // @[CSR.scala 451:15]
      end else begin
        ie_seie <= _GEN_111;
      end
    end else begin
      ie_seie <= _GEN_111;
    end
    if (reset) begin // @[CSR.scala 406:24]
      ie_stie <= 1'h0; // @[CSR.scala 406:24]
    end else if (io_rw_addr == 12'h104) begin // @[CSR.scala 446:35]
      if (wen) begin // @[CSR.scala 448:15]
        ie_stie <= wdata[5]; // @[CSR.scala 450:15]
      end else begin
        ie_stie <= _GEN_109;
      end
    end else begin
      ie_stie <= _GEN_109;
    end
    if (reset) begin // @[CSR.scala 404:24]
      ie_ssie <= 1'h0; // @[CSR.scala 404:24]
    end else if (io_rw_addr == 12'h104) begin // @[CSR.scala 446:35]
      if (wen) begin // @[CSR.scala 448:15]
        ie_ssie <= wdata[1]; // @[CSR.scala 449:15]
      end else begin
        ie_ssie <= _GEN_107;
      end
    end else begin
      ie_ssie <= _GEN_107;
    end
    if (reset) begin // @[CSR.scala 409:24]
      ie_meie <= 1'h0; // @[CSR.scala 409:24]
    end else if (io_rw_addr == 12'h304) begin // @[CSR.scala 434:35]
      if (wen) begin // @[CSR.scala 436:15]
        ie_meie <= wdata[11]; // @[CSR.scala 442:15]
      end
    end
    if (reset) begin // @[CSR.scala 407:24]
      ie_mtie <= 1'h0; // @[CSR.scala 407:24]
    end else if (io_rw_addr == 12'h304) begin // @[CSR.scala 434:35]
      if (wen) begin // @[CSR.scala 436:15]
        ie_mtie <= wdata[7]; // @[CSR.scala 440:15]
      end
    end
    if (reset) begin // @[CSR.scala 405:24]
      ie_msie <= 1'h0; // @[CSR.scala 405:24]
    end else if (io_rw_addr == 12'h304) begin // @[CSR.scala 434:35]
      if (wen) begin // @[CSR.scala 436:15]
        ie_msie <= wdata[3]; // @[CSR.scala 438:15]
      end
    end
    if (reset) begin // @[CSR.scala 387:24]
      mideleg <= 64'h0; // @[CSR.scala 387:24]
    end else if (io_rw_addr == 12'h303) begin // @[CSR.scala 388:39]
      if (wen) begin // @[CSR.scala 390:15]
        mideleg <= _mideleg_T; // @[CSR.scala 391:15]
      end
    end
    if (reset) begin // @[CSR.scala 372:24]
      medeleg <= 64'h0; // @[CSR.scala 372:24]
    end else if (io_rw_addr == 12'h302) begin // @[CSR.scala 373:39]
      if (wen) begin // @[CSR.scala 375:15]
        medeleg <= _medeleg_T; // @[CSR.scala 376:15]
      end
    end
    if (reset) begin // @[CSR.scala 342:33]
      mhartid <= 64'h0; // @[CSR.scala 342:33]
    end else if (io_rw_addr == 12'hf14) begin // @[CSR.scala 344:39]
      if (wen & mhartid_writable) begin // @[CSR.scala 346:35]
        if (2'h3 == io_rw_cmd) begin // @[Mux.scala 81:58]
          mhartid <= _wdata_T_2;
        end else begin
          mhartid <= _wdata_T_6;
        end
      end
    end
    if (reset) begin // @[CSR.scala 283:29]
      satp <= 64'h0; // @[CSR.scala 283:29]
    end else if (io_rw_addr == 12'h180) begin // @[CSR.scala 291:36]
      if (wen & satp_wen) begin // @[CSR.scala 293:27]
        if (2'h3 == io_rw_cmd) begin // @[Mux.scala 81:58]
          satp <= _wdata_T_2;
        end else begin
          satp <= _wdata_T_6;
        end
      end
    end
    if (reset) begin // @[CSR.scala 268:22]
      stval <= 64'h0; // @[CSR.scala 268:22]
    end else if (trap_to_s & trap) begin // @[CSR.scala 804:27]
      if (io_uop_exc == 3'h3) begin // @[CSR.scala 792:39]
        stval <= io_uop_pc; // @[CSR.scala 793:10]
      end else if (is_exc_from_lsu) begin // @[CSR.scala 789:25]
        stval <= io_lsu_addr; // @[CSR.scala 790:10]
      end else begin
        stval <= 64'h0; // @[CSR.scala 788:25]
      end
    end else if (io_rw_addr == 12'h143) begin // @[CSR.scala 269:37]
      if (wen) begin // @[CSR.scala 271:15]
        stval <= wdata; // @[CSR.scala 272:13]
      end
    end
    if (reset) begin // @[CSR.scala 253:23]
      scause <= 64'h0; // @[CSR.scala 253:23]
    end else if (trap_to_s & trap) begin // @[CSR.scala 804:27]
      if (is_exc) begin // @[CSR.scala 806:23]
        scause <= {{60'd0}, cause_exc};
      end else begin
        scause <= _scause_T;
      end
    end else if (io_rw_addr == 12'h142) begin // @[CSR.scala 254:38]
      if (wen) begin // @[CSR.scala 256:15]
        scause <= wdata; // @[CSR.scala 257:14]
      end
    end
    if (reset) begin // @[CSR.scala 238:21]
      sepc <= 64'h0; // @[CSR.scala 238:21]
    end else if (trap_to_s & trap) begin // @[CSR.scala 804:27]
      sepc <= io_uop_pc; // @[CSR.scala 807:17]
    end else if (io_rw_addr == 12'h141) begin // @[CSR.scala 239:36]
      if (wen) begin // @[CSR.scala 241:15]
        sepc <= wdata; // @[CSR.scala 242:12]
      end
    end
    if (reset) begin // @[CSR.scala 223:25]
      sscratch <= 64'h0; // @[CSR.scala 223:25]
    end else if (io_rw_addr == 12'h140) begin // @[CSR.scala 224:40]
      if (wen) begin // @[CSR.scala 226:15]
        if (2'h3 == io_rw_cmd) begin // @[Mux.scala 81:58]
          sscratch <= _wdata_T_2;
        end else begin
          sscratch <= _wdata_T_6;
        end
      end
    end
    if (reset) begin // @[CSR.scala 193:22]
      stvec <= 64'h0; // @[CSR.scala 193:22]
    end else if (io_rw_addr == 12'h105) begin // @[CSR.scala 194:37]
      if (wen) begin // @[CSR.scala 196:15]
        if (2'h3 == io_rw_cmd) begin // @[Mux.scala 81:58]
          stvec <= _wdata_T_2;
        end else begin
          stvec <= _wdata_T_6;
        end
      end
    end
    if (reset) begin // @[CSR.scala 86:28]
      status_fs <= 2'h0; // @[CSR.scala 86:28]
    end else if (io_rw_addr == 12'h300) begin // @[CSR.scala 164:39]
      if (wen) begin // @[CSR.scala 166:15]
        status_fs <= wdata[14:13]; // @[CSR.scala 170:19]
      end else begin
        status_fs <= _GEN_10;
      end
    end else begin
      status_fs <= _GEN_10;
    end
    if (reset) begin // @[CSR.scala 119:29]
      mstatus_tsr <= 1'h0; // @[CSR.scala 119:29]
    end else if (io_rw_addr == 12'h300) begin // @[CSR.scala 164:39]
      if (wen) begin // @[CSR.scala 166:15]
        mstatus_tsr <= wdata[22]; // @[CSR.scala 180:20]
      end
    end
    if (reset) begin // @[CSR.scala 118:29]
      mstatus_tw <= 1'h0; // @[CSR.scala 118:29]
    end else if (io_rw_addr == 12'h300) begin // @[CSR.scala 164:39]
      if (wen) begin // @[CSR.scala 166:15]
        mstatus_tw <= wdata[21]; // @[CSR.scala 179:20]
      end
    end
    if (reset) begin // @[CSR.scala 89:28]
      status_mxr <= 1'h0; // @[CSR.scala 89:28]
    end else if (io_rw_addr == 12'h300) begin // @[CSR.scala 164:39]
      if (wen) begin // @[CSR.scala 166:15]
        status_mxr <= wdata[19]; // @[CSR.scala 173:20]
      end else begin
        status_mxr <= _GEN_12;
      end
    end else begin
      status_mxr <= _GEN_12;
    end
    if (reset) begin // @[CSR.scala 88:28]
      status_sum <= 1'h0; // @[CSR.scala 88:28]
    end else if (io_rw_addr == 12'h300) begin // @[CSR.scala 164:39]
      if (wen) begin // @[CSR.scala 166:15]
        status_sum <= wdata[18]; // @[CSR.scala 172:20]
      end else begin
        status_sum <= _GEN_11;
      end
    end else begin
      status_sum <= _GEN_11;
    end
    if (reset) begin // @[CSR.scala 116:29]
      mstatus_mprv <= 1'h0; // @[CSR.scala 116:29]
    end else if (is_sret & sret_legal) begin // @[CSR.scala 671:31]
      if (_GEN_219 != 2'h3) begin // @[CSR.scala 677:34]
        mstatus_mprv <= 1'h0; // @[CSR.scala 678:20]
      end else begin
        mstatus_mprv <= _GEN_175;
      end
    end else begin
      mstatus_mprv <= _GEN_175;
    end
    if (reset) begin // @[CSR.scala 115:29]
      mstatus_mpp <= 2'h0; // @[CSR.scala 115:29]
    end else if (~trap_to_s & trap) begin // @[CSR.scala 815:28]
      mstatus_mpp <= prv; // @[CSR.scala 821:18]
    end else if (is_mret & mret_legal) begin // @[CSR.scala 658:31]
      mstatus_mpp <= 2'h0; // @[CSR.scala 663:18]
    end else if (io_rw_addr == 12'h300) begin // @[CSR.scala 164:39]
      mstatus_mpp <= _GEN_22;
    end
    status_spp <= _GEN_225[0]; // @[CSR.scala 84:{28,28}]
    if (reset) begin // @[CSR.scala 114:29]
      mstatus_mpie <= 1'h0; // @[CSR.scala 114:29]
    end else if (~trap_to_s & trap) begin // @[CSR.scala 815:28]
      mstatus_mpie <= mstatus_mie; // @[CSR.scala 819:18]
    end else begin
      mstatus_mpie <= _GEN_173;
    end
    if (reset) begin // @[CSR.scala 82:28]
      status_spie <= 1'h0; // @[CSR.scala 82:28]
    end else if (trap_to_s & trap) begin // @[CSR.scala 804:27]
      status_spie <= status_sie; // @[CSR.scala 808:17]
    end else begin
      status_spie <= _GEN_179;
    end
    if (reset) begin // @[CSR.scala 113:29]
      mstatus_mie <= 1'h0; // @[CSR.scala 113:29]
    end else if (~trap_to_s & trap) begin // @[CSR.scala 815:28]
      mstatus_mie <= 1'h0; // @[CSR.scala 820:18]
    end else if (is_mret & mret_legal) begin // @[CSR.scala 658:31]
      mstatus_mie <= mstatus_mpie; // @[CSR.scala 661:18]
    end else if (io_rw_addr == 12'h300) begin // @[CSR.scala 164:39]
      mstatus_mie <= _GEN_20;
    end
    if (reset) begin // @[CSR.scala 81:28]
      status_sie <= 1'h0; // @[CSR.scala 81:28]
    end else if (trap_to_s & trap) begin // @[CSR.scala 804:27]
      status_sie <= 1'h0; // @[CSR.scala 809:17]
    end else if (is_sret & sret_legal) begin // @[CSR.scala 671:31]
      status_sie <= status_spie; // @[CSR.scala 674:17]
    end else if (io_rw_addr == 12'h300) begin // @[CSR.scala 164:39]
      status_sie <= _GEN_14;
    end else begin
      status_sie <= _GEN_7;
    end
    mhartid_writable <= reset | _GEN_88; // @[CSR.scala 343:{33,33}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  prv = _RAND_0[1:0];
  _RAND_1 = {2{`RANDOM}};
  mcounteren = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  scounteren = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  mstatus_tvm = _RAND_3[0:0];
  _RAND_4 = {2{`RANDOM}};
  instret = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  cycle = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  ip_seip_r = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  ip_stip = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  ip_ssip = _RAND_8[0:0];
  _RAND_9 = {2{`RANDOM}};
  mtval = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  mcause = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  mepc = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  mscratch = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  mtvec = _RAND_13[63:0];
  _RAND_14 = {1{`RANDOM}};
  ie_seie = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  ie_stie = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  ie_ssie = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  ie_meie = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  ie_mtie = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  ie_msie = _RAND_19[0:0];
  _RAND_20 = {2{`RANDOM}};
  mideleg = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  medeleg = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  mhartid = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  satp = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  stval = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  scause = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  sepc = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  sscratch = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  stvec = _RAND_28[63:0];
  _RAND_29 = {1{`RANDOM}};
  status_fs = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  mstatus_tsr = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  mstatus_tw = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  status_mxr = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  status_sum = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  mstatus_mprv = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  mstatus_mpp = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  status_spp = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  mstatus_mpie = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  status_spie = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  mstatus_mie = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  status_sie = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  mhartid_writable = _RAND_41[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CachePortProxy_1(
  input         clock,
  input         reset,
  input  [1:0]  io_prv,
  input         io_sv39_en,
  input  [15:0] io_satp_asid,
  input  [43:0] io_satp_ppn,
  input         io_sfence_vma,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [38:0] io_in_req_bits_addr,
  input  [63:0] io_in_req_bits_wdata,
  input  [7:0]  io_in_req_bits_wmask,
  input         io_in_req_bits_wen,
  input  [1:0]  io_in_req_bits_len,
  input         io_in_req_bits_lrsc,
  input  [4:0]  io_in_req_bits_amo,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [63:0] io_in_resp_bits_rdata,
  output        io_in_resp_bits_page_fault,
  output        io_in_resp_bits_access_fault,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [38:0] io_out_req_bits_addr,
  output [63:0] io_out_req_bits_wdata,
  output [7:0]  io_out_req_bits_wmask,
  output        io_out_req_bits_wen,
  output [1:0]  io_out_req_bits_len,
  output        io_out_req_bits_lrsc,
  output [4:0]  io_out_req_bits_amo,
  output        io_out_resp_ready,
  input         io_out_resp_valid,
  input  [63:0] io_out_resp_bits_rdata,
  input         io_ptw_req_ready,
  output        io_ptw_req_valid,
  output [38:0] io_ptw_req_bits_addr,
  output        io_ptw_resp_ready,
  input         io_ptw_resp_valid,
  input  [63:0] io_ptw_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
`endif // RANDOMIZE_REG_INIT
  wire  tlb_clock; // @[CachePortProxy.scala 28:19]
  wire  tlb_reset; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_sfence_vma; // @[CachePortProxy.scala 28:19]
  wire [8:0] tlb_io_vaddr_vpn2; // @[CachePortProxy.scala 28:19]
  wire [8:0] tlb_io_vaddr_vpn1; // @[CachePortProxy.scala 28:19]
  wire [8:0] tlb_io_vaddr_vpn0; // @[CachePortProxy.scala 28:19]
  wire [1:0] tlb_io_rpte_ppn2; // @[CachePortProxy.scala 28:19]
  wire [8:0] tlb_io_rpte_ppn1; // @[CachePortProxy.scala 28:19]
  wire [8:0] tlb_io_rpte_ppn0; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_rpte_flag_d; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_rpte_flag_a; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_rpte_flag_u; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_rpte_flag_x; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_rpte_flag_w; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_rpte_flag_r; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_rpte_flag_v; // @[CachePortProxy.scala 28:19]
  wire [1:0] tlb_io_rlevel; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_hit; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_wen; // @[CachePortProxy.scala 28:19]
  wire [8:0] tlb_io_wvaddr_vpn2; // @[CachePortProxy.scala 28:19]
  wire [8:0] tlb_io_wvaddr_vpn1; // @[CachePortProxy.scala 28:19]
  wire [8:0] tlb_io_wvaddr_vpn0; // @[CachePortProxy.scala 28:19]
  wire [1:0] tlb_io_wpte_ppn2; // @[CachePortProxy.scala 28:19]
  wire [8:0] tlb_io_wpte_ppn1; // @[CachePortProxy.scala 28:19]
  wire [8:0] tlb_io_wpte_ppn0; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_wpte_flag_d; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_wpte_flag_a; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_wpte_flag_g; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_wpte_flag_u; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_wpte_flag_x; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_wpte_flag_w; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_wpte_flag_r; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_wpte_flag_v; // @[CachePortProxy.scala 28:19]
  wire [1:0] tlb_io_wlevel; // @[CachePortProxy.scala 28:19]
  wire [15:0] tlb_io_satp_asid; // @[CachePortProxy.scala 28:19]
  reg [2:0] state; // @[CachePortProxy.scala 21:93]
  wire  _in_req_bits_T = state == 3'h0; // @[CachePortProxy.scala 24:54]
  reg [38:0] in_req_bits_r_addr; // @[Reg.scala 35:20]
  reg [63:0] in_req_bits_r_wdata; // @[Reg.scala 35:20]
  reg [7:0] in_req_bits_r_wmask; // @[Reg.scala 35:20]
  reg  in_req_bits_r_wen; // @[Reg.scala 35:20]
  reg [1:0] in_req_bits_r_len; // @[Reg.scala 35:20]
  reg  in_req_bits_r_lrsc; // @[Reg.scala 35:20]
  reg [4:0] in_req_bits_r_amo; // @[Reg.scala 35:20]
  wire [38:0] _GEN_0 = _in_req_bits_T ? io_in_req_bits_addr : in_req_bits_r_addr; // @[Reg.scala 36:18 35:20 36:22]
  wire  _GEN_3 = _in_req_bits_T ? io_in_req_bits_wen : in_req_bits_r_wen; // @[Reg.scala 36:18 35:20 36:22]
  wire [11:0] in_vaddr_offset = _GEN_0[11:0]; // @[CachePortProxy.scala 25:46]
  wire [8:0] in_vaddr_vpn0 = _GEN_0[20:12]; // @[CachePortProxy.scala 25:46]
  wire [8:0] in_vaddr_vpn1 = _GEN_0[29:21]; // @[CachePortProxy.scala 25:46]
  wire [8:0] in_vaddr_vpn2 = _GEN_0[38:30]; // @[CachePortProxy.scala 25:46]
  wire  _atp_en_T_1 = io_prv != 2'h3 & io_sv39_en; // @[CachePortProxy.scala 38:48]
  reg  atp_en_r; // @[Reg.scala 35:20]
  wire  _GEN_7 = _in_req_bits_T ? _atp_en_T_1 : atp_en_r; // @[Reg.scala 36:18 35:20 36:22]
  wire  in_addr_boot = io_in_req_bits_addr >= 39'h10000 & io_in_req_bits_addr <= 39'h30000; // @[CachePortProxy.scala 42:50]
  wire  in_addr_clint = io_in_req_bits_addr >= 39'h2000000 & io_in_req_bits_addr <= 39'h200ffff; // @[CachePortProxy.scala 43:50]
  wire  in_addr_plic = io_in_req_bits_addr >= 39'hc000000 & io_in_req_bits_addr <= 39'hfffffff; // @[CachePortProxy.scala 44:50]
  wire  in_addr_uart = io_in_req_bits_addr >= 39'h10000000 & io_in_req_bits_addr <= 39'h1000ffff; // @[CachePortProxy.scala 45:50]
  wire  _access_fault_T_3 = ~_GEN_7; // @[CachePortProxy.scala 46:70]
  wire  _access_fault_T_9 = ~(in_addr_boot | in_addr_clint | in_addr_plic | in_addr_uart); // @[CachePortProxy.scala 47:5]
  wire  access_fault = ~io_in_req_bits_addr[31] & (io_prv == 2'h3 | ~_GEN_7) & _access_fault_T_9; // @[CachePortProxy.scala 46:79]
  reg [1:0] ptw_level; // @[CachePortProxy.scala 50:29]
  wire  ptw_pte_flag_v = io_ptw_resp_bits_rdata[0]; // @[CachePortProxy.scala 51:53]
  wire  ptw_pte_flag_r = io_ptw_resp_bits_rdata[1]; // @[CachePortProxy.scala 51:53]
  wire  ptw_pte_flag_w = io_ptw_resp_bits_rdata[2]; // @[CachePortProxy.scala 51:53]
  wire  ptw_pte_flag_x = io_ptw_resp_bits_rdata[3]; // @[CachePortProxy.scala 51:53]
  wire  ptw_pte_flag_u = io_ptw_resp_bits_rdata[4]; // @[CachePortProxy.scala 51:53]
  wire  ptw_pte_flag_g = io_ptw_resp_bits_rdata[5]; // @[CachePortProxy.scala 51:53]
  wire  ptw_pte_flag_a = io_ptw_resp_bits_rdata[6]; // @[CachePortProxy.scala 51:53]
  wire  ptw_pte_flag_d = io_ptw_resp_bits_rdata[7]; // @[CachePortProxy.scala 51:53]
  wire [8:0] ptw_pte_ppn0 = io_ptw_resp_bits_rdata[18:10]; // @[CachePortProxy.scala 51:53]
  wire [8:0] ptw_pte_ppn1 = io_ptw_resp_bits_rdata[27:19]; // @[CachePortProxy.scala 51:53]
  wire [1:0] ptw_pte_ppn2 = io_ptw_resp_bits_rdata[29:28]; // @[CachePortProxy.scala 51:53]
  wire  _ptw_pte_reg_T = io_ptw_resp_ready & io_ptw_resp_valid; // @[Decoupled.scala 51:35]
  reg [1:0] ptw_pte_reg_ppn2; // @[Reg.scala 35:20]
  reg [8:0] ptw_pte_reg_ppn1; // @[Reg.scala 35:20]
  reg [8:0] ptw_pte_reg_ppn0; // @[Reg.scala 35:20]
  reg  ptw_pte_reg_flag_d; // @[Reg.scala 35:20]
  reg  ptw_pte_reg_flag_a; // @[Reg.scala 35:20]
  reg  ptw_pte_reg_flag_g; // @[Reg.scala 35:20]
  reg  ptw_pte_reg_flag_u; // @[Reg.scala 35:20]
  reg  ptw_pte_reg_flag_x; // @[Reg.scala 35:20]
  reg  ptw_pte_reg_flag_w; // @[Reg.scala 35:20]
  reg  ptw_pte_reg_flag_r; // @[Reg.scala 35:20]
  reg  ptw_pte_reg_flag_v; // @[Reg.scala 35:20]
  wire  _ptw_complete_T_4 = ptw_pte_flag_r | ptw_pte_flag_x; // @[CachePortProxy.scala 7:37]
  wire  ptw_complete = ~ptw_pte_flag_v | ~ptw_pte_flag_r & ptw_pte_flag_w | _ptw_complete_T_4 | ptw_level == 2'h0; // @[CachePortProxy.scala 53:96]
  wire  _T_1 = io_in_req_ready & io_in_req_valid; // @[Decoupled.scala 51:35]
  wire  _T_2 = ~tlb_io_hit; // @[CachePortProxy.scala 59:24]
  wire [2:0] _GEN_20 = _GEN_7 & ~tlb_io_hit ? 3'h1 : state; // @[CachePortProxy.scala 59:37 60:17 21:93]
  wire [2:0] _GEN_21 = _T_1 ? _GEN_20 : state; // @[CachePortProxy.scala 58:28 21:93]
  wire  _T_7 = io_ptw_req_ready & io_ptw_req_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _ptw_level_T_1 = ptw_level - 2'h1; // @[CachePortProxy.scala 81:34]
  wire [2:0] _GEN_25 = ptw_complete ? 3'h3 : 3'h1; // @[CachePortProxy.scala 77:28 78:17 80:21]
  wire [1:0] _GEN_26 = ptw_complete ? ptw_level : _ptw_level_T_1; // @[CachePortProxy.scala 77:28 50:29 81:21]
  wire [2:0] _GEN_27 = _ptw_pte_reg_T ? _GEN_25 : state; // @[CachePortProxy.scala 76:30 21:93]
  wire [1:0] _GEN_28 = _ptw_pte_reg_T ? _GEN_26 : ptw_level; // @[CachePortProxy.scala 50:29 76:30]
  wire  _T_11 = io_out_req_ready & io_out_req_valid; // @[Decoupled.scala 51:35]
  wire  pte_flag_v = _in_req_bits_T ? tlb_io_rpte_flag_v : ptw_pte_reg_flag_v; // @[CachePortProxy.scala 121:18]
  wire  pte_flag_r = _in_req_bits_T ? tlb_io_rpte_flag_r : ptw_pte_reg_flag_r; // @[CachePortProxy.scala 121:18]
  wire  _T_16 = ~pte_flag_r; // @[CachePortProxy.scala 136:24]
  wire  pte_flag_w = _in_req_bits_T ? tlb_io_rpte_flag_w : ptw_pte_reg_flag_w; // @[CachePortProxy.scala 121:18]
  wire  pf1 = ~pte_flag_v | ~pte_flag_r & pte_flag_w; // @[CachePortProxy.scala 136:20]
  wire  pte_flag_x = _in_req_bits_T ? tlb_io_rpte_flag_x : ptw_pte_reg_flag_x; // @[CachePortProxy.scala 121:18]
  wire  _T_19 = pte_flag_r | pte_flag_x; // @[CachePortProxy.scala 7:37]
  wire  pte_flag_a = _in_req_bits_T ? tlb_io_rpte_flag_a : ptw_pte_reg_flag_a; // @[CachePortProxy.scala 121:18]
  wire  _T_20 = ~pte_flag_a; // @[CachePortProxy.scala 140:10]
  wire  pf2 = _T_19 & _T_20; // @[CachePortProxy.scala 139:21 132:24]
  reg [1:0] prv_r; // @[Reg.scala 35:20]
  wire [1:0] prv = _in_req_bits_T ? io_prv : prv_r; // @[Utils.scala 50:8]
  wire  pte_flag_u = _in_req_bits_T ? tlb_io_rpte_flag_u : ptw_pte_reg_flag_u; // @[CachePortProxy.scala 121:18]
  wire  _T_23 = prv == 2'h0 & ~pte_flag_u; // @[CachePortProxy.scala 143:26]
  wire  pf3 = _T_19 & _T_23; // @[CachePortProxy.scala 139:21 133:24]
  wire  pte_flag_d = _in_req_bits_T ? tlb_io_rpte_flag_d : ptw_pte_reg_flag_d; // @[CachePortProxy.scala 121:18]
  wire  _T_29 = _GEN_3 & (~pte_flag_w | _T_16 | ~pte_flag_d); // @[CachePortProxy.scala 152:28]
  wire  pf4 = _T_19 & _T_29; // @[CachePortProxy.scala 139:21 134:24]
  wire  _T_30 = state == 3'h3; // @[CachePortProxy.scala 156:16]
  wire [8:0] pte_ppn1 = _in_req_bits_T ? tlb_io_rpte_ppn1 : ptw_pte_reg_ppn1; // @[CachePortProxy.scala 121:18]
  wire [8:0] pte_ppn0 = _in_req_bits_T ? tlb_io_rpte_ppn0 : ptw_pte_reg_ppn0; // @[CachePortProxy.scala 121:18]
  wire [17:0] _T_32 = {pte_ppn1,pte_ppn0}; // @[Cat.scala 33:92]
  wire  _T_38 = ptw_level == 2'h2 & _T_32 != 18'h0 | ptw_level == 2'h1 & pte_ppn0 != 9'h0; // @[CachePortProxy.scala 157:67]
  wire  _GEN_45 = state == 3'h3 & _T_38; // @[CachePortProxy.scala 135:24 156:36]
  wire  pf5 = _T_19 & _GEN_45; // @[CachePortProxy.scala 139:21 135:24]
  wire  page_fault = pf1 | pf2 | pf3 | pf4 | pf5; // @[CachePortProxy.scala 162:42]
  wire [2:0] _GEN_29 = _T_11 | page_fault ? 3'h0 : state; // @[CachePortProxy.scala 86:43 87:15 21:93]
  wire  _T_14 = io_in_resp_ready & io_in_resp_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_30 = _T_14 ? 3'h0 : state; // @[CachePortProxy.scala 91:29 92:15 21:93]
  wire [2:0] _GEN_31 = 3'h4 == state ? _GEN_30 : state; // @[CachePortProxy.scala 56:17 21:93]
  wire [2:0] _GEN_32 = 3'h3 == state ? _GEN_29 : _GEN_31; // @[CachePortProxy.scala 56:17]
  wire [55:0] _l2_addr_T = {io_satp_ppn,in_vaddr_vpn2,3'h0}; // @[Cat.scala 33:92]
  wire [31:0] l1_addr = {ptw_pte_reg_ppn2,ptw_pte_reg_ppn1,ptw_pte_reg_ppn0,in_vaddr_vpn1,3'h0}; // @[Cat.scala 33:92]
  wire [31:0] l0_addr = {ptw_pte_reg_ppn2,ptw_pte_reg_ppn1,ptw_pte_reg_ppn0,in_vaddr_vpn0,3'h0}; // @[Cat.scala 33:92]
  wire [31:0] l2_addr = _l2_addr_T[31:0]; // @[CachePortProxy.scala 102:11 98:21]
  wire [31:0] _io_ptw_req_bits_addr_T_1 = 2'h2 == ptw_level ? l2_addr : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] _io_ptw_req_bits_addr_T_3 = 2'h1 == ptw_level ? l1_addr : _io_ptw_req_bits_addr_T_1; // @[Mux.scala 81:58]
  wire [31:0] _io_ptw_req_bits_addr_T_5 = 2'h0 == ptw_level ? l0_addr : _io_ptw_req_bits_addr_T_3; // @[Mux.scala 81:58]
  wire [1:0] pte_ppn2 = _in_req_bits_T ? tlb_io_rpte_ppn2 : ptw_pte_reg_ppn2; // @[CachePortProxy.scala 121:18]
  wire [1:0] level = _in_req_bits_T ? tlb_io_rlevel : ptw_level; // @[CachePortProxy.scala 122:18]
  wire  _tlb_io_wen_T_1 = ~page_fault; // @[CachePortProxy.scala 125:50]
  wire  _tlb_io_wen_T_2 = _T_30 & ~page_fault; // @[CachePortProxy.scala 125:47]
  wire [8:0] paddr_ppn0 = level > 2'h0 ? in_vaddr_vpn0 : pte_ppn0; // @[CachePortProxy.scala 167:22]
  wire [8:0] paddr_ppn1 = level > 2'h1 ? in_vaddr_vpn1 : pte_ppn1; // @[CachePortProxy.scala 168:22]
  wire [31:0] _io_out_req_bits_addr_T = {pte_ppn2,paddr_ppn1,paddr_ppn0,in_vaddr_offset}; // @[CachePortProxy.scala 177:43]
  wire [38:0] _io_out_req_bits_addr_WIRE = {{7'd0}, _io_out_req_bits_addr_T}; // @[CachePortProxy.scala 177:{43,43}]
  wire  _page_fault_reg_T_7 = page_fault & _GEN_7 & (_in_req_bits_T & tlb_io_hit & _T_1 | _T_30); // @[CachePortProxy.scala 182:26]
  reg  page_fault_reg; // @[Utils.scala 36:20]
  wire  _GEN_51 = _page_fault_reg_T_7 | page_fault_reg; // @[Utils.scala 41:19 36:20 41:23]
  TLB tlb ( // @[CachePortProxy.scala 28:19]
    .clock(tlb_clock),
    .reset(tlb_reset),
    .io_sfence_vma(tlb_io_sfence_vma),
    .io_vaddr_vpn2(tlb_io_vaddr_vpn2),
    .io_vaddr_vpn1(tlb_io_vaddr_vpn1),
    .io_vaddr_vpn0(tlb_io_vaddr_vpn0),
    .io_rpte_ppn2(tlb_io_rpte_ppn2),
    .io_rpte_ppn1(tlb_io_rpte_ppn1),
    .io_rpte_ppn0(tlb_io_rpte_ppn0),
    .io_rpte_flag_d(tlb_io_rpte_flag_d),
    .io_rpte_flag_a(tlb_io_rpte_flag_a),
    .io_rpte_flag_u(tlb_io_rpte_flag_u),
    .io_rpte_flag_x(tlb_io_rpte_flag_x),
    .io_rpte_flag_w(tlb_io_rpte_flag_w),
    .io_rpte_flag_r(tlb_io_rpte_flag_r),
    .io_rpte_flag_v(tlb_io_rpte_flag_v),
    .io_rlevel(tlb_io_rlevel),
    .io_hit(tlb_io_hit),
    .io_wen(tlb_io_wen),
    .io_wvaddr_vpn2(tlb_io_wvaddr_vpn2),
    .io_wvaddr_vpn1(tlb_io_wvaddr_vpn1),
    .io_wvaddr_vpn0(tlb_io_wvaddr_vpn0),
    .io_wpte_ppn2(tlb_io_wpte_ppn2),
    .io_wpte_ppn1(tlb_io_wpte_ppn1),
    .io_wpte_ppn0(tlb_io_wpte_ppn0),
    .io_wpte_flag_d(tlb_io_wpte_flag_d),
    .io_wpte_flag_a(tlb_io_wpte_flag_a),
    .io_wpte_flag_g(tlb_io_wpte_flag_g),
    .io_wpte_flag_u(tlb_io_wpte_flag_u),
    .io_wpte_flag_x(tlb_io_wpte_flag_x),
    .io_wpte_flag_w(tlb_io_wpte_flag_w),
    .io_wpte_flag_r(tlb_io_wpte_flag_r),
    .io_wpte_flag_v(tlb_io_wpte_flag_v),
    .io_wlevel(tlb_io_wlevel),
    .io_satp_asid(tlb_io_satp_asid)
  );
  assign io_in_req_ready = _in_req_bits_T & (io_out_req_ready | access_fault | _GEN_7 & (_T_2 | page_fault)); // @[CachePortProxy.scala 172:41]
  assign io_in_resp_valid = io_out_resp_valid | io_in_resp_bits_page_fault | io_in_resp_bits_access_fault; // @[CachePortProxy.scala 189:83]
  assign io_in_resp_bits_rdata = io_out_resp_bits_rdata; // @[CachePortProxy.scala 185:32]
  assign io_in_resp_bits_page_fault = page_fault_reg; // @[CachePortProxy.scala 186:32]
  assign io_in_resp_bits_access_fault = state == 3'h4; // @[CachePortProxy.scala 187:42]
  assign io_out_req_valid = _in_req_bits_T & (tlb_io_hit & _tlb_io_wen_T_1 | _access_fault_T_3 & ~access_fault) &
    io_in_req_valid | _tlb_io_wen_T_2; // @[CachePortProxy.scala 173:126]
  assign io_out_req_bits_addr = _GEN_7 ? _io_out_req_bits_addr_WIRE : _GEN_0; // @[CachePortProxy.scala 176:16 175:19 177:26]
  assign io_out_req_bits_wdata = _in_req_bits_T ? io_in_req_bits_wdata : in_req_bits_r_wdata; // @[Utils.scala 50:8]
  assign io_out_req_bits_wmask = _in_req_bits_T ? io_in_req_bits_wmask : in_req_bits_r_wmask; // @[Utils.scala 50:8]
  assign io_out_req_bits_wen = _in_req_bits_T ? io_in_req_bits_wen : in_req_bits_r_wen; // @[Utils.scala 50:8]
  assign io_out_req_bits_len = _in_req_bits_T ? io_in_req_bits_len : in_req_bits_r_len; // @[Utils.scala 50:8]
  assign io_out_req_bits_lrsc = _in_req_bits_T ? io_in_req_bits_lrsc : in_req_bits_r_lrsc; // @[Utils.scala 50:8]
  assign io_out_req_bits_amo = _in_req_bits_T ? io_in_req_bits_amo : in_req_bits_r_amo; // @[Utils.scala 50:8]
  assign io_out_resp_ready = io_in_resp_ready; // @[CachePortProxy.scala 190:32]
  assign io_ptw_req_valid = state == 3'h1; // @[CachePortProxy.scala 117:31]
  assign io_ptw_req_bits_addr = {{7'd0}, _io_ptw_req_bits_addr_T_5}; // @[CachePortProxy.scala 108:24]
  assign io_ptw_resp_ready = state == 3'h2; // @[CachePortProxy.scala 118:31]
  assign tlb_clock = clock;
  assign tlb_reset = reset;
  assign tlb_io_sfence_vma = io_sfence_vma; // @[CachePortProxy.scala 31:21]
  assign tlb_io_vaddr_vpn2 = io_in_req_bits_addr[38:30]; // @[CachePortProxy.scala 32:52]
  assign tlb_io_vaddr_vpn1 = io_in_req_bits_addr[29:21]; // @[CachePortProxy.scala 32:52]
  assign tlb_io_vaddr_vpn0 = io_in_req_bits_addr[20:12]; // @[CachePortProxy.scala 32:52]
  assign tlb_io_wen = _T_30 & ~page_fault; // @[CachePortProxy.scala 125:47]
  assign tlb_io_wvaddr_vpn2 = _GEN_0[38:30]; // @[CachePortProxy.scala 25:46]
  assign tlb_io_wvaddr_vpn1 = _GEN_0[29:21]; // @[CachePortProxy.scala 25:46]
  assign tlb_io_wvaddr_vpn0 = _GEN_0[20:12]; // @[CachePortProxy.scala 25:46]
  assign tlb_io_wpte_ppn2 = ptw_pte_reg_ppn2; // @[CachePortProxy.scala 127:17]
  assign tlb_io_wpte_ppn1 = ptw_pte_reg_ppn1; // @[CachePortProxy.scala 127:17]
  assign tlb_io_wpte_ppn0 = ptw_pte_reg_ppn0; // @[CachePortProxy.scala 127:17]
  assign tlb_io_wpte_flag_d = ptw_pte_reg_flag_d; // @[CachePortProxy.scala 127:17]
  assign tlb_io_wpte_flag_a = ptw_pte_reg_flag_a; // @[CachePortProxy.scala 127:17]
  assign tlb_io_wpte_flag_g = ptw_pte_reg_flag_g; // @[CachePortProxy.scala 127:17]
  assign tlb_io_wpte_flag_u = ptw_pte_reg_flag_u; // @[CachePortProxy.scala 127:17]
  assign tlb_io_wpte_flag_x = ptw_pte_reg_flag_x; // @[CachePortProxy.scala 127:17]
  assign tlb_io_wpte_flag_w = ptw_pte_reg_flag_w; // @[CachePortProxy.scala 127:17]
  assign tlb_io_wpte_flag_r = ptw_pte_reg_flag_r; // @[CachePortProxy.scala 127:17]
  assign tlb_io_wpte_flag_v = ptw_pte_reg_flag_v; // @[CachePortProxy.scala 127:17]
  assign tlb_io_wlevel = ptw_level; // @[CachePortProxy.scala 128:17]
  assign tlb_io_satp_asid = io_satp_asid; // @[CachePortProxy.scala 30:21]
  always @(posedge clock) begin
    if (reset) begin // @[CachePortProxy.scala 21:93]
      state <= 3'h0; // @[CachePortProxy.scala 21:93]
    end else if (3'h0 == state) begin // @[CachePortProxy.scala 56:17]
      if (io_in_req_valid) begin // @[CachePortProxy.scala 63:29]
        if (_access_fault_T_3 & access_fault) begin // @[CachePortProxy.scala 64:39]
          state <= 3'h4; // @[CachePortProxy.scala 65:17]
        end else begin
          state <= _GEN_21;
        end
      end else begin
        state <= _GEN_21;
      end
    end else if (3'h1 == state) begin // @[CachePortProxy.scala 56:17]
      if (_T_7) begin // @[CachePortProxy.scala 71:29]
        state <= 3'h2; // @[CachePortProxy.scala 72:15]
      end
    end else if (3'h2 == state) begin // @[CachePortProxy.scala 56:17]
      state <= _GEN_27;
    end else begin
      state <= _GEN_32;
    end
    if (reset) begin // @[Reg.scala 35:20]
      in_req_bits_r_addr <= 39'h0; // @[Reg.scala 35:20]
    end else if (_in_req_bits_T) begin // @[Reg.scala 36:18]
      in_req_bits_r_addr <= io_in_req_bits_addr; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      in_req_bits_r_wdata <= 64'h0; // @[Reg.scala 35:20]
    end else if (_in_req_bits_T) begin // @[Reg.scala 36:18]
      in_req_bits_r_wdata <= io_in_req_bits_wdata; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      in_req_bits_r_wmask <= 8'h0; // @[Reg.scala 35:20]
    end else if (_in_req_bits_T) begin // @[Reg.scala 36:18]
      in_req_bits_r_wmask <= io_in_req_bits_wmask; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      in_req_bits_r_wen <= 1'h0; // @[Reg.scala 35:20]
    end else if (_in_req_bits_T) begin // @[Reg.scala 36:18]
      in_req_bits_r_wen <= io_in_req_bits_wen; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      in_req_bits_r_len <= 2'h0; // @[Reg.scala 35:20]
    end else if (_in_req_bits_T) begin // @[Reg.scala 36:18]
      in_req_bits_r_len <= io_in_req_bits_len; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      in_req_bits_r_lrsc <= 1'h0; // @[Reg.scala 35:20]
    end else if (_in_req_bits_T) begin // @[Reg.scala 36:18]
      in_req_bits_r_lrsc <= io_in_req_bits_lrsc; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      in_req_bits_r_amo <= 5'h0; // @[Reg.scala 35:20]
    end else if (_in_req_bits_T) begin // @[Reg.scala 36:18]
      in_req_bits_r_amo <= io_in_req_bits_amo; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      atp_en_r <= 1'h0; // @[Reg.scala 35:20]
    end else if (_in_req_bits_T) begin // @[Reg.scala 36:18]
      atp_en_r <= _atp_en_T_1; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[CachePortProxy.scala 50:29]
      ptw_level <= 2'h0; // @[CachePortProxy.scala 50:29]
    end else if (3'h0 == state) begin // @[CachePortProxy.scala 56:17]
      ptw_level <= 2'h2; // @[CachePortProxy.scala 68:17]
    end else if (!(3'h1 == state)) begin // @[CachePortProxy.scala 56:17]
      if (3'h2 == state) begin // @[CachePortProxy.scala 56:17]
        ptw_level <= _GEN_28;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      ptw_pte_reg_ppn2 <= 2'h0; // @[Reg.scala 35:20]
    end else if (_ptw_pte_reg_T) begin // @[Reg.scala 36:18]
      ptw_pte_reg_ppn2 <= ptw_pte_ppn2; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ptw_pte_reg_ppn1 <= 9'h0; // @[Reg.scala 35:20]
    end else if (_ptw_pte_reg_T) begin // @[Reg.scala 36:18]
      ptw_pte_reg_ppn1 <= ptw_pte_ppn1; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ptw_pte_reg_ppn0 <= 9'h0; // @[Reg.scala 35:20]
    end else if (_ptw_pte_reg_T) begin // @[Reg.scala 36:18]
      ptw_pte_reg_ppn0 <= ptw_pte_ppn0; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ptw_pte_reg_flag_d <= 1'h0; // @[Reg.scala 35:20]
    end else if (_ptw_pte_reg_T) begin // @[Reg.scala 36:18]
      ptw_pte_reg_flag_d <= ptw_pte_flag_d; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ptw_pte_reg_flag_a <= 1'h0; // @[Reg.scala 35:20]
    end else if (_ptw_pte_reg_T) begin // @[Reg.scala 36:18]
      ptw_pte_reg_flag_a <= ptw_pte_flag_a; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ptw_pte_reg_flag_g <= 1'h0; // @[Reg.scala 35:20]
    end else if (_ptw_pte_reg_T) begin // @[Reg.scala 36:18]
      ptw_pte_reg_flag_g <= ptw_pte_flag_g; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ptw_pte_reg_flag_u <= 1'h0; // @[Reg.scala 35:20]
    end else if (_ptw_pte_reg_T) begin // @[Reg.scala 36:18]
      ptw_pte_reg_flag_u <= ptw_pte_flag_u; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ptw_pte_reg_flag_x <= 1'h0; // @[Reg.scala 35:20]
    end else if (_ptw_pte_reg_T) begin // @[Reg.scala 36:18]
      ptw_pte_reg_flag_x <= ptw_pte_flag_x; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ptw_pte_reg_flag_w <= 1'h0; // @[Reg.scala 35:20]
    end else if (_ptw_pte_reg_T) begin // @[Reg.scala 36:18]
      ptw_pte_reg_flag_w <= ptw_pte_flag_w; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ptw_pte_reg_flag_r <= 1'h0; // @[Reg.scala 35:20]
    end else if (_ptw_pte_reg_T) begin // @[Reg.scala 36:18]
      ptw_pte_reg_flag_r <= ptw_pte_flag_r; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ptw_pte_reg_flag_v <= 1'h0; // @[Reg.scala 35:20]
    end else if (_ptw_pte_reg_T) begin // @[Reg.scala 36:18]
      ptw_pte_reg_flag_v <= ptw_pte_flag_v; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      prv_r <= 2'h0; // @[Reg.scala 35:20]
    end else if (_in_req_bits_T) begin // @[Utils.scala 50:8]
      prv_r <= io_prv;
    end
    if (reset) begin // @[Utils.scala 36:20]
      page_fault_reg <= 1'h0; // @[Utils.scala 36:20]
    end else if (_T_14) begin // @[Utils.scala 42:18]
      page_fault_reg <= 1'h0; // @[Utils.scala 42:22]
    end else begin
      page_fault_reg <= _GEN_51;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {2{`RANDOM}};
  in_req_bits_r_addr = _RAND_1[38:0];
  _RAND_2 = {2{`RANDOM}};
  in_req_bits_r_wdata = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  in_req_bits_r_wmask = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  in_req_bits_r_wen = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  in_req_bits_r_len = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  in_req_bits_r_lrsc = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  in_req_bits_r_amo = _RAND_7[4:0];
  _RAND_8 = {1{`RANDOM}};
  atp_en_r = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  ptw_level = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  ptw_pte_reg_ppn2 = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  ptw_pte_reg_ppn1 = _RAND_11[8:0];
  _RAND_12 = {1{`RANDOM}};
  ptw_pte_reg_ppn0 = _RAND_12[8:0];
  _RAND_13 = {1{`RANDOM}};
  ptw_pte_reg_flag_d = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  ptw_pte_reg_flag_a = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  ptw_pte_reg_flag_g = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  ptw_pte_reg_flag_u = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  ptw_pte_reg_flag_x = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  ptw_pte_reg_flag_w = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  ptw_pte_reg_flag_r = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  ptw_pte_reg_flag_v = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  prv_r = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  page_fault_reg = _RAND_22[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CachePortXBar1to2(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [38:0] io_in_req_bits_addr,
  input  [63:0] io_in_req_bits_wdata,
  input  [7:0]  io_in_req_bits_wmask,
  input         io_in_req_bits_wen,
  input  [1:0]  io_in_req_bits_len,
  input         io_in_req_bits_lrsc,
  input  [4:0]  io_in_req_bits_amo,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_0_req_ready,
  output        io_out_0_req_valid,
  output [38:0] io_out_0_req_bits_addr,
  output [63:0] io_out_0_req_bits_wdata,
  output [7:0]  io_out_0_req_bits_wmask,
  output        io_out_0_req_bits_wen,
  output [1:0]  io_out_0_req_bits_len,
  output        io_out_0_req_bits_lrsc,
  output [4:0]  io_out_0_req_bits_amo,
  output        io_out_0_resp_ready,
  input         io_out_0_resp_valid,
  input  [63:0] io_out_0_resp_bits_rdata,
  input         io_out_1_req_ready,
  output        io_out_1_req_valid,
  output [38:0] io_out_1_req_bits_addr,
  output [63:0] io_out_1_req_bits_wdata,
  output [7:0]  io_out_1_req_bits_wmask,
  output        io_out_1_req_bits_wen,
  output [1:0]  io_out_1_req_bits_len,
  output        io_out_1_resp_ready,
  input         io_out_1_resp_valid,
  input  [63:0] io_out_1_resp_bits_rdata,
  input         io_to_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  _to_1_r_T = io_in_req_ready & io_in_req_valid; // @[Decoupled.scala 51:35]
  reg  to_1_r; // @[Reg.scala 35:20]
  assign io_in_req_ready = io_to_1 ? io_out_1_req_ready : io_out_0_req_ready; // @[Bus.scala 100:29]
  assign io_in_resp_valid = to_1_r ? io_out_1_resp_valid : io_out_0_resp_valid; // @[Bus.scala 104:30]
  assign io_in_resp_bits_rdata = to_1_r ? io_out_1_resp_bits_rdata : io_out_0_resp_bits_rdata; // @[Bus.scala 103:30]
  assign io_out_0_req_valid = io_in_req_valid & ~io_to_1; // @[Bus.scala 98:42]
  assign io_out_0_req_bits_addr = io_in_req_bits_addr; // @[Bus.scala 96:23]
  assign io_out_0_req_bits_wdata = io_in_req_bits_wdata; // @[Bus.scala 96:23]
  assign io_out_0_req_bits_wmask = io_in_req_bits_wmask; // @[Bus.scala 96:23]
  assign io_out_0_req_bits_wen = io_in_req_bits_wen; // @[Bus.scala 96:23]
  assign io_out_0_req_bits_len = io_in_req_bits_len; // @[Bus.scala 96:23]
  assign io_out_0_req_bits_lrsc = io_in_req_bits_lrsc; // @[Bus.scala 96:23]
  assign io_out_0_req_bits_amo = io_in_req_bits_amo; // @[Bus.scala 96:23]
  assign io_out_0_resp_ready = io_in_resp_ready; // @[Bus.scala 106:24]
  assign io_out_1_req_valid = io_in_req_valid & io_to_1; // @[Bus.scala 99:42]
  assign io_out_1_req_bits_addr = io_in_req_bits_addr; // @[Bus.scala 97:23]
  assign io_out_1_req_bits_wdata = io_in_req_bits_wdata; // @[Bus.scala 97:23]
  assign io_out_1_req_bits_wmask = io_in_req_bits_wmask; // @[Bus.scala 97:23]
  assign io_out_1_req_bits_wen = io_in_req_bits_wen; // @[Bus.scala 97:23]
  assign io_out_1_req_bits_len = io_in_req_bits_len; // @[Bus.scala 97:23]
  assign io_out_1_resp_ready = io_in_resp_ready; // @[Bus.scala 107:24]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 35:20]
      to_1_r <= 1'h0; // @[Reg.scala 35:20]
    end else if (_to_1_r_T) begin // @[Reg.scala 36:18]
      to_1_r <= io_to_1; // @[Reg.scala 36:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  to_1_r = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PipelineReg_1(
  input         clock,
  input         reset,
  input         io_in_uop_valid,
  input  [4:0]  io_in_uop_rd_index,
  input         io_in_uop_rd_wen,
  input  [63:0] io_in_rd_data,
  output        io_out_uop_valid,
  output [4:0]  io_out_uop_rd_index,
  output        io_out_uop_rd_wen,
  output [63:0] io_out_rd_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg  reg_uop_valid; // @[Reg.scala 35:20]
  reg [4:0] reg_uop_rd_index; // @[Reg.scala 35:20]
  reg  reg_uop_rd_wen; // @[Reg.scala 35:20]
  reg [63:0] reg_rd_data; // @[Reg.scala 35:20]
  assign io_out_uop_valid = reg_uop_valid; // @[DataType.scala 41:10]
  assign io_out_uop_rd_index = reg_uop_rd_index; // @[DataType.scala 41:10]
  assign io_out_uop_rd_wen = reg_uop_rd_wen; // @[DataType.scala 41:10]
  assign io_out_rd_data = reg_rd_data; // @[DataType.scala 41:10]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 35:20]
      reg_uop_valid <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      reg_uop_valid <= io_in_uop_valid;
    end
    if (reset) begin // @[Reg.scala 35:20]
      reg_uop_rd_index <= 5'h0; // @[Reg.scala 35:20]
    end else begin
      reg_uop_rd_index <= io_in_uop_rd_index;
    end
    if (reset) begin // @[Reg.scala 35:20]
      reg_uop_rd_wen <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      reg_uop_rd_wen <= io_in_uop_rd_wen;
    end
    if (reset) begin // @[Reg.scala 35:20]
      reg_rd_data <= 64'h0; // @[Reg.scala 35:20]
    end else begin
      reg_rd_data <= io_in_rd_data;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_uop_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  reg_uop_rd_index = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  reg_uop_rd_wen = _RAND_2[0:0];
  _RAND_3 = {2{`RANDOM}};
  reg_rd_data = _RAND_3[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Core(
  input         clock,
  input         reset,
  input         io_imem_req_ready,
  output        io_imem_req_valid,
  output [38:0] io_imem_req_bits_addr,
  output        io_imem_resp_ready,
  input         io_imem_resp_valid,
  input  [63:0] io_imem_resp_bits_rdata,
  input         io_dmem_req_ready,
  output        io_dmem_req_valid,
  output [38:0] io_dmem_req_bits_addr,
  output [63:0] io_dmem_req_bits_wdata,
  output [7:0]  io_dmem_req_bits_wmask,
  output        io_dmem_req_bits_wen,
  output [1:0]  io_dmem_req_bits_len,
  output        io_dmem_req_bits_lrsc,
  output [4:0]  io_dmem_req_bits_amo,
  output        io_dmem_resp_ready,
  input         io_dmem_resp_valid,
  input  [63:0] io_dmem_resp_bits_rdata,
  input         io_iptw_req_ready,
  output        io_iptw_req_valid,
  output [38:0] io_iptw_req_bits_addr,
  output        io_iptw_resp_ready,
  input         io_iptw_resp_valid,
  input  [63:0] io_iptw_resp_bits_rdata,
  input         io_dptw_req_ready,
  output        io_dptw_req_valid,
  output [38:0] io_dptw_req_bits_addr,
  output        io_dptw_resp_ready,
  input         io_dptw_resp_valid,
  input  [63:0] io_dptw_resp_bits_rdata,
  input         io_uncache_req_ready,
  output        io_uncache_req_valid,
  output [38:0] io_uncache_req_bits_addr,
  output [63:0] io_uncache_req_bits_wdata,
  output [7:0]  io_uncache_req_bits_wmask,
  output        io_uncache_req_bits_wen,
  output [1:0]  io_uncache_req_bits_len,
  output        io_uncache_resp_ready,
  input         io_uncache_resp_valid,
  input  [63:0] io_uncache_resp_bits_rdata,
  output        io_fence_i,
  input         io_intr_mtip,
  input         io_intr_msip,
  input         io_intr_meip,
  input         io_intr_seip
);
  wire  ifu_clock; // @[Core.scala 27:19]
  wire  ifu_reset; // @[Core.scala 27:19]
  wire  ifu_io_jmp_packet_valid; // @[Core.scala 27:19]
  wire [63:0] ifu_io_jmp_packet_target; // @[Core.scala 27:19]
  wire  ifu_io_jmp_packet_bp_update; // @[Core.scala 27:19]
  wire  ifu_io_jmp_packet_bp_taken; // @[Core.scala 27:19]
  wire [63:0] ifu_io_jmp_packet_bp_pc; // @[Core.scala 27:19]
  wire  ifu_io_imem_req_ready; // @[Core.scala 27:19]
  wire  ifu_io_imem_req_valid; // @[Core.scala 27:19]
  wire [38:0] ifu_io_imem_req_bits_addr; // @[Core.scala 27:19]
  wire  ifu_io_imem_resp_ready; // @[Core.scala 27:19]
  wire  ifu_io_imem_resp_valid; // @[Core.scala 27:19]
  wire [63:0] ifu_io_imem_resp_bits_rdata; // @[Core.scala 27:19]
  wire  ifu_io_imem_resp_bits_page_fault; // @[Core.scala 27:19]
  wire  ifu_io_imem_resp_bits_access_fault; // @[Core.scala 27:19]
  wire [63:0] ifu_io_out_pc; // @[Core.scala 27:19]
  wire [31:0] ifu_io_out_instr; // @[Core.scala 27:19]
  wire  ifu_io_out_valid; // @[Core.scala 27:19]
  wire  ifu_io_out_page_fault; // @[Core.scala 27:19]
  wire  ifu_io_out_access_fault; // @[Core.scala 27:19]
  wire [63:0] ifu_io_out_bp_npc; // @[Core.scala 27:19]
  wire  ifu_io_stall_b; // @[Core.scala 27:19]
  wire  imem_proxy_clock; // @[Core.scala 28:26]
  wire  imem_proxy_reset; // @[Core.scala 28:26]
  wire [1:0] imem_proxy_io_prv; // @[Core.scala 28:26]
  wire  imem_proxy_io_sv39_en; // @[Core.scala 28:26]
  wire [15:0] imem_proxy_io_satp_asid; // @[Core.scala 28:26]
  wire [43:0] imem_proxy_io_satp_ppn; // @[Core.scala 28:26]
  wire  imem_proxy_io_sfence_vma; // @[Core.scala 28:26]
  wire  imem_proxy_io_in_req_ready; // @[Core.scala 28:26]
  wire  imem_proxy_io_in_req_valid; // @[Core.scala 28:26]
  wire [38:0] imem_proxy_io_in_req_bits_addr; // @[Core.scala 28:26]
  wire  imem_proxy_io_in_resp_ready; // @[Core.scala 28:26]
  wire  imem_proxy_io_in_resp_valid; // @[Core.scala 28:26]
  wire [63:0] imem_proxy_io_in_resp_bits_rdata; // @[Core.scala 28:26]
  wire  imem_proxy_io_in_resp_bits_page_fault; // @[Core.scala 28:26]
  wire  imem_proxy_io_in_resp_bits_access_fault; // @[Core.scala 28:26]
  wire  imem_proxy_io_out_req_ready; // @[Core.scala 28:26]
  wire  imem_proxy_io_out_req_valid; // @[Core.scala 28:26]
  wire [38:0] imem_proxy_io_out_req_bits_addr; // @[Core.scala 28:26]
  wire  imem_proxy_io_out_resp_ready; // @[Core.scala 28:26]
  wire  imem_proxy_io_out_resp_valid; // @[Core.scala 28:26]
  wire [63:0] imem_proxy_io_out_resp_bits_rdata; // @[Core.scala 28:26]
  wire  imem_proxy_io_ptw_req_ready; // @[Core.scala 28:26]
  wire  imem_proxy_io_ptw_req_valid; // @[Core.scala 28:26]
  wire [38:0] imem_proxy_io_ptw_req_bits_addr; // @[Core.scala 28:26]
  wire  imem_proxy_io_ptw_resp_ready; // @[Core.scala 28:26]
  wire  imem_proxy_io_ptw_resp_valid; // @[Core.scala 28:26]
  wire [63:0] imem_proxy_io_ptw_resp_bits_rdata; // @[Core.scala 28:26]
  wire  instr_buffer_clock; // @[Core.scala 54:28]
  wire  instr_buffer_reset; // @[Core.scala 54:28]
  wire  instr_buffer_io_enq_ready; // @[Core.scala 54:28]
  wire  instr_buffer_io_enq_valid; // @[Core.scala 54:28]
  wire [63:0] instr_buffer_io_enq_bits_pc; // @[Core.scala 54:28]
  wire [31:0] instr_buffer_io_enq_bits_instr; // @[Core.scala 54:28]
  wire  instr_buffer_io_enq_bits_page_fault; // @[Core.scala 54:28]
  wire  instr_buffer_io_enq_bits_access_fault; // @[Core.scala 54:28]
  wire [63:0] instr_buffer_io_enq_bits_bp_npc; // @[Core.scala 54:28]
  wire  instr_buffer_io_deq_ready; // @[Core.scala 54:28]
  wire  instr_buffer_io_deq_valid; // @[Core.scala 54:28]
  wire [63:0] instr_buffer_io_deq_bits_pc; // @[Core.scala 54:28]
  wire [31:0] instr_buffer_io_deq_bits_instr; // @[Core.scala 54:28]
  wire  instr_buffer_io_deq_bits_page_fault; // @[Core.scala 54:28]
  wire  instr_buffer_io_deq_bits_access_fault; // @[Core.scala 54:28]
  wire [63:0] instr_buffer_io_deq_bits_bp_npc; // @[Core.scala 54:28]
  wire  instr_buffer_io_flush; // @[Core.scala 54:28]
  wire [63:0] decode_io_in_pc; // @[Core.scala 63:22]
  wire [31:0] decode_io_in_instr; // @[Core.scala 63:22]
  wire  decode_io_in_valid; // @[Core.scala 63:22]
  wire  decode_io_in_page_fault; // @[Core.scala 63:22]
  wire  decode_io_in_access_fault; // @[Core.scala 63:22]
  wire  decode_io_out_valid; // @[Core.scala 63:22]
  wire [2:0] decode_io_out_exc; // @[Core.scala 63:22]
  wire [63:0] decode_io_out_pc; // @[Core.scala 63:22]
  wire [63:0] decode_io_out_npc; // @[Core.scala 63:22]
  wire [31:0] decode_io_out_instr; // @[Core.scala 63:22]
  wire [2:0] decode_io_out_fu; // @[Core.scala 63:22]
  wire [3:0] decode_io_out_alu_op; // @[Core.scala 63:22]
  wire [1:0] decode_io_out_jmp_op; // @[Core.scala 63:22]
  wire [3:0] decode_io_out_mdu_op; // @[Core.scala 63:22]
  wire [4:0] decode_io_out_lsu_op; // @[Core.scala 63:22]
  wire [1:0] decode_io_out_mem_len; // @[Core.scala 63:22]
  wire [1:0] decode_io_out_csr_op; // @[Core.scala 63:22]
  wire [2:0] decode_io_out_sys_op; // @[Core.scala 63:22]
  wire [1:0] decode_io_out_rs1_src; // @[Core.scala 63:22]
  wire [1:0] decode_io_out_rs2_src; // @[Core.scala 63:22]
  wire [4:0] decode_io_out_rs1_index; // @[Core.scala 63:22]
  wire [4:0] decode_io_out_rs2_index; // @[Core.scala 63:22]
  wire [4:0] decode_io_out_rd_index; // @[Core.scala 63:22]
  wire  decode_io_out_rd_wen; // @[Core.scala 63:22]
  wire [31:0] decode_io_out_imm; // @[Core.scala 63:22]
  wire  decode_io_out_dw; // @[Core.scala 63:22]
  wire  rf_clock; // @[Core.scala 67:18]
  wire  rf_reset; // @[Core.scala 67:18]
  wire [4:0] rf_io_rs1_index; // @[Core.scala 67:18]
  wire [4:0] rf_io_rs2_index; // @[Core.scala 67:18]
  wire [63:0] rf_io_rs1_data; // @[Core.scala 67:18]
  wire [63:0] rf_io_rs2_data; // @[Core.scala 67:18]
  wire [4:0] rf_io_rd_index; // @[Core.scala 67:18]
  wire [63:0] rf_io_rd_data; // @[Core.scala 67:18]
  wire  rf_io_rd_wen; // @[Core.scala 67:18]
  wire  id_ex_clock; // @[Core.scala 74:35]
  wire  id_ex_reset; // @[Core.scala 74:35]
  wire  id_ex_io_in_uop_valid; // @[Core.scala 74:35]
  wire [2:0] id_ex_io_in_uop_exc; // @[Core.scala 74:35]
  wire [63:0] id_ex_io_in_uop_pc; // @[Core.scala 74:35]
  wire [63:0] id_ex_io_in_uop_npc; // @[Core.scala 74:35]
  wire [31:0] id_ex_io_in_uop_instr; // @[Core.scala 74:35]
  wire [2:0] id_ex_io_in_uop_fu; // @[Core.scala 74:35]
  wire [3:0] id_ex_io_in_uop_alu_op; // @[Core.scala 74:35]
  wire [1:0] id_ex_io_in_uop_jmp_op; // @[Core.scala 74:35]
  wire [3:0] id_ex_io_in_uop_mdu_op; // @[Core.scala 74:35]
  wire [4:0] id_ex_io_in_uop_lsu_op; // @[Core.scala 74:35]
  wire [1:0] id_ex_io_in_uop_mem_len; // @[Core.scala 74:35]
  wire [1:0] id_ex_io_in_uop_csr_op; // @[Core.scala 74:35]
  wire [2:0] id_ex_io_in_uop_sys_op; // @[Core.scala 74:35]
  wire [4:0] id_ex_io_in_uop_rd_index; // @[Core.scala 74:35]
  wire  id_ex_io_in_uop_rd_wen; // @[Core.scala 74:35]
  wire [31:0] id_ex_io_in_uop_imm; // @[Core.scala 74:35]
  wire  id_ex_io_in_uop_dw; // @[Core.scala 74:35]
  wire [63:0] id_ex_io_in_rs1_data; // @[Core.scala 74:35]
  wire [63:0] id_ex_io_in_rs2_data; // @[Core.scala 74:35]
  wire [63:0] id_ex_io_in_rs2_data_from_rf; // @[Core.scala 74:35]
  wire [63:0] id_ex_io_in_bp_npc; // @[Core.scala 74:35]
  wire  id_ex_io_out_uop_valid; // @[Core.scala 74:35]
  wire [2:0] id_ex_io_out_uop_exc; // @[Core.scala 74:35]
  wire [63:0] id_ex_io_out_uop_pc; // @[Core.scala 74:35]
  wire [63:0] id_ex_io_out_uop_npc; // @[Core.scala 74:35]
  wire [31:0] id_ex_io_out_uop_instr; // @[Core.scala 74:35]
  wire [2:0] id_ex_io_out_uop_fu; // @[Core.scala 74:35]
  wire [3:0] id_ex_io_out_uop_alu_op; // @[Core.scala 74:35]
  wire [1:0] id_ex_io_out_uop_jmp_op; // @[Core.scala 74:35]
  wire [3:0] id_ex_io_out_uop_mdu_op; // @[Core.scala 74:35]
  wire [4:0] id_ex_io_out_uop_lsu_op; // @[Core.scala 74:35]
  wire [1:0] id_ex_io_out_uop_mem_len; // @[Core.scala 74:35]
  wire [1:0] id_ex_io_out_uop_csr_op; // @[Core.scala 74:35]
  wire [2:0] id_ex_io_out_uop_sys_op; // @[Core.scala 74:35]
  wire [4:0] id_ex_io_out_uop_rd_index; // @[Core.scala 74:35]
  wire  id_ex_io_out_uop_rd_wen; // @[Core.scala 74:35]
  wire [31:0] id_ex_io_out_uop_imm; // @[Core.scala 74:35]
  wire  id_ex_io_out_uop_dw; // @[Core.scala 74:35]
  wire [63:0] id_ex_io_out_rs1_data; // @[Core.scala 74:35]
  wire [63:0] id_ex_io_out_rs2_data; // @[Core.scala 74:35]
  wire [63:0] id_ex_io_out_rs2_data_from_rf; // @[Core.scala 74:35]
  wire [63:0] id_ex_io_out_bp_npc; // @[Core.scala 74:35]
  wire  id_ex_io_en; // @[Core.scala 74:35]
  wire  id_ex_io_flush; // @[Core.scala 74:35]
  wire [3:0] alu_io_uop_alu_op; // @[Core.scala 85:19]
  wire [1:0] alu_io_uop_jmp_op; // @[Core.scala 85:19]
  wire  alu_io_uop_dw; // @[Core.scala 85:19]
  wire [63:0] alu_io_in1; // @[Core.scala 85:19]
  wire [63:0] alu_io_in2; // @[Core.scala 85:19]
  wire [63:0] alu_io_out; // @[Core.scala 85:19]
  wire [63:0] alu_io_adder_out; // @[Core.scala 85:19]
  wire  alu_io_cmp_out; // @[Core.scala 85:19]
  wire  lsu_clock; // @[Core.scala 108:19]
  wire  lsu_reset; // @[Core.scala 108:19]
  wire [4:0] lsu_io_uop_lsu_op; // @[Core.scala 108:19]
  wire [1:0] lsu_io_uop_mem_len; // @[Core.scala 108:19]
  wire  lsu_io_is_mem; // @[Core.scala 108:19]
  wire  lsu_io_is_store; // @[Core.scala 108:19]
  wire  lsu_io_is_amo; // @[Core.scala 108:19]
  wire [63:0] lsu_io_addr; // @[Core.scala 108:19]
  wire [63:0] lsu_io_wdata; // @[Core.scala 108:19]
  wire [63:0] lsu_io_rdata; // @[Core.scala 108:19]
  wire  lsu_io_valid; // @[Core.scala 108:19]
  wire [3:0] lsu_io_exc_code; // @[Core.scala 108:19]
  wire  lsu_io_dmem_req_ready; // @[Core.scala 108:19]
  wire  lsu_io_dmem_req_valid; // @[Core.scala 108:19]
  wire [38:0] lsu_io_dmem_req_bits_addr; // @[Core.scala 108:19]
  wire [63:0] lsu_io_dmem_req_bits_wdata; // @[Core.scala 108:19]
  wire [7:0] lsu_io_dmem_req_bits_wmask; // @[Core.scala 108:19]
  wire  lsu_io_dmem_req_bits_wen; // @[Core.scala 108:19]
  wire [1:0] lsu_io_dmem_req_bits_len; // @[Core.scala 108:19]
  wire  lsu_io_dmem_req_bits_lrsc; // @[Core.scala 108:19]
  wire [4:0] lsu_io_dmem_req_bits_amo; // @[Core.scala 108:19]
  wire  lsu_io_dmem_resp_ready; // @[Core.scala 108:19]
  wire  lsu_io_dmem_resp_valid; // @[Core.scala 108:19]
  wire [63:0] lsu_io_dmem_resp_bits_rdata; // @[Core.scala 108:19]
  wire  lsu_io_dmem_resp_bits_page_fault; // @[Core.scala 108:19]
  wire  lsu_io_dmem_resp_bits_access_fault; // @[Core.scala 108:19]
  wire  lsu_io_ready; // @[Core.scala 108:19]
  wire  mdu_clock; // @[Core.scala 116:19]
  wire  mdu_reset; // @[Core.scala 116:19]
  wire  mdu_io_uop_valid; // @[Core.scala 116:19]
  wire [3:0] mdu_io_uop_mdu_op; // @[Core.scala 116:19]
  wire  mdu_io_uop_dw; // @[Core.scala 116:19]
  wire  mdu_io_is_mdu; // @[Core.scala 116:19]
  wire [63:0] mdu_io_in1; // @[Core.scala 116:19]
  wire [63:0] mdu_io_in2; // @[Core.scala 116:19]
  wire [63:0] mdu_io_out; // @[Core.scala 116:19]
  wire  mdu_io_valid; // @[Core.scala 116:19]
  wire  mdu_io_ready; // @[Core.scala 116:19]
  wire  csr_clock; // @[Core.scala 122:19]
  wire  csr_reset; // @[Core.scala 122:19]
  wire  csr_io_uop_valid; // @[Core.scala 122:19]
  wire [2:0] csr_io_uop_exc; // @[Core.scala 122:19]
  wire [63:0] csr_io_uop_pc; // @[Core.scala 122:19]
  wire [63:0] csr_io_uop_npc; // @[Core.scala 122:19]
  wire [2:0] csr_io_uop_fu; // @[Core.scala 122:19]
  wire [2:0] csr_io_uop_sys_op; // @[Core.scala 122:19]
  wire [11:0] csr_io_rw_addr; // @[Core.scala 122:19]
  wire [1:0] csr_io_rw_cmd; // @[Core.scala 122:19]
  wire [63:0] csr_io_rw_wdata; // @[Core.scala 122:19]
  wire [63:0] csr_io_rw_rdata; // @[Core.scala 122:19]
  wire  csr_io_rw_valid; // @[Core.scala 122:19]
  wire [1:0] csr_io_prv; // @[Core.scala 122:19]
  wire  csr_io_mprv; // @[Core.scala 122:19]
  wire [1:0] csr_io_mpp; // @[Core.scala 122:19]
  wire  csr_io_sv39_en; // @[Core.scala 122:19]
  wire [15:0] csr_io_satp_asid; // @[Core.scala 122:19]
  wire [43:0] csr_io_satp_ppn; // @[Core.scala 122:19]
  wire  csr_io_sfence_vma; // @[Core.scala 122:19]
  wire  csr_io_fence_i; // @[Core.scala 122:19]
  wire  csr_io_jmp_packet_valid; // @[Core.scala 122:19]
  wire [63:0] csr_io_jmp_packet_target; // @[Core.scala 122:19]
  wire [63:0] csr_io_lsu_addr; // @[Core.scala 122:19]
  wire [3:0] csr_io_lsu_exc_code; // @[Core.scala 122:19]
  wire  csr_io_interrupt_mtip; // @[Core.scala 122:19]
  wire  csr_io_interrupt_msip; // @[Core.scala 122:19]
  wire  csr_io_interrupt_meip; // @[Core.scala 122:19]
  wire  csr_io_interrupt_seip; // @[Core.scala 122:19]
  wire  csr_io_is_int; // @[Core.scala 122:19]
  wire  csr_io_commit; // @[Core.scala 122:19]
  wire  dmem_proxy_clock; // @[Core.scala 142:26]
  wire  dmem_proxy_reset; // @[Core.scala 142:26]
  wire [1:0] dmem_proxy_io_prv; // @[Core.scala 142:26]
  wire  dmem_proxy_io_sv39_en; // @[Core.scala 142:26]
  wire [15:0] dmem_proxy_io_satp_asid; // @[Core.scala 142:26]
  wire [43:0] dmem_proxy_io_satp_ppn; // @[Core.scala 142:26]
  wire  dmem_proxy_io_sfence_vma; // @[Core.scala 142:26]
  wire  dmem_proxy_io_in_req_ready; // @[Core.scala 142:26]
  wire  dmem_proxy_io_in_req_valid; // @[Core.scala 142:26]
  wire [38:0] dmem_proxy_io_in_req_bits_addr; // @[Core.scala 142:26]
  wire [63:0] dmem_proxy_io_in_req_bits_wdata; // @[Core.scala 142:26]
  wire [7:0] dmem_proxy_io_in_req_bits_wmask; // @[Core.scala 142:26]
  wire  dmem_proxy_io_in_req_bits_wen; // @[Core.scala 142:26]
  wire [1:0] dmem_proxy_io_in_req_bits_len; // @[Core.scala 142:26]
  wire  dmem_proxy_io_in_req_bits_lrsc; // @[Core.scala 142:26]
  wire [4:0] dmem_proxy_io_in_req_bits_amo; // @[Core.scala 142:26]
  wire  dmem_proxy_io_in_resp_ready; // @[Core.scala 142:26]
  wire  dmem_proxy_io_in_resp_valid; // @[Core.scala 142:26]
  wire [63:0] dmem_proxy_io_in_resp_bits_rdata; // @[Core.scala 142:26]
  wire  dmem_proxy_io_in_resp_bits_page_fault; // @[Core.scala 142:26]
  wire  dmem_proxy_io_in_resp_bits_access_fault; // @[Core.scala 142:26]
  wire  dmem_proxy_io_out_req_ready; // @[Core.scala 142:26]
  wire  dmem_proxy_io_out_req_valid; // @[Core.scala 142:26]
  wire [38:0] dmem_proxy_io_out_req_bits_addr; // @[Core.scala 142:26]
  wire [63:0] dmem_proxy_io_out_req_bits_wdata; // @[Core.scala 142:26]
  wire [7:0] dmem_proxy_io_out_req_bits_wmask; // @[Core.scala 142:26]
  wire  dmem_proxy_io_out_req_bits_wen; // @[Core.scala 142:26]
  wire [1:0] dmem_proxy_io_out_req_bits_len; // @[Core.scala 142:26]
  wire  dmem_proxy_io_out_req_bits_lrsc; // @[Core.scala 142:26]
  wire [4:0] dmem_proxy_io_out_req_bits_amo; // @[Core.scala 142:26]
  wire  dmem_proxy_io_out_resp_ready; // @[Core.scala 142:26]
  wire  dmem_proxy_io_out_resp_valid; // @[Core.scala 142:26]
  wire [63:0] dmem_proxy_io_out_resp_bits_rdata; // @[Core.scala 142:26]
  wire  dmem_proxy_io_ptw_req_ready; // @[Core.scala 142:26]
  wire  dmem_proxy_io_ptw_req_valid; // @[Core.scala 142:26]
  wire [38:0] dmem_proxy_io_ptw_req_bits_addr; // @[Core.scala 142:26]
  wire  dmem_proxy_io_ptw_resp_ready; // @[Core.scala 142:26]
  wire  dmem_proxy_io_ptw_resp_valid; // @[Core.scala 142:26]
  wire [63:0] dmem_proxy_io_ptw_resp_bits_rdata; // @[Core.scala 142:26]
  wire  c2_xbar_clock; // @[Core.scala 164:23]
  wire  c2_xbar_reset; // @[Core.scala 164:23]
  wire  c2_xbar_io_in_req_ready; // @[Core.scala 164:23]
  wire  c2_xbar_io_in_req_valid; // @[Core.scala 164:23]
  wire [38:0] c2_xbar_io_in_req_bits_addr; // @[Core.scala 164:23]
  wire [63:0] c2_xbar_io_in_req_bits_wdata; // @[Core.scala 164:23]
  wire [7:0] c2_xbar_io_in_req_bits_wmask; // @[Core.scala 164:23]
  wire  c2_xbar_io_in_req_bits_wen; // @[Core.scala 164:23]
  wire [1:0] c2_xbar_io_in_req_bits_len; // @[Core.scala 164:23]
  wire  c2_xbar_io_in_req_bits_lrsc; // @[Core.scala 164:23]
  wire [4:0] c2_xbar_io_in_req_bits_amo; // @[Core.scala 164:23]
  wire  c2_xbar_io_in_resp_ready; // @[Core.scala 164:23]
  wire  c2_xbar_io_in_resp_valid; // @[Core.scala 164:23]
  wire [63:0] c2_xbar_io_in_resp_bits_rdata; // @[Core.scala 164:23]
  wire  c2_xbar_io_out_0_req_ready; // @[Core.scala 164:23]
  wire  c2_xbar_io_out_0_req_valid; // @[Core.scala 164:23]
  wire [38:0] c2_xbar_io_out_0_req_bits_addr; // @[Core.scala 164:23]
  wire [63:0] c2_xbar_io_out_0_req_bits_wdata; // @[Core.scala 164:23]
  wire [7:0] c2_xbar_io_out_0_req_bits_wmask; // @[Core.scala 164:23]
  wire  c2_xbar_io_out_0_req_bits_wen; // @[Core.scala 164:23]
  wire [1:0] c2_xbar_io_out_0_req_bits_len; // @[Core.scala 164:23]
  wire  c2_xbar_io_out_0_req_bits_lrsc; // @[Core.scala 164:23]
  wire [4:0] c2_xbar_io_out_0_req_bits_amo; // @[Core.scala 164:23]
  wire  c2_xbar_io_out_0_resp_ready; // @[Core.scala 164:23]
  wire  c2_xbar_io_out_0_resp_valid; // @[Core.scala 164:23]
  wire [63:0] c2_xbar_io_out_0_resp_bits_rdata; // @[Core.scala 164:23]
  wire  c2_xbar_io_out_1_req_ready; // @[Core.scala 164:23]
  wire  c2_xbar_io_out_1_req_valid; // @[Core.scala 164:23]
  wire [38:0] c2_xbar_io_out_1_req_bits_addr; // @[Core.scala 164:23]
  wire [63:0] c2_xbar_io_out_1_req_bits_wdata; // @[Core.scala 164:23]
  wire [7:0] c2_xbar_io_out_1_req_bits_wmask; // @[Core.scala 164:23]
  wire  c2_xbar_io_out_1_req_bits_wen; // @[Core.scala 164:23]
  wire [1:0] c2_xbar_io_out_1_req_bits_len; // @[Core.scala 164:23]
  wire  c2_xbar_io_out_1_resp_ready; // @[Core.scala 164:23]
  wire  c2_xbar_io_out_1_resp_valid; // @[Core.scala 164:23]
  wire [63:0] c2_xbar_io_out_1_resp_bits_rdata; // @[Core.scala 164:23]
  wire  c2_xbar_io_to_1; // @[Core.scala 164:23]
  wire  ex_wb_clock; // @[Core.scala 172:21]
  wire  ex_wb_reset; // @[Core.scala 172:21]
  wire  ex_wb_io_in_uop_valid; // @[Core.scala 172:21]
  wire [4:0] ex_wb_io_in_uop_rd_index; // @[Core.scala 172:21]
  wire  ex_wb_io_in_uop_rd_wen; // @[Core.scala 172:21]
  wire [63:0] ex_wb_io_in_rd_data; // @[Core.scala 172:21]
  wire  ex_wb_io_out_uop_valid; // @[Core.scala 172:21]
  wire [4:0] ex_wb_io_out_uop_rd_index; // @[Core.scala 172:21]
  wire  ex_wb_io_out_uop_rd_wen; // @[Core.scala 172:21]
  wire [63:0] ex_wb_io_out_rd_data; // @[Core.scala 172:21]
  wire  alu_jmp_packet_bp_update = id_ex_io_out_uop_valid & alu_io_uop_jmp_op != 2'h0; // @[Core.scala 96:54]
  wire  _alu_jmp_packet_target_T_5 = ~alu_io_uop_jmp_op[1] & alu_io_uop_jmp_op[0]; // @[Constant.scala 52:47]
  wire [31:0] _alu_jmp_packet_target_T_8 = id_ex_io_out_uop_imm[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _alu_jmp_packet_target_T_9 = {_alu_jmp_packet_target_T_8,id_ex_io_out_uop_imm}; // @[Cat.scala 33:92]
  wire [63:0] _alu_jmp_packet_target_T_11 = id_ex_io_out_uop_pc + _alu_jmp_packet_target_T_9; // @[Core.scala 93:45]
  wire [63:0] _alu_jmp_packet_target_T_12 = alu_io_cmp_out ? _alu_jmp_packet_target_T_11 : id_ex_io_out_uop_npc; // @[Core.scala 93:8]
  wire [63:0] alu_jmp_packet_target = _alu_jmp_packet_target_T_5 ? _alu_jmp_packet_target_T_12 : alu_io_adder_out; // @[Core.scala 91:31]
  wire  alu_jmp_packet_valid = alu_jmp_packet_bp_update & alu_jmp_packet_target != id_ex_io_out_bp_npc; // @[Core.scala 90:52]
  wire  sys_jmp_packet_valid = csr_io_jmp_packet_valid; // @[Core.scala 127:23 42:28]
  wire [63:0] sys_jmp_packet_target = csr_io_jmp_packet_target; // @[Core.scala 127:23 42:28]
  wire [63:0] alu_br_out = id_ex_io_out_uop_jmp_op[1] ? id_ex_io_out_uop_npc : alu_io_out; // @[Core.scala 100:23]
  wire  is_mem = id_ex_io_out_uop_fu == 3'h3 & id_ex_io_out_uop_valid; // @[Core.scala 102:58]
  wire  is_mdu = id_ex_io_out_uop_fu == 3'h2 & id_ex_io_out_uop_valid; // @[Core.scala 103:58]
  wire  is_csr = id_ex_io_out_uop_fu == 3'h4 & id_ex_io_out_uop_valid; // @[Core.scala 104:58]
  wire [1:0] prv = csr_io_prv; // @[Core.scala 128:23 19:24]
  wire  _ex_wb_io_in_uop_valid_T_3 = is_mdu & mdu_io_valid; // @[Core.scala 176:15]
  wire  _ex_wb_io_in_uop_valid_T_4 = is_mem & lsu_io_valid & lsu_io_exc_code == 4'h0 | _ex_wb_io_in_uop_valid_T_3; // @[Core.scala 175:59]
  wire  _ex_wb_io_in_uop_valid_T_5 = is_csr & csr_io_rw_valid; // @[Core.scala 177:15]
  wire  _ex_wb_io_in_uop_valid_T_6 = _ex_wb_io_in_uop_valid_T_4 | _ex_wb_io_in_uop_valid_T_5; // @[Core.scala 176:32]
  wire  _ex_wb_io_in_uop_valid_T_12 = ~is_mem & ~is_mdu & ~is_csr & id_ex_io_out_uop_valid; // @[Core.scala 178:38]
  wire  _ex_wb_io_in_uop_valid_T_13 = _ex_wb_io_in_uop_valid_T_6 | _ex_wb_io_in_uop_valid_T_12; // @[Core.scala 177:35]
  wire [63:0] _ex_wb_io_in_rd_data_T_1 = 3'h3 == id_ex_io_out_uop_fu ? lsu_io_rdata : alu_br_out; // @[Mux.scala 81:58]
  wire [63:0] _ex_wb_io_in_rd_data_T_3 = 3'h2 == id_ex_io_out_uop_fu ? mdu_io_out : _ex_wb_io_in_rd_data_T_1; // @[Mux.scala 81:58]
  wire  need_rs1 = decode_io_out_rs1_src == 2'h2; // @[Core.scala 202:40]
  wire  need_rs2 = decode_io_out_rs2_src == 2'h2; // @[Core.scala 203:40]
  wire  _need_rs2_from_rf_T_5 = ~decode_io_out_lsu_op[4] & decode_io_out_lsu_op[0]; // @[Constant.scala 82:45]
  wire  need_rs2_from_rf = _need_rs2_from_rf_T_5 | decode_io_out_lsu_op[4] | decode_io_out_fu == 3'h2; // @[Core.scala 205:66]
  wire  _T = need_rs1 & id_ex_io_out_uop_rd_wen; // @[Core.scala 208:14]
  wire  _T_2 = _T & decode_io_out_rs1_index == id_ex_io_out_uop_rd_index; // @[Core.scala 209:7]
  wire  _T_4 = _T_2 & decode_io_out_rs1_index != 5'h0; // @[Core.scala 210:7]
  wire [95:0] _id_rs1_data_T_1 = {32'h0,instr_buffer_io_deq_bits_pc}; // @[Cat.scala 33:92]
  wire [31:0] _id_rs1_data_T_4 = decode_io_out_imm[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _id_rs1_data_T_5 = {_id_rs1_data_T_4,decode_io_out_imm}; // @[Cat.scala 33:92]
  wire [95:0] _id_rs1_data_T_7 = 2'h1 == decode_io_out_rs1_src ? _id_rs1_data_T_1 : 96'h0; // @[Mux.scala 81:58]
  wire [95:0] _id_rs1_data_T_9 = 2'h2 == decode_io_out_rs1_src ? {{32'd0}, rf_io_rs1_data} : _id_rs1_data_T_7; // @[Mux.scala 81:58]
  wire [95:0] _id_rs1_data_T_11 = 2'h3 == decode_io_out_rs1_src ? {{32'd0}, _id_rs1_data_T_5} : _id_rs1_data_T_9; // @[Mux.scala 81:58]
  wire [95:0] _GEN_0 = _T_4 ? {{32'd0}, ex_wb_io_in_rd_data} : _id_rs1_data_T_11; // @[Core.scala 211:5 212:17 214:17]
  wire  _T_5 = need_rs2 & id_ex_io_out_uop_rd_wen; // @[Core.scala 226:14]
  wire  _T_6 = decode_io_out_rs2_index == id_ex_io_out_uop_rd_index; // @[Core.scala 227:34]
  wire  _T_7 = _T_5 & decode_io_out_rs2_index == id_ex_io_out_uop_rd_index; // @[Core.scala 227:7]
  wire  _T_8 = decode_io_out_rs2_index != 5'h0; // @[Core.scala 228:34]
  wire  _T_9 = _T_7 & decode_io_out_rs2_index != 5'h0; // @[Core.scala 228:7]
  wire [95:0] _id_rs2_data_T_7 = 2'h1 == decode_io_out_rs2_src ? _id_rs1_data_T_1 : 96'h0; // @[Mux.scala 81:58]
  wire [95:0] _id_rs2_data_T_9 = 2'h2 == decode_io_out_rs2_src ? {{32'd0}, rf_io_rs2_data} : _id_rs2_data_T_7; // @[Mux.scala 81:58]
  wire [95:0] _id_rs2_data_T_11 = 2'h3 == decode_io_out_rs2_src ? {{32'd0}, _id_rs1_data_T_5} : _id_rs2_data_T_9; // @[Mux.scala 81:58]
  wire [95:0] _GEN_1 = _T_9 ? {{32'd0}, ex_wb_io_in_rd_data} : _id_rs2_data_T_11; // @[Core.scala 229:5 230:17 232:17]
  wire  _T_10 = need_rs2_from_rf & id_ex_io_out_uop_rd_wen; // @[Core.scala 244:22]
  wire  _T_12 = _T_10 & _T_6; // @[Core.scala 245:7]
  wire  _T_14 = _T_12 & _T_8; // @[Core.scala 246:7]
  IFU ifu ( // @[Core.scala 27:19]
    .clock(ifu_clock),
    .reset(ifu_reset),
    .io_jmp_packet_valid(ifu_io_jmp_packet_valid),
    .io_jmp_packet_target(ifu_io_jmp_packet_target),
    .io_jmp_packet_bp_update(ifu_io_jmp_packet_bp_update),
    .io_jmp_packet_bp_taken(ifu_io_jmp_packet_bp_taken),
    .io_jmp_packet_bp_pc(ifu_io_jmp_packet_bp_pc),
    .io_imem_req_ready(ifu_io_imem_req_ready),
    .io_imem_req_valid(ifu_io_imem_req_valid),
    .io_imem_req_bits_addr(ifu_io_imem_req_bits_addr),
    .io_imem_resp_ready(ifu_io_imem_resp_ready),
    .io_imem_resp_valid(ifu_io_imem_resp_valid),
    .io_imem_resp_bits_rdata(ifu_io_imem_resp_bits_rdata),
    .io_imem_resp_bits_page_fault(ifu_io_imem_resp_bits_page_fault),
    .io_imem_resp_bits_access_fault(ifu_io_imem_resp_bits_access_fault),
    .io_out_pc(ifu_io_out_pc),
    .io_out_instr(ifu_io_out_instr),
    .io_out_valid(ifu_io_out_valid),
    .io_out_page_fault(ifu_io_out_page_fault),
    .io_out_access_fault(ifu_io_out_access_fault),
    .io_out_bp_npc(ifu_io_out_bp_npc),
    .io_stall_b(ifu_io_stall_b)
  );
  CachePortProxy imem_proxy ( // @[Core.scala 28:26]
    .clock(imem_proxy_clock),
    .reset(imem_proxy_reset),
    .io_prv(imem_proxy_io_prv),
    .io_sv39_en(imem_proxy_io_sv39_en),
    .io_satp_asid(imem_proxy_io_satp_asid),
    .io_satp_ppn(imem_proxy_io_satp_ppn),
    .io_sfence_vma(imem_proxy_io_sfence_vma),
    .io_in_req_ready(imem_proxy_io_in_req_ready),
    .io_in_req_valid(imem_proxy_io_in_req_valid),
    .io_in_req_bits_addr(imem_proxy_io_in_req_bits_addr),
    .io_in_resp_ready(imem_proxy_io_in_resp_ready),
    .io_in_resp_valid(imem_proxy_io_in_resp_valid),
    .io_in_resp_bits_rdata(imem_proxy_io_in_resp_bits_rdata),
    .io_in_resp_bits_page_fault(imem_proxy_io_in_resp_bits_page_fault),
    .io_in_resp_bits_access_fault(imem_proxy_io_in_resp_bits_access_fault),
    .io_out_req_ready(imem_proxy_io_out_req_ready),
    .io_out_req_valid(imem_proxy_io_out_req_valid),
    .io_out_req_bits_addr(imem_proxy_io_out_req_bits_addr),
    .io_out_resp_ready(imem_proxy_io_out_resp_ready),
    .io_out_resp_valid(imem_proxy_io_out_resp_valid),
    .io_out_resp_bits_rdata(imem_proxy_io_out_resp_bits_rdata),
    .io_ptw_req_ready(imem_proxy_io_ptw_req_ready),
    .io_ptw_req_valid(imem_proxy_io_ptw_req_valid),
    .io_ptw_req_bits_addr(imem_proxy_io_ptw_req_bits_addr),
    .io_ptw_resp_ready(imem_proxy_io_ptw_resp_ready),
    .io_ptw_resp_valid(imem_proxy_io_ptw_resp_valid),
    .io_ptw_resp_bits_rdata(imem_proxy_io_ptw_resp_bits_rdata)
  );
  Queue_2 instr_buffer ( // @[Core.scala 54:28]
    .clock(instr_buffer_clock),
    .reset(instr_buffer_reset),
    .io_enq_ready(instr_buffer_io_enq_ready),
    .io_enq_valid(instr_buffer_io_enq_valid),
    .io_enq_bits_pc(instr_buffer_io_enq_bits_pc),
    .io_enq_bits_instr(instr_buffer_io_enq_bits_instr),
    .io_enq_bits_page_fault(instr_buffer_io_enq_bits_page_fault),
    .io_enq_bits_access_fault(instr_buffer_io_enq_bits_access_fault),
    .io_enq_bits_bp_npc(instr_buffer_io_enq_bits_bp_npc),
    .io_deq_ready(instr_buffer_io_deq_ready),
    .io_deq_valid(instr_buffer_io_deq_valid),
    .io_deq_bits_pc(instr_buffer_io_deq_bits_pc),
    .io_deq_bits_instr(instr_buffer_io_deq_bits_instr),
    .io_deq_bits_page_fault(instr_buffer_io_deq_bits_page_fault),
    .io_deq_bits_access_fault(instr_buffer_io_deq_bits_access_fault),
    .io_deq_bits_bp_npc(instr_buffer_io_deq_bits_bp_npc),
    .io_flush(instr_buffer_io_flush)
  );
  Decode decode ( // @[Core.scala 63:22]
    .io_in_pc(decode_io_in_pc),
    .io_in_instr(decode_io_in_instr),
    .io_in_valid(decode_io_in_valid),
    .io_in_page_fault(decode_io_in_page_fault),
    .io_in_access_fault(decode_io_in_access_fault),
    .io_out_valid(decode_io_out_valid),
    .io_out_exc(decode_io_out_exc),
    .io_out_pc(decode_io_out_pc),
    .io_out_npc(decode_io_out_npc),
    .io_out_instr(decode_io_out_instr),
    .io_out_fu(decode_io_out_fu),
    .io_out_alu_op(decode_io_out_alu_op),
    .io_out_jmp_op(decode_io_out_jmp_op),
    .io_out_mdu_op(decode_io_out_mdu_op),
    .io_out_lsu_op(decode_io_out_lsu_op),
    .io_out_mem_len(decode_io_out_mem_len),
    .io_out_csr_op(decode_io_out_csr_op),
    .io_out_sys_op(decode_io_out_sys_op),
    .io_out_rs1_src(decode_io_out_rs1_src),
    .io_out_rs2_src(decode_io_out_rs2_src),
    .io_out_rs1_index(decode_io_out_rs1_index),
    .io_out_rs2_index(decode_io_out_rs2_index),
    .io_out_rd_index(decode_io_out_rd_index),
    .io_out_rd_wen(decode_io_out_rd_wen),
    .io_out_imm(decode_io_out_imm),
    .io_out_dw(decode_io_out_dw)
  );
  RegFile rf ( // @[Core.scala 67:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_rs1_index(rf_io_rs1_index),
    .io_rs2_index(rf_io_rs2_index),
    .io_rs1_data(rf_io_rs1_data),
    .io_rs2_data(rf_io_rs2_data),
    .io_rd_index(rf_io_rd_index),
    .io_rd_data(rf_io_rd_data),
    .io_rd_wen(rf_io_rd_wen)
  );
  PipelineReg id_ex ( // @[Core.scala 74:35]
    .clock(id_ex_clock),
    .reset(id_ex_reset),
    .io_in_uop_valid(id_ex_io_in_uop_valid),
    .io_in_uop_exc(id_ex_io_in_uop_exc),
    .io_in_uop_pc(id_ex_io_in_uop_pc),
    .io_in_uop_npc(id_ex_io_in_uop_npc),
    .io_in_uop_instr(id_ex_io_in_uop_instr),
    .io_in_uop_fu(id_ex_io_in_uop_fu),
    .io_in_uop_alu_op(id_ex_io_in_uop_alu_op),
    .io_in_uop_jmp_op(id_ex_io_in_uop_jmp_op),
    .io_in_uop_mdu_op(id_ex_io_in_uop_mdu_op),
    .io_in_uop_lsu_op(id_ex_io_in_uop_lsu_op),
    .io_in_uop_mem_len(id_ex_io_in_uop_mem_len),
    .io_in_uop_csr_op(id_ex_io_in_uop_csr_op),
    .io_in_uop_sys_op(id_ex_io_in_uop_sys_op),
    .io_in_uop_rd_index(id_ex_io_in_uop_rd_index),
    .io_in_uop_rd_wen(id_ex_io_in_uop_rd_wen),
    .io_in_uop_imm(id_ex_io_in_uop_imm),
    .io_in_uop_dw(id_ex_io_in_uop_dw),
    .io_in_rs1_data(id_ex_io_in_rs1_data),
    .io_in_rs2_data(id_ex_io_in_rs2_data),
    .io_in_rs2_data_from_rf(id_ex_io_in_rs2_data_from_rf),
    .io_in_bp_npc(id_ex_io_in_bp_npc),
    .io_out_uop_valid(id_ex_io_out_uop_valid),
    .io_out_uop_exc(id_ex_io_out_uop_exc),
    .io_out_uop_pc(id_ex_io_out_uop_pc),
    .io_out_uop_npc(id_ex_io_out_uop_npc),
    .io_out_uop_instr(id_ex_io_out_uop_instr),
    .io_out_uop_fu(id_ex_io_out_uop_fu),
    .io_out_uop_alu_op(id_ex_io_out_uop_alu_op),
    .io_out_uop_jmp_op(id_ex_io_out_uop_jmp_op),
    .io_out_uop_mdu_op(id_ex_io_out_uop_mdu_op),
    .io_out_uop_lsu_op(id_ex_io_out_uop_lsu_op),
    .io_out_uop_mem_len(id_ex_io_out_uop_mem_len),
    .io_out_uop_csr_op(id_ex_io_out_uop_csr_op),
    .io_out_uop_sys_op(id_ex_io_out_uop_sys_op),
    .io_out_uop_rd_index(id_ex_io_out_uop_rd_index),
    .io_out_uop_rd_wen(id_ex_io_out_uop_rd_wen),
    .io_out_uop_imm(id_ex_io_out_uop_imm),
    .io_out_uop_dw(id_ex_io_out_uop_dw),
    .io_out_rs1_data(id_ex_io_out_rs1_data),
    .io_out_rs2_data(id_ex_io_out_rs2_data),
    .io_out_rs2_data_from_rf(id_ex_io_out_rs2_data_from_rf),
    .io_out_bp_npc(id_ex_io_out_bp_npc),
    .io_en(id_ex_io_en),
    .io_flush(id_ex_io_flush)
  );
  ALU alu ( // @[Core.scala 85:19]
    .io_uop_alu_op(alu_io_uop_alu_op),
    .io_uop_jmp_op(alu_io_uop_jmp_op),
    .io_uop_dw(alu_io_uop_dw),
    .io_in1(alu_io_in1),
    .io_in2(alu_io_in2),
    .io_out(alu_io_out),
    .io_adder_out(alu_io_adder_out),
    .io_cmp_out(alu_io_cmp_out)
  );
  LSU lsu ( // @[Core.scala 108:19]
    .clock(lsu_clock),
    .reset(lsu_reset),
    .io_uop_lsu_op(lsu_io_uop_lsu_op),
    .io_uop_mem_len(lsu_io_uop_mem_len),
    .io_is_mem(lsu_io_is_mem),
    .io_is_store(lsu_io_is_store),
    .io_is_amo(lsu_io_is_amo),
    .io_addr(lsu_io_addr),
    .io_wdata(lsu_io_wdata),
    .io_rdata(lsu_io_rdata),
    .io_valid(lsu_io_valid),
    .io_exc_code(lsu_io_exc_code),
    .io_dmem_req_ready(lsu_io_dmem_req_ready),
    .io_dmem_req_valid(lsu_io_dmem_req_valid),
    .io_dmem_req_bits_addr(lsu_io_dmem_req_bits_addr),
    .io_dmem_req_bits_wdata(lsu_io_dmem_req_bits_wdata),
    .io_dmem_req_bits_wmask(lsu_io_dmem_req_bits_wmask),
    .io_dmem_req_bits_wen(lsu_io_dmem_req_bits_wen),
    .io_dmem_req_bits_len(lsu_io_dmem_req_bits_len),
    .io_dmem_req_bits_lrsc(lsu_io_dmem_req_bits_lrsc),
    .io_dmem_req_bits_amo(lsu_io_dmem_req_bits_amo),
    .io_dmem_resp_ready(lsu_io_dmem_resp_ready),
    .io_dmem_resp_valid(lsu_io_dmem_resp_valid),
    .io_dmem_resp_bits_rdata(lsu_io_dmem_resp_bits_rdata),
    .io_dmem_resp_bits_page_fault(lsu_io_dmem_resp_bits_page_fault),
    .io_dmem_resp_bits_access_fault(lsu_io_dmem_resp_bits_access_fault),
    .io_ready(lsu_io_ready)
  );
  MDU mdu ( // @[Core.scala 116:19]
    .clock(mdu_clock),
    .reset(mdu_reset),
    .io_uop_valid(mdu_io_uop_valid),
    .io_uop_mdu_op(mdu_io_uop_mdu_op),
    .io_uop_dw(mdu_io_uop_dw),
    .io_is_mdu(mdu_io_is_mdu),
    .io_in1(mdu_io_in1),
    .io_in2(mdu_io_in2),
    .io_out(mdu_io_out),
    .io_valid(mdu_io_valid),
    .io_ready(mdu_io_ready)
  );
  CSR csr ( // @[Core.scala 122:19]
    .clock(csr_clock),
    .reset(csr_reset),
    .io_uop_valid(csr_io_uop_valid),
    .io_uop_exc(csr_io_uop_exc),
    .io_uop_pc(csr_io_uop_pc),
    .io_uop_npc(csr_io_uop_npc),
    .io_uop_fu(csr_io_uop_fu),
    .io_uop_sys_op(csr_io_uop_sys_op),
    .io_rw_addr(csr_io_rw_addr),
    .io_rw_cmd(csr_io_rw_cmd),
    .io_rw_wdata(csr_io_rw_wdata),
    .io_rw_rdata(csr_io_rw_rdata),
    .io_rw_valid(csr_io_rw_valid),
    .io_prv(csr_io_prv),
    .io_mprv(csr_io_mprv),
    .io_mpp(csr_io_mpp),
    .io_sv39_en(csr_io_sv39_en),
    .io_satp_asid(csr_io_satp_asid),
    .io_satp_ppn(csr_io_satp_ppn),
    .io_sfence_vma(csr_io_sfence_vma),
    .io_fence_i(csr_io_fence_i),
    .io_jmp_packet_valid(csr_io_jmp_packet_valid),
    .io_jmp_packet_target(csr_io_jmp_packet_target),
    .io_lsu_addr(csr_io_lsu_addr),
    .io_lsu_exc_code(csr_io_lsu_exc_code),
    .io_interrupt_mtip(csr_io_interrupt_mtip),
    .io_interrupt_msip(csr_io_interrupt_msip),
    .io_interrupt_meip(csr_io_interrupt_meip),
    .io_interrupt_seip(csr_io_interrupt_seip),
    .io_is_int(csr_io_is_int),
    .io_commit(csr_io_commit)
  );
  CachePortProxy_1 dmem_proxy ( // @[Core.scala 142:26]
    .clock(dmem_proxy_clock),
    .reset(dmem_proxy_reset),
    .io_prv(dmem_proxy_io_prv),
    .io_sv39_en(dmem_proxy_io_sv39_en),
    .io_satp_asid(dmem_proxy_io_satp_asid),
    .io_satp_ppn(dmem_proxy_io_satp_ppn),
    .io_sfence_vma(dmem_proxy_io_sfence_vma),
    .io_in_req_ready(dmem_proxy_io_in_req_ready),
    .io_in_req_valid(dmem_proxy_io_in_req_valid),
    .io_in_req_bits_addr(dmem_proxy_io_in_req_bits_addr),
    .io_in_req_bits_wdata(dmem_proxy_io_in_req_bits_wdata),
    .io_in_req_bits_wmask(dmem_proxy_io_in_req_bits_wmask),
    .io_in_req_bits_wen(dmem_proxy_io_in_req_bits_wen),
    .io_in_req_bits_len(dmem_proxy_io_in_req_bits_len),
    .io_in_req_bits_lrsc(dmem_proxy_io_in_req_bits_lrsc),
    .io_in_req_bits_amo(dmem_proxy_io_in_req_bits_amo),
    .io_in_resp_ready(dmem_proxy_io_in_resp_ready),
    .io_in_resp_valid(dmem_proxy_io_in_resp_valid),
    .io_in_resp_bits_rdata(dmem_proxy_io_in_resp_bits_rdata),
    .io_in_resp_bits_page_fault(dmem_proxy_io_in_resp_bits_page_fault),
    .io_in_resp_bits_access_fault(dmem_proxy_io_in_resp_bits_access_fault),
    .io_out_req_ready(dmem_proxy_io_out_req_ready),
    .io_out_req_valid(dmem_proxy_io_out_req_valid),
    .io_out_req_bits_addr(dmem_proxy_io_out_req_bits_addr),
    .io_out_req_bits_wdata(dmem_proxy_io_out_req_bits_wdata),
    .io_out_req_bits_wmask(dmem_proxy_io_out_req_bits_wmask),
    .io_out_req_bits_wen(dmem_proxy_io_out_req_bits_wen),
    .io_out_req_bits_len(dmem_proxy_io_out_req_bits_len),
    .io_out_req_bits_lrsc(dmem_proxy_io_out_req_bits_lrsc),
    .io_out_req_bits_amo(dmem_proxy_io_out_req_bits_amo),
    .io_out_resp_ready(dmem_proxy_io_out_resp_ready),
    .io_out_resp_valid(dmem_proxy_io_out_resp_valid),
    .io_out_resp_bits_rdata(dmem_proxy_io_out_resp_bits_rdata),
    .io_ptw_req_ready(dmem_proxy_io_ptw_req_ready),
    .io_ptw_req_valid(dmem_proxy_io_ptw_req_valid),
    .io_ptw_req_bits_addr(dmem_proxy_io_ptw_req_bits_addr),
    .io_ptw_resp_ready(dmem_proxy_io_ptw_resp_ready),
    .io_ptw_resp_valid(dmem_proxy_io_ptw_resp_valid),
    .io_ptw_resp_bits_rdata(dmem_proxy_io_ptw_resp_bits_rdata)
  );
  CachePortXBar1to2 c2_xbar ( // @[Core.scala 164:23]
    .clock(c2_xbar_clock),
    .reset(c2_xbar_reset),
    .io_in_req_ready(c2_xbar_io_in_req_ready),
    .io_in_req_valid(c2_xbar_io_in_req_valid),
    .io_in_req_bits_addr(c2_xbar_io_in_req_bits_addr),
    .io_in_req_bits_wdata(c2_xbar_io_in_req_bits_wdata),
    .io_in_req_bits_wmask(c2_xbar_io_in_req_bits_wmask),
    .io_in_req_bits_wen(c2_xbar_io_in_req_bits_wen),
    .io_in_req_bits_len(c2_xbar_io_in_req_bits_len),
    .io_in_req_bits_lrsc(c2_xbar_io_in_req_bits_lrsc),
    .io_in_req_bits_amo(c2_xbar_io_in_req_bits_amo),
    .io_in_resp_ready(c2_xbar_io_in_resp_ready),
    .io_in_resp_valid(c2_xbar_io_in_resp_valid),
    .io_in_resp_bits_rdata(c2_xbar_io_in_resp_bits_rdata),
    .io_out_0_req_ready(c2_xbar_io_out_0_req_ready),
    .io_out_0_req_valid(c2_xbar_io_out_0_req_valid),
    .io_out_0_req_bits_addr(c2_xbar_io_out_0_req_bits_addr),
    .io_out_0_req_bits_wdata(c2_xbar_io_out_0_req_bits_wdata),
    .io_out_0_req_bits_wmask(c2_xbar_io_out_0_req_bits_wmask),
    .io_out_0_req_bits_wen(c2_xbar_io_out_0_req_bits_wen),
    .io_out_0_req_bits_len(c2_xbar_io_out_0_req_bits_len),
    .io_out_0_req_bits_lrsc(c2_xbar_io_out_0_req_bits_lrsc),
    .io_out_0_req_bits_amo(c2_xbar_io_out_0_req_bits_amo),
    .io_out_0_resp_ready(c2_xbar_io_out_0_resp_ready),
    .io_out_0_resp_valid(c2_xbar_io_out_0_resp_valid),
    .io_out_0_resp_bits_rdata(c2_xbar_io_out_0_resp_bits_rdata),
    .io_out_1_req_ready(c2_xbar_io_out_1_req_ready),
    .io_out_1_req_valid(c2_xbar_io_out_1_req_valid),
    .io_out_1_req_bits_addr(c2_xbar_io_out_1_req_bits_addr),
    .io_out_1_req_bits_wdata(c2_xbar_io_out_1_req_bits_wdata),
    .io_out_1_req_bits_wmask(c2_xbar_io_out_1_req_bits_wmask),
    .io_out_1_req_bits_wen(c2_xbar_io_out_1_req_bits_wen),
    .io_out_1_req_bits_len(c2_xbar_io_out_1_req_bits_len),
    .io_out_1_resp_ready(c2_xbar_io_out_1_resp_ready),
    .io_out_1_resp_valid(c2_xbar_io_out_1_resp_valid),
    .io_out_1_resp_bits_rdata(c2_xbar_io_out_1_resp_bits_rdata),
    .io_to_1(c2_xbar_io_to_1)
  );
  PipelineReg_1 ex_wb ( // @[Core.scala 172:21]
    .clock(ex_wb_clock),
    .reset(ex_wb_reset),
    .io_in_uop_valid(ex_wb_io_in_uop_valid),
    .io_in_uop_rd_index(ex_wb_io_in_uop_rd_index),
    .io_in_uop_rd_wen(ex_wb_io_in_uop_rd_wen),
    .io_in_rd_data(ex_wb_io_in_rd_data),
    .io_out_uop_valid(ex_wb_io_out_uop_valid),
    .io_out_uop_rd_index(ex_wb_io_out_uop_rd_index),
    .io_out_uop_rd_wen(ex_wb_io_out_uop_rd_wen),
    .io_out_rd_data(ex_wb_io_out_rd_data)
  );
  assign io_imem_req_valid = imem_proxy_io_out_req_valid; // @[Core.scala 33:28]
  assign io_imem_req_bits_addr = imem_proxy_io_out_req_bits_addr; // @[Core.scala 33:28]
  assign io_imem_resp_ready = imem_proxy_io_out_resp_ready; // @[Core.scala 33:28]
  assign io_dmem_req_valid = c2_xbar_io_out_0_req_valid; // @[Core.scala 169:20]
  assign io_dmem_req_bits_addr = c2_xbar_io_out_0_req_bits_addr; // @[Core.scala 169:20]
  assign io_dmem_req_bits_wdata = c2_xbar_io_out_0_req_bits_wdata; // @[Core.scala 169:20]
  assign io_dmem_req_bits_wmask = c2_xbar_io_out_0_req_bits_wmask; // @[Core.scala 169:20]
  assign io_dmem_req_bits_wen = c2_xbar_io_out_0_req_bits_wen; // @[Core.scala 169:20]
  assign io_dmem_req_bits_len = c2_xbar_io_out_0_req_bits_len; // @[Core.scala 169:20]
  assign io_dmem_req_bits_lrsc = c2_xbar_io_out_0_req_bits_lrsc; // @[Core.scala 169:20]
  assign io_dmem_req_bits_amo = c2_xbar_io_out_0_req_bits_amo; // @[Core.scala 169:20]
  assign io_dmem_resp_ready = c2_xbar_io_out_0_resp_ready; // @[Core.scala 169:20]
  assign io_iptw_req_valid = imem_proxy_io_ptw_req_valid; // @[Core.scala 34:28]
  assign io_iptw_req_bits_addr = imem_proxy_io_ptw_req_bits_addr; // @[Core.scala 34:28]
  assign io_iptw_resp_ready = imem_proxy_io_ptw_resp_ready; // @[Core.scala 34:28]
  assign io_dptw_req_valid = dmem_proxy_io_ptw_req_valid; // @[Core.scala 166:20]
  assign io_dptw_req_bits_addr = dmem_proxy_io_ptw_req_bits_addr; // @[Core.scala 166:20]
  assign io_dptw_resp_ready = dmem_proxy_io_ptw_resp_ready; // @[Core.scala 166:20]
  assign io_uncache_req_valid = c2_xbar_io_out_1_req_valid; // @[Core.scala 170:20]
  assign io_uncache_req_bits_addr = c2_xbar_io_out_1_req_bits_addr; // @[Core.scala 170:20]
  assign io_uncache_req_bits_wdata = c2_xbar_io_out_1_req_bits_wdata; // @[Core.scala 170:20]
  assign io_uncache_req_bits_wmask = c2_xbar_io_out_1_req_bits_wmask; // @[Core.scala 170:20]
  assign io_uncache_req_bits_wen = c2_xbar_io_out_1_req_bits_wen; // @[Core.scala 170:20]
  assign io_uncache_req_bits_len = c2_xbar_io_out_1_req_bits_len; // @[Core.scala 170:20]
  assign io_uncache_resp_ready = c2_xbar_io_out_1_resp_ready; // @[Core.scala 170:20]
  assign io_fence_i = csr_io_fence_i; // @[Core.scala 136:23]
  assign ifu_clock = clock;
  assign ifu_reset = reset;
  assign ifu_io_jmp_packet_valid = alu_jmp_packet_valid | sys_jmp_packet_valid; // @[Core.scala 43:55]
  assign ifu_io_jmp_packet_target = sys_jmp_packet_valid ? sys_jmp_packet_target : alu_jmp_packet_target; // @[Core.scala 44:37]
  assign ifu_io_jmp_packet_bp_update = id_ex_io_out_uop_valid & alu_io_uop_jmp_op != 2'h0; // @[Core.scala 96:54]
  assign ifu_io_jmp_packet_bp_taken = _alu_jmp_packet_target_T_5 ? alu_io_cmp_out : alu_io_uop_jmp_op[1]; // @[Core.scala 97:34]
  assign ifu_io_jmp_packet_bp_pc = id_ex_io_out_uop_pc; // @[Core.scala 41:28 98:28]
  assign ifu_io_imem_req_ready = imem_proxy_io_in_req_ready; // @[Core.scala 32:28]
  assign ifu_io_imem_resp_valid = imem_proxy_io_in_resp_valid; // @[Core.scala 32:28]
  assign ifu_io_imem_resp_bits_rdata = imem_proxy_io_in_resp_bits_rdata; // @[Core.scala 32:28]
  assign ifu_io_imem_resp_bits_page_fault = imem_proxy_io_in_resp_bits_page_fault; // @[Core.scala 32:28]
  assign ifu_io_imem_resp_bits_access_fault = imem_proxy_io_in_resp_bits_access_fault; // @[Core.scala 32:28]
  assign ifu_io_stall_b = instr_buffer_io_enq_ready; // @[Core.scala 55:29]
  assign imem_proxy_clock = clock;
  assign imem_proxy_reset = reset;
  assign imem_proxy_io_prv = csr_io_prv; // @[Core.scala 128:23 19:24]
  assign imem_proxy_io_sv39_en = csr_io_sv39_en; // @[Core.scala 129:23 20:24]
  assign imem_proxy_io_satp_asid = csr_io_satp_asid; // @[Core.scala 130:23 21:24]
  assign imem_proxy_io_satp_ppn = csr_io_satp_ppn; // @[Core.scala 131:23 22:24]
  assign imem_proxy_io_sfence_vma = csr_io_sfence_vma; // @[Core.scala 132:23 23:24]
  assign imem_proxy_io_in_req_valid = ifu_io_imem_req_valid; // @[Core.scala 32:28]
  assign imem_proxy_io_in_req_bits_addr = ifu_io_imem_req_bits_addr; // @[Core.scala 32:28]
  assign imem_proxy_io_in_resp_ready = ifu_io_imem_resp_ready; // @[Core.scala 32:28]
  assign imem_proxy_io_out_req_ready = io_imem_req_ready; // @[Core.scala 33:28]
  assign imem_proxy_io_out_resp_valid = io_imem_resp_valid; // @[Core.scala 33:28]
  assign imem_proxy_io_out_resp_bits_rdata = io_imem_resp_bits_rdata; // @[Core.scala 33:28]
  assign imem_proxy_io_ptw_req_ready = io_iptw_req_ready; // @[Core.scala 34:28]
  assign imem_proxy_io_ptw_resp_valid = io_iptw_resp_valid; // @[Core.scala 34:28]
  assign imem_proxy_io_ptw_resp_bits_rdata = io_iptw_resp_bits_rdata; // @[Core.scala 34:28]
  assign instr_buffer_clock = clock;
  assign instr_buffer_reset = reset;
  assign instr_buffer_io_enq_valid = ifu_io_out_valid; // @[Core.scala 57:29]
  assign instr_buffer_io_enq_bits_pc = ifu_io_out_pc; // @[Core.scala 56:29]
  assign instr_buffer_io_enq_bits_instr = ifu_io_out_instr; // @[Core.scala 56:29]
  assign instr_buffer_io_enq_bits_page_fault = ifu_io_out_page_fault; // @[Core.scala 56:29]
  assign instr_buffer_io_enq_bits_access_fault = ifu_io_out_access_fault; // @[Core.scala 56:29]
  assign instr_buffer_io_enq_bits_bp_npc = ifu_io_out_bp_npc; // @[Core.scala 56:29]
  assign instr_buffer_io_deq_ready = lsu_io_ready & mdu_io_ready; // @[Core.scala 255:27]
  assign instr_buffer_io_flush = alu_jmp_packet_valid | sys_jmp_packet_valid; // @[Core.scala 256:35]
  assign decode_io_in_pc = instr_buffer_io_deq_bits_pc; // @[Core.scala 64:22]
  assign decode_io_in_instr = instr_buffer_io_deq_bits_instr; // @[Core.scala 64:22]
  assign decode_io_in_valid = instr_buffer_io_deq_ready & instr_buffer_io_deq_valid; // @[Decoupled.scala 51:35]
  assign decode_io_in_page_fault = instr_buffer_io_deq_bits_page_fault; // @[Core.scala 64:22]
  assign decode_io_in_access_fault = instr_buffer_io_deq_bits_access_fault; // @[Core.scala 64:22]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_rs1_index = decode_io_out_rs1_index; // @[Core.scala 68:19]
  assign rf_io_rs2_index = decode_io_out_rs2_index; // @[Core.scala 69:19]
  assign rf_io_rd_index = ex_wb_io_out_uop_rd_index; // @[Core.scala 197:18]
  assign rf_io_rd_data = ex_wb_io_out_rd_data; // @[Core.scala 198:18]
  assign rf_io_rd_wen = ex_wb_io_out_uop_valid & ex_wb_io_out_uop_rd_wen; // @[Core.scala 196:38]
  assign id_ex_clock = clock;
  assign id_ex_reset = reset;
  assign id_ex_io_in_uop_valid = decode_io_out_valid; // @[Core.scala 75:32]
  assign id_ex_io_in_uop_exc = decode_io_out_exc; // @[Core.scala 75:32]
  assign id_ex_io_in_uop_pc = decode_io_out_pc; // @[Core.scala 75:32]
  assign id_ex_io_in_uop_npc = decode_io_out_npc; // @[Core.scala 75:32]
  assign id_ex_io_in_uop_instr = decode_io_out_instr; // @[Core.scala 75:32]
  assign id_ex_io_in_uop_fu = decode_io_out_fu; // @[Core.scala 75:32]
  assign id_ex_io_in_uop_alu_op = decode_io_out_alu_op; // @[Core.scala 75:32]
  assign id_ex_io_in_uop_jmp_op = decode_io_out_jmp_op; // @[Core.scala 75:32]
  assign id_ex_io_in_uop_mdu_op = decode_io_out_mdu_op; // @[Core.scala 75:32]
  assign id_ex_io_in_uop_lsu_op = decode_io_out_lsu_op; // @[Core.scala 75:32]
  assign id_ex_io_in_uop_mem_len = decode_io_out_mem_len; // @[Core.scala 75:32]
  assign id_ex_io_in_uop_csr_op = decode_io_out_csr_op; // @[Core.scala 75:32]
  assign id_ex_io_in_uop_sys_op = decode_io_out_sys_op; // @[Core.scala 75:32]
  assign id_ex_io_in_uop_rd_index = decode_io_out_rd_index; // @[Core.scala 75:32]
  assign id_ex_io_in_uop_rd_wen = decode_io_out_rd_wen; // @[Core.scala 75:32]
  assign id_ex_io_in_uop_imm = decode_io_out_imm; // @[Core.scala 75:32]
  assign id_ex_io_in_uop_dw = decode_io_out_dw; // @[Core.scala 75:32]
  assign id_ex_io_in_rs1_data = _GEN_0[63:0]; // @[Core.scala 71:33]
  assign id_ex_io_in_rs2_data = _GEN_1[63:0]; // @[Core.scala 72:33]
  assign id_ex_io_in_rs2_data_from_rf = _T_14 ? ex_wb_io_in_rd_data : rf_io_rs2_data; // @[Core.scala 247:5 248:25 250:25]
  assign id_ex_io_in_bp_npc = instr_buffer_io_deq_bits_bp_npc; // @[Core.scala 79:32]
  assign id_ex_io_en = lsu_io_ready & mdu_io_ready; // @[Core.scala 255:27]
  assign id_ex_io_flush = alu_jmp_packet_valid | sys_jmp_packet_valid; // @[Core.scala 256:35]
  assign alu_io_uop_alu_op = id_ex_io_out_uop_alu_op; // @[Core.scala 86:14]
  assign alu_io_uop_jmp_op = id_ex_io_out_uop_jmp_op; // @[Core.scala 86:14]
  assign alu_io_uop_dw = id_ex_io_out_uop_dw; // @[Core.scala 86:14]
  assign alu_io_in1 = id_ex_io_out_rs1_data; // @[Core.scala 87:14]
  assign alu_io_in2 = id_ex_io_out_rs2_data; // @[Core.scala 88:14]
  assign lsu_clock = clock;
  assign lsu_reset = reset;
  assign lsu_io_uop_lsu_op = id_ex_io_out_uop_lsu_op; // @[Core.scala 109:19]
  assign lsu_io_uop_mem_len = id_ex_io_out_uop_mem_len; // @[Core.scala 109:19]
  assign lsu_io_is_mem = id_ex_io_out_uop_fu == 3'h3 & id_ex_io_out_uop_valid; // @[Core.scala 102:58]
  assign lsu_io_is_store = ~id_ex_io_out_uop_lsu_op[4] & id_ex_io_out_uop_lsu_op[0]; // @[Constant.scala 82:45]
  assign lsu_io_is_amo = id_ex_io_out_uop_lsu_op[4]; // @[Constant.scala 81:33]
  assign lsu_io_addr = id_ex_io_out_uop_jmp_op[1] ? id_ex_io_out_uop_npc : alu_io_out; // @[Core.scala 100:23]
  assign lsu_io_wdata = id_ex_io_out_rs2_data_from_rf; // @[Core.scala 114:19]
  assign lsu_io_dmem_req_ready = dmem_proxy_io_in_req_ready; // @[Core.scala 165:20]
  assign lsu_io_dmem_resp_valid = dmem_proxy_io_in_resp_valid; // @[Core.scala 165:20]
  assign lsu_io_dmem_resp_bits_rdata = dmem_proxy_io_in_resp_bits_rdata; // @[Core.scala 165:20]
  assign lsu_io_dmem_resp_bits_page_fault = dmem_proxy_io_in_resp_bits_page_fault; // @[Core.scala 165:20]
  assign lsu_io_dmem_resp_bits_access_fault = dmem_proxy_io_in_resp_bits_access_fault; // @[Core.scala 165:20]
  assign mdu_clock = clock;
  assign mdu_reset = reset;
  assign mdu_io_uop_valid = id_ex_io_out_uop_valid; // @[Core.scala 117:17]
  assign mdu_io_uop_mdu_op = id_ex_io_out_uop_mdu_op; // @[Core.scala 117:17]
  assign mdu_io_uop_dw = id_ex_io_out_uop_dw; // @[Core.scala 117:17]
  assign mdu_io_is_mdu = id_ex_io_out_uop_fu == 3'h2 & id_ex_io_out_uop_valid; // @[Core.scala 103:58]
  assign mdu_io_in1 = id_ex_io_out_rs1_data; // @[Core.scala 119:17]
  assign mdu_io_in2 = id_ex_io_out_rs2_data_from_rf; // @[Core.scala 120:17]
  assign csr_clock = clock;
  assign csr_reset = reset;
  assign csr_io_uop_valid = id_ex_io_out_uop_valid; // @[Core.scala 123:23]
  assign csr_io_uop_exc = id_ex_io_out_uop_exc; // @[Core.scala 123:23]
  assign csr_io_uop_pc = id_ex_io_out_uop_pc; // @[Core.scala 123:23]
  assign csr_io_uop_npc = id_ex_io_out_uop_npc; // @[Core.scala 123:23]
  assign csr_io_uop_fu = id_ex_io_out_uop_fu; // @[Core.scala 123:23]
  assign csr_io_uop_sys_op = id_ex_io_out_uop_sys_op; // @[Core.scala 123:23]
  assign csr_io_rw_addr = id_ex_io_out_uop_instr[31:20]; // @[Core.scala 124:48]
  assign csr_io_rw_cmd = id_ex_io_out_uop_csr_op; // @[Core.scala 125:23]
  assign csr_io_rw_wdata = id_ex_io_out_rs1_data; // @[Core.scala 126:23]
  assign csr_io_lsu_addr = lsu_io_addr; // @[Core.scala 133:23]
  assign csr_io_lsu_exc_code = lsu_io_exc_code; // @[Core.scala 134:23]
  assign csr_io_interrupt_mtip = io_intr_mtip; // @[Core.scala 135:23]
  assign csr_io_interrupt_msip = io_intr_msip; // @[Core.scala 135:23]
  assign csr_io_interrupt_meip = io_intr_meip; // @[Core.scala 135:23]
  assign csr_io_interrupt_seip = io_intr_seip; // @[Core.scala 135:23]
  assign csr_io_commit = ex_wb_io_out_uop_valid; // @[Core.scala 262:17]
  assign dmem_proxy_clock = clock;
  assign dmem_proxy_reset = reset;
  assign dmem_proxy_io_prv = csr_io_mprv ? csr_io_mpp : prv; // @[Core.scala 146:34]
  assign dmem_proxy_io_sv39_en = csr_io_sv39_en; // @[Core.scala 129:23 20:24]
  assign dmem_proxy_io_satp_asid = csr_io_satp_asid; // @[Core.scala 130:23 21:24]
  assign dmem_proxy_io_satp_ppn = csr_io_satp_ppn; // @[Core.scala 131:23 22:24]
  assign dmem_proxy_io_sfence_vma = csr_io_sfence_vma; // @[Core.scala 132:23 23:24]
  assign dmem_proxy_io_in_req_valid = lsu_io_dmem_req_valid; // @[Core.scala 165:20]
  assign dmem_proxy_io_in_req_bits_addr = lsu_io_dmem_req_bits_addr; // @[Core.scala 165:20]
  assign dmem_proxy_io_in_req_bits_wdata = lsu_io_dmem_req_bits_wdata; // @[Core.scala 165:20]
  assign dmem_proxy_io_in_req_bits_wmask = lsu_io_dmem_req_bits_wmask; // @[Core.scala 165:20]
  assign dmem_proxy_io_in_req_bits_wen = lsu_io_dmem_req_bits_wen; // @[Core.scala 165:20]
  assign dmem_proxy_io_in_req_bits_len = lsu_io_dmem_req_bits_len; // @[Core.scala 165:20]
  assign dmem_proxy_io_in_req_bits_lrsc = lsu_io_dmem_req_bits_lrsc; // @[Core.scala 165:20]
  assign dmem_proxy_io_in_req_bits_amo = lsu_io_dmem_req_bits_amo; // @[Core.scala 165:20]
  assign dmem_proxy_io_in_resp_ready = lsu_io_dmem_resp_ready; // @[Core.scala 165:20]
  assign dmem_proxy_io_out_req_ready = c2_xbar_io_in_req_ready; // @[Core.scala 167:20]
  assign dmem_proxy_io_out_resp_valid = c2_xbar_io_in_resp_valid; // @[Core.scala 167:20]
  assign dmem_proxy_io_out_resp_bits_rdata = c2_xbar_io_in_resp_bits_rdata; // @[Core.scala 167:20]
  assign dmem_proxy_io_ptw_req_ready = io_dptw_req_ready; // @[Core.scala 166:20]
  assign dmem_proxy_io_ptw_resp_valid = io_dptw_resp_valid; // @[Core.scala 166:20]
  assign dmem_proxy_io_ptw_resp_bits_rdata = io_dptw_resp_bits_rdata; // @[Core.scala 166:20]
  assign c2_xbar_clock = clock;
  assign c2_xbar_reset = reset;
  assign c2_xbar_io_in_req_valid = dmem_proxy_io_out_req_valid; // @[Core.scala 167:20]
  assign c2_xbar_io_in_req_bits_addr = dmem_proxy_io_out_req_bits_addr; // @[Core.scala 167:20]
  assign c2_xbar_io_in_req_bits_wdata = dmem_proxy_io_out_req_bits_wdata; // @[Core.scala 167:20]
  assign c2_xbar_io_in_req_bits_wmask = dmem_proxy_io_out_req_bits_wmask; // @[Core.scala 167:20]
  assign c2_xbar_io_in_req_bits_wen = dmem_proxy_io_out_req_bits_wen; // @[Core.scala 167:20]
  assign c2_xbar_io_in_req_bits_len = dmem_proxy_io_out_req_bits_len; // @[Core.scala 167:20]
  assign c2_xbar_io_in_req_bits_lrsc = dmem_proxy_io_out_req_bits_lrsc; // @[Core.scala 167:20]
  assign c2_xbar_io_in_req_bits_amo = dmem_proxy_io_out_req_bits_amo; // @[Core.scala 167:20]
  assign c2_xbar_io_in_resp_ready = dmem_proxy_io_out_resp_ready; // @[Core.scala 167:20]
  assign c2_xbar_io_out_0_req_ready = io_dmem_req_ready; // @[Core.scala 169:20]
  assign c2_xbar_io_out_0_resp_valid = io_dmem_resp_valid; // @[Core.scala 169:20]
  assign c2_xbar_io_out_0_resp_bits_rdata = io_dmem_resp_bits_rdata; // @[Core.scala 169:20]
  assign c2_xbar_io_out_1_req_ready = io_uncache_req_ready; // @[Core.scala 170:20]
  assign c2_xbar_io_out_1_resp_valid = io_uncache_resp_valid; // @[Core.scala 170:20]
  assign c2_xbar_io_out_1_resp_bits_rdata = io_uncache_resp_bits_rdata; // @[Core.scala 170:20]
  assign c2_xbar_io_to_1 = ~dmem_proxy_io_out_req_bits_addr[31]; // @[Core.scala 168:23]
  assign ex_wb_clock = clock;
  assign ex_wb_reset = reset;
  assign ex_wb_io_in_uop_valid = _ex_wb_io_in_uop_valid_T_13 & ~csr_io_is_int; // @[Core.scala 179:5]
  assign ex_wb_io_in_uop_rd_index = id_ex_io_out_uop_rd_index; // @[Core.scala 173:19]
  assign ex_wb_io_in_uop_rd_wen = id_ex_io_out_uop_rd_wen; // @[Core.scala 173:19]
  assign ex_wb_io_in_rd_data = 3'h4 == id_ex_io_out_uop_fu ? csr_io_rw_rdata : _ex_wb_io_in_rd_data_T_3; // @[Mux.scala 81:58]
endmodule
module RRArbiter(
  input         clock,
  input         io_in_0_valid,
  input  [38:0] io_in_0_bits_addr,
  input  [63:0] io_in_0_bits_wdata,
  input  [7:0]  io_in_0_bits_wmask,
  input         io_in_0_bits_wen,
  input  [1:0]  io_in_0_bits_len,
  input         io_in_0_bits_lrsc,
  input  [4:0]  io_in_0_bits_amo,
  input         io_in_1_valid,
  input  [38:0] io_in_1_bits_addr,
  input         io_in_2_valid,
  input  [38:0] io_in_2_bits_addr,
  input         io_out_ready,
  output        io_out_valid,
  output [38:0] io_out_bits_addr,
  output [63:0] io_out_bits_wdata,
  output [7:0]  io_out_bits_wmask,
  output        io_out_bits_wen,
  output [1:0]  io_out_bits_len,
  output        io_out_bits_lrsc,
  output [4:0]  io_out_bits_amo,
  output [1:0]  io_chosen
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  _GEN_1 = 2'h1 == io_chosen ? io_in_1_valid : io_in_0_valid; // @[Arbiter.scala 55:{16,16}]
  wire [38:0] _GEN_4 = 2'h1 == io_chosen ? io_in_1_bits_addr : io_in_0_bits_addr; // @[Arbiter.scala 56:{15,15}]
  wire [63:0] _GEN_7 = 2'h1 == io_chosen ? 64'h0 : io_in_0_bits_wdata; // @[Arbiter.scala 56:{15,15}]
  wire [7:0] _GEN_10 = 2'h1 == io_chosen ? 8'h0 : io_in_0_bits_wmask; // @[Arbiter.scala 56:{15,15}]
  wire  _GEN_13 = 2'h1 == io_chosen ? 1'h0 : io_in_0_bits_wen; // @[Arbiter.scala 56:{15,15}]
  wire [1:0] _GEN_16 = 2'h1 == io_chosen ? 2'h0 : io_in_0_bits_len; // @[Arbiter.scala 56:{15,15}]
  wire  _GEN_19 = 2'h1 == io_chosen ? 1'h0 : io_in_0_bits_lrsc; // @[Arbiter.scala 56:{15,15}]
  wire [4:0] _GEN_22 = 2'h1 == io_chosen ? 5'h0 : io_in_0_bits_amo; // @[Arbiter.scala 56:{15,15}]
  wire  _ctrl_validMask_grantMask_lastGrant_T = io_out_ready & io_out_valid; // @[Decoupled.scala 51:35]
  reg [1:0] lastGrant; // @[Reg.scala 19:16]
  wire  grantMask_1 = 2'h1 > lastGrant; // @[Arbiter.scala 81:49]
  wire  grantMask_2 = 2'h2 > lastGrant; // @[Arbiter.scala 81:49]
  wire  validMask_1 = io_in_1_valid & grantMask_1; // @[Arbiter.scala 82:76]
  wire  validMask_2 = io_in_2_valid & grantMask_2; // @[Arbiter.scala 82:76]
  wire [1:0] _GEN_25 = io_in_1_valid ? 2'h1 : 2'h2; // @[Arbiter.scala 91:{26,35} 89:41]
  wire [1:0] _GEN_26 = io_in_0_valid ? 2'h0 : _GEN_25; // @[Arbiter.scala 91:{26,35}]
  wire [1:0] _GEN_27 = validMask_2 ? 2'h2 : _GEN_26; // @[Arbiter.scala 93:{24,33}]
  assign io_out_valid = 2'h2 == io_chosen ? io_in_2_valid : _GEN_1; // @[Arbiter.scala 55:{16,16}]
  assign io_out_bits_addr = 2'h2 == io_chosen ? io_in_2_bits_addr : _GEN_4; // @[Arbiter.scala 56:{15,15}]
  assign io_out_bits_wdata = 2'h2 == io_chosen ? 64'h0 : _GEN_7; // @[Arbiter.scala 56:{15,15}]
  assign io_out_bits_wmask = 2'h2 == io_chosen ? 8'h0 : _GEN_10; // @[Arbiter.scala 56:{15,15}]
  assign io_out_bits_wen = 2'h2 == io_chosen ? 1'h0 : _GEN_13; // @[Arbiter.scala 56:{15,15}]
  assign io_out_bits_len = 2'h2 == io_chosen ? 2'h0 : _GEN_16; // @[Arbiter.scala 56:{15,15}]
  assign io_out_bits_lrsc = 2'h2 == io_chosen ? 1'h0 : _GEN_19; // @[Arbiter.scala 56:{15,15}]
  assign io_out_bits_amo = 2'h2 == io_chosen ? 5'h0 : _GEN_22; // @[Arbiter.scala 56:{15,15}]
  assign io_chosen = validMask_1 ? 2'h1 : _GEN_27; // @[Arbiter.scala 93:{24,33}]
  always @(posedge clock) begin
    if (_ctrl_validMask_grantMask_lastGrant_T) begin // @[Reg.scala 20:18]
      lastGrant <= io_chosen; // @[Reg.scala 20:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lastGrant = _RAND_0[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_3(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [1:0] io_enq_bits,
  input        io_deq_ready,
  output       io_deq_valid,
  output [1:0] io_deq_bits
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] ram [0:3]; // @[Decoupled.scala 273:95]
  wire  ram_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire [1:0] ram_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [1:0] ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_MPORT_en; // @[Decoupled.scala 273:95]
  reg [1:0] enq_ptr_value; // @[Counter.scala 61:40]
  reg [1:0] deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _value_T_1 = enq_ptr_value + 2'h1; // @[Counter.scala 77:24]
  wire [1:0] _value_T_3 = deq_ptr_value + 2'h1; // @[Counter.scala 77:24]
  assign ram_io_deq_bits_MPORT_en = 1'h1;
  assign ram_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_MPORT_data = io_enq_bits;
  assign ram_MPORT_addr = enq_ptr_value;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits = ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  always @(posedge clock) begin
    if (ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 2'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 2'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram[initvar] = _RAND_0[1:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enq_ptr_value = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  deq_ptr_value = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CachePortXBarNto1(
  input         clock,
  input         reset,
  output        io_in_0_req_ready,
  input         io_in_0_req_valid,
  input  [38:0] io_in_0_req_bits_addr,
  input  [63:0] io_in_0_req_bits_wdata,
  input  [7:0]  io_in_0_req_bits_wmask,
  input         io_in_0_req_bits_wen,
  input  [1:0]  io_in_0_req_bits_len,
  input         io_in_0_req_bits_lrsc,
  input  [4:0]  io_in_0_req_bits_amo,
  input         io_in_0_resp_ready,
  output        io_in_0_resp_valid,
  output [63:0] io_in_0_resp_bits_rdata,
  output        io_in_1_req_ready,
  input         io_in_1_req_valid,
  input  [38:0] io_in_1_req_bits_addr,
  input         io_in_1_resp_ready,
  output        io_in_1_resp_valid,
  output [63:0] io_in_1_resp_bits_rdata,
  output        io_in_2_req_ready,
  input         io_in_2_req_valid,
  input  [38:0] io_in_2_req_bits_addr,
  input         io_in_2_resp_ready,
  output        io_in_2_resp_valid,
  output [63:0] io_in_2_resp_bits_rdata,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [38:0] io_out_req_bits_addr,
  output [63:0] io_out_req_bits_wdata,
  output [7:0]  io_out_req_bits_wmask,
  output        io_out_req_bits_wen,
  output [1:0]  io_out_req_bits_len,
  output        io_out_req_bits_lrsc,
  output [4:0]  io_out_req_bits_amo,
  output        io_out_resp_ready,
  input         io_out_resp_valid,
  input  [63:0] io_out_resp_bits_rdata
);
  wire  arbiter_clock; // @[Bus.scala 47:23]
  wire  arbiter_io_in_0_valid; // @[Bus.scala 47:23]
  wire [38:0] arbiter_io_in_0_bits_addr; // @[Bus.scala 47:23]
  wire [63:0] arbiter_io_in_0_bits_wdata; // @[Bus.scala 47:23]
  wire [7:0] arbiter_io_in_0_bits_wmask; // @[Bus.scala 47:23]
  wire  arbiter_io_in_0_bits_wen; // @[Bus.scala 47:23]
  wire [1:0] arbiter_io_in_0_bits_len; // @[Bus.scala 47:23]
  wire  arbiter_io_in_0_bits_lrsc; // @[Bus.scala 47:23]
  wire [4:0] arbiter_io_in_0_bits_amo; // @[Bus.scala 47:23]
  wire  arbiter_io_in_1_valid; // @[Bus.scala 47:23]
  wire [38:0] arbiter_io_in_1_bits_addr; // @[Bus.scala 47:23]
  wire  arbiter_io_in_2_valid; // @[Bus.scala 47:23]
  wire [38:0] arbiter_io_in_2_bits_addr; // @[Bus.scala 47:23]
  wire  arbiter_io_out_ready; // @[Bus.scala 47:23]
  wire  arbiter_io_out_valid; // @[Bus.scala 47:23]
  wire [38:0] arbiter_io_out_bits_addr; // @[Bus.scala 47:23]
  wire [63:0] arbiter_io_out_bits_wdata; // @[Bus.scala 47:23]
  wire [7:0] arbiter_io_out_bits_wmask; // @[Bus.scala 47:23]
  wire  arbiter_io_out_bits_wen; // @[Bus.scala 47:23]
  wire [1:0] arbiter_io_out_bits_len; // @[Bus.scala 47:23]
  wire  arbiter_io_out_bits_lrsc; // @[Bus.scala 47:23]
  wire [4:0] arbiter_io_out_bits_amo; // @[Bus.scala 47:23]
  wire [1:0] arbiter_io_chosen; // @[Bus.scala 47:23]
  wire  id_queue_clock; // @[Bus.scala 54:24]
  wire  id_queue_reset; // @[Bus.scala 54:24]
  wire  id_queue_io_enq_ready; // @[Bus.scala 54:24]
  wire  id_queue_io_enq_valid; // @[Bus.scala 54:24]
  wire [1:0] id_queue_io_enq_bits; // @[Bus.scala 54:24]
  wire  id_queue_io_deq_ready; // @[Bus.scala 54:24]
  wire  id_queue_io_deq_valid; // @[Bus.scala 54:24]
  wire [1:0] id_queue_io_deq_bits; // @[Bus.scala 54:24]
  wire  _GEN_0 = id_queue_io_deq_valid & id_queue_io_deq_bits == 2'h0 & io_in_0_resp_ready; // @[Bus.scala 75:25 78:67 79:27]
  wire  _GEN_2 = id_queue_io_deq_valid & id_queue_io_deq_bits == 2'h1 ? io_in_1_resp_ready : _GEN_0; // @[Bus.scala 78:67 79:27]
  RRArbiter arbiter ( // @[Bus.scala 47:23]
    .clock(arbiter_clock),
    .io_in_0_valid(arbiter_io_in_0_valid),
    .io_in_0_bits_addr(arbiter_io_in_0_bits_addr),
    .io_in_0_bits_wdata(arbiter_io_in_0_bits_wdata),
    .io_in_0_bits_wmask(arbiter_io_in_0_bits_wmask),
    .io_in_0_bits_wen(arbiter_io_in_0_bits_wen),
    .io_in_0_bits_len(arbiter_io_in_0_bits_len),
    .io_in_0_bits_lrsc(arbiter_io_in_0_bits_lrsc),
    .io_in_0_bits_amo(arbiter_io_in_0_bits_amo),
    .io_in_1_valid(arbiter_io_in_1_valid),
    .io_in_1_bits_addr(arbiter_io_in_1_bits_addr),
    .io_in_2_valid(arbiter_io_in_2_valid),
    .io_in_2_bits_addr(arbiter_io_in_2_bits_addr),
    .io_out_ready(arbiter_io_out_ready),
    .io_out_valid(arbiter_io_out_valid),
    .io_out_bits_addr(arbiter_io_out_bits_addr),
    .io_out_bits_wdata(arbiter_io_out_bits_wdata),
    .io_out_bits_wmask(arbiter_io_out_bits_wmask),
    .io_out_bits_wen(arbiter_io_out_bits_wen),
    .io_out_bits_len(arbiter_io_out_bits_len),
    .io_out_bits_lrsc(arbiter_io_out_bits_lrsc),
    .io_out_bits_amo(arbiter_io_out_bits_amo),
    .io_chosen(arbiter_io_chosen)
  );
  Queue_3 id_queue ( // @[Bus.scala 54:24]
    .clock(id_queue_clock),
    .reset(id_queue_reset),
    .io_enq_ready(id_queue_io_enq_ready),
    .io_enq_valid(id_queue_io_enq_valid),
    .io_enq_bits(id_queue_io_enq_bits),
    .io_deq_ready(id_queue_io_deq_ready),
    .io_deq_valid(id_queue_io_deq_valid),
    .io_deq_bits(id_queue_io_deq_bits)
  );
  assign io_in_0_req_ready = arbiter_io_chosen == 2'h0 & io_out_req_ready & id_queue_io_enq_ready; // @[Bus.scala 61:75]
  assign io_in_0_resp_valid = id_queue_io_deq_valid & id_queue_io_deq_bits == 2'h0 & io_out_resp_valid; // @[Bus.scala 74:25 78:67 80:27]
  assign io_in_0_resp_bits_rdata = io_out_resp_bits_rdata; // @[Bus.scala 73:25]
  assign io_in_1_req_ready = arbiter_io_chosen == 2'h1 & io_out_req_ready & id_queue_io_enq_ready; // @[Bus.scala 61:75]
  assign io_in_1_resp_valid = id_queue_io_deq_valid & id_queue_io_deq_bits == 2'h1 & io_out_resp_valid; // @[Bus.scala 74:25 78:67 80:27]
  assign io_in_1_resp_bits_rdata = io_out_resp_bits_rdata; // @[Bus.scala 73:25]
  assign io_in_2_req_ready = arbiter_io_chosen == 2'h2 & io_out_req_ready & id_queue_io_enq_ready; // @[Bus.scala 61:75]
  assign io_in_2_resp_valid = id_queue_io_deq_valid & id_queue_io_deq_bits == 2'h2 & io_out_resp_valid; // @[Bus.scala 74:25 78:67 80:27]
  assign io_in_2_resp_bits_rdata = io_out_resp_bits_rdata; // @[Bus.scala 73:25]
  assign io_out_req_valid = arbiter_io_out_valid; // @[Bus.scala 66:15]
  assign io_out_req_bits_addr = arbiter_io_out_bits_addr; // @[Bus.scala 65:15]
  assign io_out_req_bits_wdata = arbiter_io_out_bits_wdata; // @[Bus.scala 65:15]
  assign io_out_req_bits_wmask = arbiter_io_out_bits_wmask; // @[Bus.scala 65:15]
  assign io_out_req_bits_wen = arbiter_io_out_bits_wen; // @[Bus.scala 65:15]
  assign io_out_req_bits_len = arbiter_io_out_bits_len; // @[Bus.scala 65:15]
  assign io_out_req_bits_lrsc = arbiter_io_out_bits_lrsc; // @[Bus.scala 65:15]
  assign io_out_req_bits_amo = arbiter_io_out_bits_amo; // @[Bus.scala 65:15]
  assign io_out_resp_ready = id_queue_io_deq_valid & id_queue_io_deq_bits == 2'h2 ? io_in_2_resp_ready : _GEN_2; // @[Bus.scala 78:67 79:27]
  assign arbiter_clock = clock;
  assign arbiter_io_in_0_valid = io_in_0_req_valid; // @[Bus.scala 50:22]
  assign arbiter_io_in_0_bits_addr = io_in_0_req_bits_addr; // @[Bus.scala 50:22]
  assign arbiter_io_in_0_bits_wdata = io_in_0_req_bits_wdata; // @[Bus.scala 50:22]
  assign arbiter_io_in_0_bits_wmask = io_in_0_req_bits_wmask; // @[Bus.scala 50:22]
  assign arbiter_io_in_0_bits_wen = io_in_0_req_bits_wen; // @[Bus.scala 50:22]
  assign arbiter_io_in_0_bits_len = io_in_0_req_bits_len; // @[Bus.scala 50:22]
  assign arbiter_io_in_0_bits_lrsc = io_in_0_req_bits_lrsc; // @[Bus.scala 50:22]
  assign arbiter_io_in_0_bits_amo = io_in_0_req_bits_amo; // @[Bus.scala 50:22]
  assign arbiter_io_in_1_valid = io_in_1_req_valid; // @[Bus.scala 50:22]
  assign arbiter_io_in_1_bits_addr = io_in_1_req_bits_addr; // @[Bus.scala 50:22]
  assign arbiter_io_in_2_valid = io_in_2_req_valid; // @[Bus.scala 50:22]
  assign arbiter_io_in_2_bits_addr = io_in_2_req_bits_addr; // @[Bus.scala 50:22]
  assign arbiter_io_out_ready = io_out_req_ready; // @[Bus.scala 67:15]
  assign id_queue_clock = clock;
  assign id_queue_reset = reset;
  assign id_queue_io_enq_valid = io_out_req_ready & io_out_req_valid; // @[Decoupled.scala 51:35]
  assign id_queue_io_enq_bits = arbiter_io_chosen; // @[Bus.scala 56:25]
  assign id_queue_io_deq_ready = io_out_resp_ready & io_out_resp_valid; // @[Decoupled.scala 51:35]
endmodule
module SoCImp(
  input          clock,
  input          reset,
  input          auto_out_a_ready,
  output         auto_out_a_valid,
  output [2:0]   auto_out_a_bits_opcode,
  output [2:0]   auto_out_a_bits_param,
  output [2:0]   auto_out_a_bits_size,
  output [3:0]   auto_out_a_bits_source,
  output [31:0]  auto_out_a_bits_address,
  output [31:0]  auto_out_a_bits_mask,
  output [255:0] auto_out_a_bits_data,
  output         auto_out_b_ready,
  input          auto_out_b_valid,
  input  [2:0]   auto_out_b_bits_size,
  input  [3:0]   auto_out_b_bits_source,
  input  [31:0]  auto_out_b_bits_address,
  input          auto_out_c_ready,
  output         auto_out_c_valid,
  output [2:0]   auto_out_c_bits_opcode,
  output [2:0]   auto_out_c_bits_param,
  output [2:0]   auto_out_c_bits_size,
  output [3:0]   auto_out_c_bits_source,
  output [31:0]  auto_out_c_bits_address,
  output [255:0] auto_out_c_bits_data,
  output         auto_out_d_ready,
  input          auto_out_d_valid,
  input  [2:0]   auto_out_d_bits_opcode,
  input  [2:0]   auto_out_d_bits_size,
  input  [3:0]   auto_out_d_bits_source,
  input  [5:0]   auto_out_d_bits_sink,
  input  [255:0] auto_out_d_bits_data,
  input          auto_out_e_ready,
  output         auto_out_e_valid,
  output [5:0]   auto_out_e_bits_sink,
  input          io_intr_mtip,
  input          io_intr_msip,
  input          io_intr_meip,
  input          io_intr_seip
);
  wire  icache_clock; // @[SoC.scala 27:27]
  wire  icache_reset; // @[SoC.scala 27:27]
  wire  icache_auto_out_a_ready; // @[SoC.scala 27:27]
  wire  icache_auto_out_a_valid; // @[SoC.scala 27:27]
  wire [1:0] icache_auto_out_a_bits_source; // @[SoC.scala 27:27]
  wire [31:0] icache_auto_out_a_bits_address; // @[SoC.scala 27:27]
  wire  icache_auto_out_d_ready; // @[SoC.scala 27:27]
  wire  icache_auto_out_d_valid; // @[SoC.scala 27:27]
  wire [255:0] icache_auto_out_d_bits_data; // @[SoC.scala 27:27]
  wire  icache_io_cache_req_ready; // @[SoC.scala 27:27]
  wire  icache_io_cache_req_valid; // @[SoC.scala 27:27]
  wire [38:0] icache_io_cache_req_bits_addr; // @[SoC.scala 27:27]
  wire  icache_io_cache_resp_ready; // @[SoC.scala 27:27]
  wire  icache_io_cache_resp_valid; // @[SoC.scala 27:27]
  wire [63:0] icache_io_cache_resp_bits_rdata; // @[SoC.scala 27:27]
  wire  icache_io_fence_i; // @[SoC.scala 27:27]
  wire  dcache_clock; // @[SoC.scala 28:27]
  wire  dcache_reset; // @[SoC.scala 28:27]
  wire  dcache_auto_out_a_ready; // @[SoC.scala 28:27]
  wire  dcache_auto_out_a_valid; // @[SoC.scala 28:27]
  wire [1:0] dcache_auto_out_a_bits_source; // @[SoC.scala 28:27]
  wire [31:0] dcache_auto_out_a_bits_address; // @[SoC.scala 28:27]
  wire  dcache_auto_out_b_ready; // @[SoC.scala 28:27]
  wire  dcache_auto_out_b_valid; // @[SoC.scala 28:27]
  wire [2:0] dcache_auto_out_b_bits_size; // @[SoC.scala 28:27]
  wire [1:0] dcache_auto_out_b_bits_source; // @[SoC.scala 28:27]
  wire [31:0] dcache_auto_out_b_bits_address; // @[SoC.scala 28:27]
  wire  dcache_auto_out_c_ready; // @[SoC.scala 28:27]
  wire  dcache_auto_out_c_valid; // @[SoC.scala 28:27]
  wire [2:0] dcache_auto_out_c_bits_opcode; // @[SoC.scala 28:27]
  wire [2:0] dcache_auto_out_c_bits_param; // @[SoC.scala 28:27]
  wire [2:0] dcache_auto_out_c_bits_size; // @[SoC.scala 28:27]
  wire [1:0] dcache_auto_out_c_bits_source; // @[SoC.scala 28:27]
  wire [31:0] dcache_auto_out_c_bits_address; // @[SoC.scala 28:27]
  wire [255:0] dcache_auto_out_c_bits_data; // @[SoC.scala 28:27]
  wire  dcache_auto_out_d_ready; // @[SoC.scala 28:27]
  wire  dcache_auto_out_d_valid; // @[SoC.scala 28:27]
  wire [5:0] dcache_auto_out_d_bits_sink; // @[SoC.scala 28:27]
  wire [255:0] dcache_auto_out_d_bits_data; // @[SoC.scala 28:27]
  wire  dcache_auto_out_e_ready; // @[SoC.scala 28:27]
  wire  dcache_auto_out_e_valid; // @[SoC.scala 28:27]
  wire [5:0] dcache_auto_out_e_bits_sink; // @[SoC.scala 28:27]
  wire  dcache_io_cache_req_ready; // @[SoC.scala 28:27]
  wire  dcache_io_cache_req_valid; // @[SoC.scala 28:27]
  wire [38:0] dcache_io_cache_req_bits_addr; // @[SoC.scala 28:27]
  wire [63:0] dcache_io_cache_req_bits_wdata; // @[SoC.scala 28:27]
  wire [7:0] dcache_io_cache_req_bits_wmask; // @[SoC.scala 28:27]
  wire  dcache_io_cache_req_bits_wen; // @[SoC.scala 28:27]
  wire [1:0] dcache_io_cache_req_bits_len; // @[SoC.scala 28:27]
  wire  dcache_io_cache_req_bits_lrsc; // @[SoC.scala 28:27]
  wire [4:0] dcache_io_cache_req_bits_amo; // @[SoC.scala 28:27]
  wire  dcache_io_cache_resp_ready; // @[SoC.scala 28:27]
  wire  dcache_io_cache_resp_valid; // @[SoC.scala 28:27]
  wire [63:0] dcache_io_cache_resp_bits_rdata; // @[SoC.scala 28:27]
  wire  uncache_clock; // @[SoC.scala 29:27]
  wire  uncache_reset; // @[SoC.scala 29:27]
  wire  uncache_auto_out_a_ready; // @[SoC.scala 29:27]
  wire  uncache_auto_out_a_valid; // @[SoC.scala 29:27]
  wire [2:0] uncache_auto_out_a_bits_opcode; // @[SoC.scala 29:27]
  wire [2:0] uncache_auto_out_a_bits_size; // @[SoC.scala 29:27]
  wire [1:0] uncache_auto_out_a_bits_source; // @[SoC.scala 29:27]
  wire [31:0] uncache_auto_out_a_bits_address; // @[SoC.scala 29:27]
  wire [7:0] uncache_auto_out_a_bits_mask; // @[SoC.scala 29:27]
  wire [63:0] uncache_auto_out_a_bits_data; // @[SoC.scala 29:27]
  wire  uncache_auto_out_d_ready; // @[SoC.scala 29:27]
  wire  uncache_auto_out_d_valid; // @[SoC.scala 29:27]
  wire [63:0] uncache_auto_out_d_bits_data; // @[SoC.scala 29:27]
  wire  uncache_io_in_req_ready; // @[SoC.scala 29:27]
  wire  uncache_io_in_req_valid; // @[SoC.scala 29:27]
  wire [38:0] uncache_io_in_req_bits_addr; // @[SoC.scala 29:27]
  wire [63:0] uncache_io_in_req_bits_wdata; // @[SoC.scala 29:27]
  wire [7:0] uncache_io_in_req_bits_wmask; // @[SoC.scala 29:27]
  wire  uncache_io_in_req_bits_wen; // @[SoC.scala 29:27]
  wire [1:0] uncache_io_in_req_bits_len; // @[SoC.scala 29:27]
  wire  uncache_io_in_resp_ready; // @[SoC.scala 29:27]
  wire  uncache_io_in_resp_valid; // @[SoC.scala 29:27]
  wire [63:0] uncache_io_in_resp_bits_rdata; // @[SoC.scala 29:27]
  wire  xbar_clock; // @[SoC.scala 30:27]
  wire  xbar_reset; // @[SoC.scala 30:27]
  wire  xbar_auto_in_2_a_ready; // @[SoC.scala 30:27]
  wire  xbar_auto_in_2_a_valid; // @[SoC.scala 30:27]
  wire [1:0] xbar_auto_in_2_a_bits_source; // @[SoC.scala 30:27]
  wire [31:0] xbar_auto_in_2_a_bits_address; // @[SoC.scala 30:27]
  wire  xbar_auto_in_2_b_ready; // @[SoC.scala 30:27]
  wire  xbar_auto_in_2_b_valid; // @[SoC.scala 30:27]
  wire [2:0] xbar_auto_in_2_b_bits_size; // @[SoC.scala 30:27]
  wire [1:0] xbar_auto_in_2_b_bits_source; // @[SoC.scala 30:27]
  wire [31:0] xbar_auto_in_2_b_bits_address; // @[SoC.scala 30:27]
  wire  xbar_auto_in_2_c_ready; // @[SoC.scala 30:27]
  wire  xbar_auto_in_2_c_valid; // @[SoC.scala 30:27]
  wire [2:0] xbar_auto_in_2_c_bits_opcode; // @[SoC.scala 30:27]
  wire [2:0] xbar_auto_in_2_c_bits_param; // @[SoC.scala 30:27]
  wire [2:0] xbar_auto_in_2_c_bits_size; // @[SoC.scala 30:27]
  wire [1:0] xbar_auto_in_2_c_bits_source; // @[SoC.scala 30:27]
  wire [31:0] xbar_auto_in_2_c_bits_address; // @[SoC.scala 30:27]
  wire [255:0] xbar_auto_in_2_c_bits_data; // @[SoC.scala 30:27]
  wire  xbar_auto_in_2_d_ready; // @[SoC.scala 30:27]
  wire  xbar_auto_in_2_d_valid; // @[SoC.scala 30:27]
  wire [5:0] xbar_auto_in_2_d_bits_sink; // @[SoC.scala 30:27]
  wire [255:0] xbar_auto_in_2_d_bits_data; // @[SoC.scala 30:27]
  wire  xbar_auto_in_2_e_ready; // @[SoC.scala 30:27]
  wire  xbar_auto_in_2_e_valid; // @[SoC.scala 30:27]
  wire [5:0] xbar_auto_in_2_e_bits_sink; // @[SoC.scala 30:27]
  wire  xbar_auto_in_1_a_ready; // @[SoC.scala 30:27]
  wire  xbar_auto_in_1_a_valid; // @[SoC.scala 30:27]
  wire [2:0] xbar_auto_in_1_a_bits_opcode; // @[SoC.scala 30:27]
  wire [2:0] xbar_auto_in_1_a_bits_size; // @[SoC.scala 30:27]
  wire [1:0] xbar_auto_in_1_a_bits_source; // @[SoC.scala 30:27]
  wire [31:0] xbar_auto_in_1_a_bits_address; // @[SoC.scala 30:27]
  wire [31:0] xbar_auto_in_1_a_bits_mask; // @[SoC.scala 30:27]
  wire [255:0] xbar_auto_in_1_a_bits_data; // @[SoC.scala 30:27]
  wire  xbar_auto_in_1_d_ready; // @[SoC.scala 30:27]
  wire  xbar_auto_in_1_d_valid; // @[SoC.scala 30:27]
  wire [2:0] xbar_auto_in_1_d_bits_opcode; // @[SoC.scala 30:27]
  wire [2:0] xbar_auto_in_1_d_bits_size; // @[SoC.scala 30:27]
  wire [1:0] xbar_auto_in_1_d_bits_source; // @[SoC.scala 30:27]
  wire [255:0] xbar_auto_in_1_d_bits_data; // @[SoC.scala 30:27]
  wire  xbar_auto_in_0_a_ready; // @[SoC.scala 30:27]
  wire  xbar_auto_in_0_a_valid; // @[SoC.scala 30:27]
  wire [1:0] xbar_auto_in_0_a_bits_source; // @[SoC.scala 30:27]
  wire [31:0] xbar_auto_in_0_a_bits_address; // @[SoC.scala 30:27]
  wire  xbar_auto_in_0_d_ready; // @[SoC.scala 30:27]
  wire  xbar_auto_in_0_d_valid; // @[SoC.scala 30:27]
  wire [255:0] xbar_auto_in_0_d_bits_data; // @[SoC.scala 30:27]
  wire  xbar_auto_out_a_ready; // @[SoC.scala 30:27]
  wire  xbar_auto_out_a_valid; // @[SoC.scala 30:27]
  wire [2:0] xbar_auto_out_a_bits_opcode; // @[SoC.scala 30:27]
  wire [2:0] xbar_auto_out_a_bits_param; // @[SoC.scala 30:27]
  wire [2:0] xbar_auto_out_a_bits_size; // @[SoC.scala 30:27]
  wire [3:0] xbar_auto_out_a_bits_source; // @[SoC.scala 30:27]
  wire [31:0] xbar_auto_out_a_bits_address; // @[SoC.scala 30:27]
  wire [31:0] xbar_auto_out_a_bits_mask; // @[SoC.scala 30:27]
  wire [255:0] xbar_auto_out_a_bits_data; // @[SoC.scala 30:27]
  wire  xbar_auto_out_b_ready; // @[SoC.scala 30:27]
  wire  xbar_auto_out_b_valid; // @[SoC.scala 30:27]
  wire [2:0] xbar_auto_out_b_bits_size; // @[SoC.scala 30:27]
  wire [3:0] xbar_auto_out_b_bits_source; // @[SoC.scala 30:27]
  wire [31:0] xbar_auto_out_b_bits_address; // @[SoC.scala 30:27]
  wire  xbar_auto_out_c_ready; // @[SoC.scala 30:27]
  wire  xbar_auto_out_c_valid; // @[SoC.scala 30:27]
  wire [2:0] xbar_auto_out_c_bits_opcode; // @[SoC.scala 30:27]
  wire [2:0] xbar_auto_out_c_bits_param; // @[SoC.scala 30:27]
  wire [2:0] xbar_auto_out_c_bits_size; // @[SoC.scala 30:27]
  wire [3:0] xbar_auto_out_c_bits_source; // @[SoC.scala 30:27]
  wire [31:0] xbar_auto_out_c_bits_address; // @[SoC.scala 30:27]
  wire [255:0] xbar_auto_out_c_bits_data; // @[SoC.scala 30:27]
  wire  xbar_auto_out_d_ready; // @[SoC.scala 30:27]
  wire  xbar_auto_out_d_valid; // @[SoC.scala 30:27]
  wire [2:0] xbar_auto_out_d_bits_opcode; // @[SoC.scala 30:27]
  wire [2:0] xbar_auto_out_d_bits_size; // @[SoC.scala 30:27]
  wire [3:0] xbar_auto_out_d_bits_source; // @[SoC.scala 30:27]
  wire [5:0] xbar_auto_out_d_bits_sink; // @[SoC.scala 30:27]
  wire [255:0] xbar_auto_out_d_bits_data; // @[SoC.scala 30:27]
  wire  xbar_auto_out_e_ready; // @[SoC.scala 30:27]
  wire  xbar_auto_out_e_valid; // @[SoC.scala 30:27]
  wire [5:0] xbar_auto_out_e_bits_sink; // @[SoC.scala 30:27]
  wire  widget_clock; // @[WidthWidget.scala 220:28]
  wire  widget_reset; // @[WidthWidget.scala 220:28]
  wire  widget_auto_in_a_ready; // @[WidthWidget.scala 220:28]
  wire  widget_auto_in_a_valid; // @[WidthWidget.scala 220:28]
  wire [2:0] widget_auto_in_a_bits_opcode; // @[WidthWidget.scala 220:28]
  wire [2:0] widget_auto_in_a_bits_size; // @[WidthWidget.scala 220:28]
  wire [1:0] widget_auto_in_a_bits_source; // @[WidthWidget.scala 220:28]
  wire [31:0] widget_auto_in_a_bits_address; // @[WidthWidget.scala 220:28]
  wire [7:0] widget_auto_in_a_bits_mask; // @[WidthWidget.scala 220:28]
  wire [63:0] widget_auto_in_a_bits_data; // @[WidthWidget.scala 220:28]
  wire  widget_auto_in_d_ready; // @[WidthWidget.scala 220:28]
  wire  widget_auto_in_d_valid; // @[WidthWidget.scala 220:28]
  wire [63:0] widget_auto_in_d_bits_data; // @[WidthWidget.scala 220:28]
  wire  widget_auto_out_a_ready; // @[WidthWidget.scala 220:28]
  wire  widget_auto_out_a_valid; // @[WidthWidget.scala 220:28]
  wire [2:0] widget_auto_out_a_bits_opcode; // @[WidthWidget.scala 220:28]
  wire [2:0] widget_auto_out_a_bits_size; // @[WidthWidget.scala 220:28]
  wire [1:0] widget_auto_out_a_bits_source; // @[WidthWidget.scala 220:28]
  wire [31:0] widget_auto_out_a_bits_address; // @[WidthWidget.scala 220:28]
  wire [31:0] widget_auto_out_a_bits_mask; // @[WidthWidget.scala 220:28]
  wire [255:0] widget_auto_out_a_bits_data; // @[WidthWidget.scala 220:28]
  wire  widget_auto_out_d_ready; // @[WidthWidget.scala 220:28]
  wire  widget_auto_out_d_valid; // @[WidthWidget.scala 220:28]
  wire [2:0] widget_auto_out_d_bits_opcode; // @[WidthWidget.scala 220:28]
  wire [2:0] widget_auto_out_d_bits_size; // @[WidthWidget.scala 220:28]
  wire [1:0] widget_auto_out_d_bits_source; // @[WidthWidget.scala 220:28]
  wire [255:0] widget_auto_out_d_bits_data; // @[WidthWidget.scala 220:28]
  wire  core_clock; // @[SoC.scala 40:22]
  wire  core_reset; // @[SoC.scala 40:22]
  wire  core_io_imem_req_ready; // @[SoC.scala 40:22]
  wire  core_io_imem_req_valid; // @[SoC.scala 40:22]
  wire [38:0] core_io_imem_req_bits_addr; // @[SoC.scala 40:22]
  wire  core_io_imem_resp_ready; // @[SoC.scala 40:22]
  wire  core_io_imem_resp_valid; // @[SoC.scala 40:22]
  wire [63:0] core_io_imem_resp_bits_rdata; // @[SoC.scala 40:22]
  wire  core_io_dmem_req_ready; // @[SoC.scala 40:22]
  wire  core_io_dmem_req_valid; // @[SoC.scala 40:22]
  wire [38:0] core_io_dmem_req_bits_addr; // @[SoC.scala 40:22]
  wire [63:0] core_io_dmem_req_bits_wdata; // @[SoC.scala 40:22]
  wire [7:0] core_io_dmem_req_bits_wmask; // @[SoC.scala 40:22]
  wire  core_io_dmem_req_bits_wen; // @[SoC.scala 40:22]
  wire [1:0] core_io_dmem_req_bits_len; // @[SoC.scala 40:22]
  wire  core_io_dmem_req_bits_lrsc; // @[SoC.scala 40:22]
  wire [4:0] core_io_dmem_req_bits_amo; // @[SoC.scala 40:22]
  wire  core_io_dmem_resp_ready; // @[SoC.scala 40:22]
  wire  core_io_dmem_resp_valid; // @[SoC.scala 40:22]
  wire [63:0] core_io_dmem_resp_bits_rdata; // @[SoC.scala 40:22]
  wire  core_io_iptw_req_ready; // @[SoC.scala 40:22]
  wire  core_io_iptw_req_valid; // @[SoC.scala 40:22]
  wire [38:0] core_io_iptw_req_bits_addr; // @[SoC.scala 40:22]
  wire  core_io_iptw_resp_ready; // @[SoC.scala 40:22]
  wire  core_io_iptw_resp_valid; // @[SoC.scala 40:22]
  wire [63:0] core_io_iptw_resp_bits_rdata; // @[SoC.scala 40:22]
  wire  core_io_dptw_req_ready; // @[SoC.scala 40:22]
  wire  core_io_dptw_req_valid; // @[SoC.scala 40:22]
  wire [38:0] core_io_dptw_req_bits_addr; // @[SoC.scala 40:22]
  wire  core_io_dptw_resp_ready; // @[SoC.scala 40:22]
  wire  core_io_dptw_resp_valid; // @[SoC.scala 40:22]
  wire [63:0] core_io_dptw_resp_bits_rdata; // @[SoC.scala 40:22]
  wire  core_io_uncache_req_ready; // @[SoC.scala 40:22]
  wire  core_io_uncache_req_valid; // @[SoC.scala 40:22]
  wire [38:0] core_io_uncache_req_bits_addr; // @[SoC.scala 40:22]
  wire [63:0] core_io_uncache_req_bits_wdata; // @[SoC.scala 40:22]
  wire [7:0] core_io_uncache_req_bits_wmask; // @[SoC.scala 40:22]
  wire  core_io_uncache_req_bits_wen; // @[SoC.scala 40:22]
  wire [1:0] core_io_uncache_req_bits_len; // @[SoC.scala 40:22]
  wire  core_io_uncache_resp_ready; // @[SoC.scala 40:22]
  wire  core_io_uncache_resp_valid; // @[SoC.scala 40:22]
  wire [63:0] core_io_uncache_resp_bits_rdata; // @[SoC.scala 40:22]
  wire  core_io_fence_i; // @[SoC.scala 40:22]
  wire  core_io_intr_mtip; // @[SoC.scala 40:22]
  wire  core_io_intr_msip; // @[SoC.scala 40:22]
  wire  core_io_intr_meip; // @[SoC.scala 40:22]
  wire  core_io_intr_seip; // @[SoC.scala 40:22]
  wire  xbar_1_clock; // @[SoC.scala 50:22]
  wire  xbar_1_reset; // @[SoC.scala 50:22]
  wire  xbar_1_io_in_0_req_ready; // @[SoC.scala 50:22]
  wire  xbar_1_io_in_0_req_valid; // @[SoC.scala 50:22]
  wire [38:0] xbar_1_io_in_0_req_bits_addr; // @[SoC.scala 50:22]
  wire [63:0] xbar_1_io_in_0_req_bits_wdata; // @[SoC.scala 50:22]
  wire [7:0] xbar_1_io_in_0_req_bits_wmask; // @[SoC.scala 50:22]
  wire  xbar_1_io_in_0_req_bits_wen; // @[SoC.scala 50:22]
  wire [1:0] xbar_1_io_in_0_req_bits_len; // @[SoC.scala 50:22]
  wire  xbar_1_io_in_0_req_bits_lrsc; // @[SoC.scala 50:22]
  wire [4:0] xbar_1_io_in_0_req_bits_amo; // @[SoC.scala 50:22]
  wire  xbar_1_io_in_0_resp_ready; // @[SoC.scala 50:22]
  wire  xbar_1_io_in_0_resp_valid; // @[SoC.scala 50:22]
  wire [63:0] xbar_1_io_in_0_resp_bits_rdata; // @[SoC.scala 50:22]
  wire  xbar_1_io_in_1_req_ready; // @[SoC.scala 50:22]
  wire  xbar_1_io_in_1_req_valid; // @[SoC.scala 50:22]
  wire [38:0] xbar_1_io_in_1_req_bits_addr; // @[SoC.scala 50:22]
  wire  xbar_1_io_in_1_resp_ready; // @[SoC.scala 50:22]
  wire  xbar_1_io_in_1_resp_valid; // @[SoC.scala 50:22]
  wire [63:0] xbar_1_io_in_1_resp_bits_rdata; // @[SoC.scala 50:22]
  wire  xbar_1_io_in_2_req_ready; // @[SoC.scala 50:22]
  wire  xbar_1_io_in_2_req_valid; // @[SoC.scala 50:22]
  wire [38:0] xbar_1_io_in_2_req_bits_addr; // @[SoC.scala 50:22]
  wire  xbar_1_io_in_2_resp_ready; // @[SoC.scala 50:22]
  wire  xbar_1_io_in_2_resp_valid; // @[SoC.scala 50:22]
  wire [63:0] xbar_1_io_in_2_resp_bits_rdata; // @[SoC.scala 50:22]
  wire  xbar_1_io_out_req_ready; // @[SoC.scala 50:22]
  wire  xbar_1_io_out_req_valid; // @[SoC.scala 50:22]
  wire [38:0] xbar_1_io_out_req_bits_addr; // @[SoC.scala 50:22]
  wire [63:0] xbar_1_io_out_req_bits_wdata; // @[SoC.scala 50:22]
  wire [7:0] xbar_1_io_out_req_bits_wmask; // @[SoC.scala 50:22]
  wire  xbar_1_io_out_req_bits_wen; // @[SoC.scala 50:22]
  wire [1:0] xbar_1_io_out_req_bits_len; // @[SoC.scala 50:22]
  wire  xbar_1_io_out_req_bits_lrsc; // @[SoC.scala 50:22]
  wire [4:0] xbar_1_io_out_req_bits_amo; // @[SoC.scala 50:22]
  wire  xbar_1_io_out_resp_ready; // @[SoC.scala 50:22]
  wire  xbar_1_io_out_resp_valid; // @[SoC.scala 50:22]
  wire [63:0] xbar_1_io_out_resp_bits_rdata; // @[SoC.scala 50:22]
  ICache icache ( // @[SoC.scala 27:27]
    .clock(icache_clock),
    .reset(icache_reset),
    .auto_out_a_ready(icache_auto_out_a_ready),
    .auto_out_a_valid(icache_auto_out_a_valid),
    .auto_out_a_bits_source(icache_auto_out_a_bits_source),
    .auto_out_a_bits_address(icache_auto_out_a_bits_address),
    .auto_out_d_ready(icache_auto_out_d_ready),
    .auto_out_d_valid(icache_auto_out_d_valid),
    .auto_out_d_bits_data(icache_auto_out_d_bits_data),
    .io_cache_req_ready(icache_io_cache_req_ready),
    .io_cache_req_valid(icache_io_cache_req_valid),
    .io_cache_req_bits_addr(icache_io_cache_req_bits_addr),
    .io_cache_resp_ready(icache_io_cache_resp_ready),
    .io_cache_resp_valid(icache_io_cache_resp_valid),
    .io_cache_resp_bits_rdata(icache_io_cache_resp_bits_rdata),
    .io_fence_i(icache_io_fence_i)
  );
  DCache dcache ( // @[SoC.scala 28:27]
    .clock(dcache_clock),
    .reset(dcache_reset),
    .auto_out_a_ready(dcache_auto_out_a_ready),
    .auto_out_a_valid(dcache_auto_out_a_valid),
    .auto_out_a_bits_source(dcache_auto_out_a_bits_source),
    .auto_out_a_bits_address(dcache_auto_out_a_bits_address),
    .auto_out_b_ready(dcache_auto_out_b_ready),
    .auto_out_b_valid(dcache_auto_out_b_valid),
    .auto_out_b_bits_size(dcache_auto_out_b_bits_size),
    .auto_out_b_bits_source(dcache_auto_out_b_bits_source),
    .auto_out_b_bits_address(dcache_auto_out_b_bits_address),
    .auto_out_c_ready(dcache_auto_out_c_ready),
    .auto_out_c_valid(dcache_auto_out_c_valid),
    .auto_out_c_bits_opcode(dcache_auto_out_c_bits_opcode),
    .auto_out_c_bits_param(dcache_auto_out_c_bits_param),
    .auto_out_c_bits_size(dcache_auto_out_c_bits_size),
    .auto_out_c_bits_source(dcache_auto_out_c_bits_source),
    .auto_out_c_bits_address(dcache_auto_out_c_bits_address),
    .auto_out_c_bits_data(dcache_auto_out_c_bits_data),
    .auto_out_d_ready(dcache_auto_out_d_ready),
    .auto_out_d_valid(dcache_auto_out_d_valid),
    .auto_out_d_bits_sink(dcache_auto_out_d_bits_sink),
    .auto_out_d_bits_data(dcache_auto_out_d_bits_data),
    .auto_out_e_ready(dcache_auto_out_e_ready),
    .auto_out_e_valid(dcache_auto_out_e_valid),
    .auto_out_e_bits_sink(dcache_auto_out_e_bits_sink),
    .io_cache_req_ready(dcache_io_cache_req_ready),
    .io_cache_req_valid(dcache_io_cache_req_valid),
    .io_cache_req_bits_addr(dcache_io_cache_req_bits_addr),
    .io_cache_req_bits_wdata(dcache_io_cache_req_bits_wdata),
    .io_cache_req_bits_wmask(dcache_io_cache_req_bits_wmask),
    .io_cache_req_bits_wen(dcache_io_cache_req_bits_wen),
    .io_cache_req_bits_len(dcache_io_cache_req_bits_len),
    .io_cache_req_bits_lrsc(dcache_io_cache_req_bits_lrsc),
    .io_cache_req_bits_amo(dcache_io_cache_req_bits_amo),
    .io_cache_resp_ready(dcache_io_cache_resp_ready),
    .io_cache_resp_valid(dcache_io_cache_resp_valid),
    .io_cache_resp_bits_rdata(dcache_io_cache_resp_bits_rdata)
  );
  Uncache uncache ( // @[SoC.scala 29:27]
    .clock(uncache_clock),
    .reset(uncache_reset),
    .auto_out_a_ready(uncache_auto_out_a_ready),
    .auto_out_a_valid(uncache_auto_out_a_valid),
    .auto_out_a_bits_opcode(uncache_auto_out_a_bits_opcode),
    .auto_out_a_bits_size(uncache_auto_out_a_bits_size),
    .auto_out_a_bits_source(uncache_auto_out_a_bits_source),
    .auto_out_a_bits_address(uncache_auto_out_a_bits_address),
    .auto_out_a_bits_mask(uncache_auto_out_a_bits_mask),
    .auto_out_a_bits_data(uncache_auto_out_a_bits_data),
    .auto_out_d_ready(uncache_auto_out_d_ready),
    .auto_out_d_valid(uncache_auto_out_d_valid),
    .auto_out_d_bits_data(uncache_auto_out_d_bits_data),
    .io_in_req_ready(uncache_io_in_req_ready),
    .io_in_req_valid(uncache_io_in_req_valid),
    .io_in_req_bits_addr(uncache_io_in_req_bits_addr),
    .io_in_req_bits_wdata(uncache_io_in_req_bits_wdata),
    .io_in_req_bits_wmask(uncache_io_in_req_bits_wmask),
    .io_in_req_bits_wen(uncache_io_in_req_bits_wen),
    .io_in_req_bits_len(uncache_io_in_req_bits_len),
    .io_in_resp_ready(uncache_io_in_resp_ready),
    .io_in_resp_valid(uncache_io_in_resp_valid),
    .io_in_resp_bits_rdata(uncache_io_in_resp_bits_rdata)
  );
  TLXbar xbar ( // @[SoC.scala 30:27]
    .clock(xbar_clock),
    .reset(xbar_reset),
    .auto_in_2_a_ready(xbar_auto_in_2_a_ready),
    .auto_in_2_a_valid(xbar_auto_in_2_a_valid),
    .auto_in_2_a_bits_source(xbar_auto_in_2_a_bits_source),
    .auto_in_2_a_bits_address(xbar_auto_in_2_a_bits_address),
    .auto_in_2_b_ready(xbar_auto_in_2_b_ready),
    .auto_in_2_b_valid(xbar_auto_in_2_b_valid),
    .auto_in_2_b_bits_size(xbar_auto_in_2_b_bits_size),
    .auto_in_2_b_bits_source(xbar_auto_in_2_b_bits_source),
    .auto_in_2_b_bits_address(xbar_auto_in_2_b_bits_address),
    .auto_in_2_c_ready(xbar_auto_in_2_c_ready),
    .auto_in_2_c_valid(xbar_auto_in_2_c_valid),
    .auto_in_2_c_bits_opcode(xbar_auto_in_2_c_bits_opcode),
    .auto_in_2_c_bits_param(xbar_auto_in_2_c_bits_param),
    .auto_in_2_c_bits_size(xbar_auto_in_2_c_bits_size),
    .auto_in_2_c_bits_source(xbar_auto_in_2_c_bits_source),
    .auto_in_2_c_bits_address(xbar_auto_in_2_c_bits_address),
    .auto_in_2_c_bits_data(xbar_auto_in_2_c_bits_data),
    .auto_in_2_d_ready(xbar_auto_in_2_d_ready),
    .auto_in_2_d_valid(xbar_auto_in_2_d_valid),
    .auto_in_2_d_bits_sink(xbar_auto_in_2_d_bits_sink),
    .auto_in_2_d_bits_data(xbar_auto_in_2_d_bits_data),
    .auto_in_2_e_ready(xbar_auto_in_2_e_ready),
    .auto_in_2_e_valid(xbar_auto_in_2_e_valid),
    .auto_in_2_e_bits_sink(xbar_auto_in_2_e_bits_sink),
    .auto_in_1_a_ready(xbar_auto_in_1_a_ready),
    .auto_in_1_a_valid(xbar_auto_in_1_a_valid),
    .auto_in_1_a_bits_opcode(xbar_auto_in_1_a_bits_opcode),
    .auto_in_1_a_bits_size(xbar_auto_in_1_a_bits_size),
    .auto_in_1_a_bits_source(xbar_auto_in_1_a_bits_source),
    .auto_in_1_a_bits_address(xbar_auto_in_1_a_bits_address),
    .auto_in_1_a_bits_mask(xbar_auto_in_1_a_bits_mask),
    .auto_in_1_a_bits_data(xbar_auto_in_1_a_bits_data),
    .auto_in_1_d_ready(xbar_auto_in_1_d_ready),
    .auto_in_1_d_valid(xbar_auto_in_1_d_valid),
    .auto_in_1_d_bits_opcode(xbar_auto_in_1_d_bits_opcode),
    .auto_in_1_d_bits_size(xbar_auto_in_1_d_bits_size),
    .auto_in_1_d_bits_source(xbar_auto_in_1_d_bits_source),
    .auto_in_1_d_bits_data(xbar_auto_in_1_d_bits_data),
    .auto_in_0_a_ready(xbar_auto_in_0_a_ready),
    .auto_in_0_a_valid(xbar_auto_in_0_a_valid),
    .auto_in_0_a_bits_source(xbar_auto_in_0_a_bits_source),
    .auto_in_0_a_bits_address(xbar_auto_in_0_a_bits_address),
    .auto_in_0_d_ready(xbar_auto_in_0_d_ready),
    .auto_in_0_d_valid(xbar_auto_in_0_d_valid),
    .auto_in_0_d_bits_data(xbar_auto_in_0_d_bits_data),
    .auto_out_a_ready(xbar_auto_out_a_ready),
    .auto_out_a_valid(xbar_auto_out_a_valid),
    .auto_out_a_bits_opcode(xbar_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(xbar_auto_out_a_bits_param),
    .auto_out_a_bits_size(xbar_auto_out_a_bits_size),
    .auto_out_a_bits_source(xbar_auto_out_a_bits_source),
    .auto_out_a_bits_address(xbar_auto_out_a_bits_address),
    .auto_out_a_bits_mask(xbar_auto_out_a_bits_mask),
    .auto_out_a_bits_data(xbar_auto_out_a_bits_data),
    .auto_out_b_ready(xbar_auto_out_b_ready),
    .auto_out_b_valid(xbar_auto_out_b_valid),
    .auto_out_b_bits_size(xbar_auto_out_b_bits_size),
    .auto_out_b_bits_source(xbar_auto_out_b_bits_source),
    .auto_out_b_bits_address(xbar_auto_out_b_bits_address),
    .auto_out_c_ready(xbar_auto_out_c_ready),
    .auto_out_c_valid(xbar_auto_out_c_valid),
    .auto_out_c_bits_opcode(xbar_auto_out_c_bits_opcode),
    .auto_out_c_bits_param(xbar_auto_out_c_bits_param),
    .auto_out_c_bits_size(xbar_auto_out_c_bits_size),
    .auto_out_c_bits_source(xbar_auto_out_c_bits_source),
    .auto_out_c_bits_address(xbar_auto_out_c_bits_address),
    .auto_out_c_bits_data(xbar_auto_out_c_bits_data),
    .auto_out_d_ready(xbar_auto_out_d_ready),
    .auto_out_d_valid(xbar_auto_out_d_valid),
    .auto_out_d_bits_opcode(xbar_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(xbar_auto_out_d_bits_size),
    .auto_out_d_bits_source(xbar_auto_out_d_bits_source),
    .auto_out_d_bits_sink(xbar_auto_out_d_bits_sink),
    .auto_out_d_bits_data(xbar_auto_out_d_bits_data),
    .auto_out_e_ready(xbar_auto_out_e_ready),
    .auto_out_e_valid(xbar_auto_out_e_valid),
    .auto_out_e_bits_sink(xbar_auto_out_e_bits_sink)
  );
  TLWidthWidget widget ( // @[WidthWidget.scala 220:28]
    .clock(widget_clock),
    .reset(widget_reset),
    .auto_in_a_ready(widget_auto_in_a_ready),
    .auto_in_a_valid(widget_auto_in_a_valid),
    .auto_in_a_bits_opcode(widget_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(widget_auto_in_a_bits_size),
    .auto_in_a_bits_source(widget_auto_in_a_bits_source),
    .auto_in_a_bits_address(widget_auto_in_a_bits_address),
    .auto_in_a_bits_mask(widget_auto_in_a_bits_mask),
    .auto_in_a_bits_data(widget_auto_in_a_bits_data),
    .auto_in_d_ready(widget_auto_in_d_ready),
    .auto_in_d_valid(widget_auto_in_d_valid),
    .auto_in_d_bits_data(widget_auto_in_d_bits_data),
    .auto_out_a_ready(widget_auto_out_a_ready),
    .auto_out_a_valid(widget_auto_out_a_valid),
    .auto_out_a_bits_opcode(widget_auto_out_a_bits_opcode),
    .auto_out_a_bits_size(widget_auto_out_a_bits_size),
    .auto_out_a_bits_source(widget_auto_out_a_bits_source),
    .auto_out_a_bits_address(widget_auto_out_a_bits_address),
    .auto_out_a_bits_mask(widget_auto_out_a_bits_mask),
    .auto_out_a_bits_data(widget_auto_out_a_bits_data),
    .auto_out_d_ready(widget_auto_out_d_ready),
    .auto_out_d_valid(widget_auto_out_d_valid),
    .auto_out_d_bits_opcode(widget_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(widget_auto_out_d_bits_size),
    .auto_out_d_bits_source(widget_auto_out_d_bits_source),
    .auto_out_d_bits_data(widget_auto_out_d_bits_data)
  );
  Core core ( // @[SoC.scala 40:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_imem_req_ready(core_io_imem_req_ready),
    .io_imem_req_valid(core_io_imem_req_valid),
    .io_imem_req_bits_addr(core_io_imem_req_bits_addr),
    .io_imem_resp_ready(core_io_imem_resp_ready),
    .io_imem_resp_valid(core_io_imem_resp_valid),
    .io_imem_resp_bits_rdata(core_io_imem_resp_bits_rdata),
    .io_dmem_req_ready(core_io_dmem_req_ready),
    .io_dmem_req_valid(core_io_dmem_req_valid),
    .io_dmem_req_bits_addr(core_io_dmem_req_bits_addr),
    .io_dmem_req_bits_wdata(core_io_dmem_req_bits_wdata),
    .io_dmem_req_bits_wmask(core_io_dmem_req_bits_wmask),
    .io_dmem_req_bits_wen(core_io_dmem_req_bits_wen),
    .io_dmem_req_bits_len(core_io_dmem_req_bits_len),
    .io_dmem_req_bits_lrsc(core_io_dmem_req_bits_lrsc),
    .io_dmem_req_bits_amo(core_io_dmem_req_bits_amo),
    .io_dmem_resp_ready(core_io_dmem_resp_ready),
    .io_dmem_resp_valid(core_io_dmem_resp_valid),
    .io_dmem_resp_bits_rdata(core_io_dmem_resp_bits_rdata),
    .io_iptw_req_ready(core_io_iptw_req_ready),
    .io_iptw_req_valid(core_io_iptw_req_valid),
    .io_iptw_req_bits_addr(core_io_iptw_req_bits_addr),
    .io_iptw_resp_ready(core_io_iptw_resp_ready),
    .io_iptw_resp_valid(core_io_iptw_resp_valid),
    .io_iptw_resp_bits_rdata(core_io_iptw_resp_bits_rdata),
    .io_dptw_req_ready(core_io_dptw_req_ready),
    .io_dptw_req_valid(core_io_dptw_req_valid),
    .io_dptw_req_bits_addr(core_io_dptw_req_bits_addr),
    .io_dptw_resp_ready(core_io_dptw_resp_ready),
    .io_dptw_resp_valid(core_io_dptw_resp_valid),
    .io_dptw_resp_bits_rdata(core_io_dptw_resp_bits_rdata),
    .io_uncache_req_ready(core_io_uncache_req_ready),
    .io_uncache_req_valid(core_io_uncache_req_valid),
    .io_uncache_req_bits_addr(core_io_uncache_req_bits_addr),
    .io_uncache_req_bits_wdata(core_io_uncache_req_bits_wdata),
    .io_uncache_req_bits_wmask(core_io_uncache_req_bits_wmask),
    .io_uncache_req_bits_wen(core_io_uncache_req_bits_wen),
    .io_uncache_req_bits_len(core_io_uncache_req_bits_len),
    .io_uncache_resp_ready(core_io_uncache_resp_ready),
    .io_uncache_resp_valid(core_io_uncache_resp_valid),
    .io_uncache_resp_bits_rdata(core_io_uncache_resp_bits_rdata),
    .io_fence_i(core_io_fence_i),
    .io_intr_mtip(core_io_intr_mtip),
    .io_intr_msip(core_io_intr_msip),
    .io_intr_meip(core_io_intr_meip),
    .io_intr_seip(core_io_intr_seip)
  );
  CachePortXBarNto1 xbar_1 ( // @[SoC.scala 50:22]
    .clock(xbar_1_clock),
    .reset(xbar_1_reset),
    .io_in_0_req_ready(xbar_1_io_in_0_req_ready),
    .io_in_0_req_valid(xbar_1_io_in_0_req_valid),
    .io_in_0_req_bits_addr(xbar_1_io_in_0_req_bits_addr),
    .io_in_0_req_bits_wdata(xbar_1_io_in_0_req_bits_wdata),
    .io_in_0_req_bits_wmask(xbar_1_io_in_0_req_bits_wmask),
    .io_in_0_req_bits_wen(xbar_1_io_in_0_req_bits_wen),
    .io_in_0_req_bits_len(xbar_1_io_in_0_req_bits_len),
    .io_in_0_req_bits_lrsc(xbar_1_io_in_0_req_bits_lrsc),
    .io_in_0_req_bits_amo(xbar_1_io_in_0_req_bits_amo),
    .io_in_0_resp_ready(xbar_1_io_in_0_resp_ready),
    .io_in_0_resp_valid(xbar_1_io_in_0_resp_valid),
    .io_in_0_resp_bits_rdata(xbar_1_io_in_0_resp_bits_rdata),
    .io_in_1_req_ready(xbar_1_io_in_1_req_ready),
    .io_in_1_req_valid(xbar_1_io_in_1_req_valid),
    .io_in_1_req_bits_addr(xbar_1_io_in_1_req_bits_addr),
    .io_in_1_resp_ready(xbar_1_io_in_1_resp_ready),
    .io_in_1_resp_valid(xbar_1_io_in_1_resp_valid),
    .io_in_1_resp_bits_rdata(xbar_1_io_in_1_resp_bits_rdata),
    .io_in_2_req_ready(xbar_1_io_in_2_req_ready),
    .io_in_2_req_valid(xbar_1_io_in_2_req_valid),
    .io_in_2_req_bits_addr(xbar_1_io_in_2_req_bits_addr),
    .io_in_2_resp_ready(xbar_1_io_in_2_resp_ready),
    .io_in_2_resp_valid(xbar_1_io_in_2_resp_valid),
    .io_in_2_resp_bits_rdata(xbar_1_io_in_2_resp_bits_rdata),
    .io_out_req_ready(xbar_1_io_out_req_ready),
    .io_out_req_valid(xbar_1_io_out_req_valid),
    .io_out_req_bits_addr(xbar_1_io_out_req_bits_addr),
    .io_out_req_bits_wdata(xbar_1_io_out_req_bits_wdata),
    .io_out_req_bits_wmask(xbar_1_io_out_req_bits_wmask),
    .io_out_req_bits_wen(xbar_1_io_out_req_bits_wen),
    .io_out_req_bits_len(xbar_1_io_out_req_bits_len),
    .io_out_req_bits_lrsc(xbar_1_io_out_req_bits_lrsc),
    .io_out_req_bits_amo(xbar_1_io_out_req_bits_amo),
    .io_out_resp_ready(xbar_1_io_out_resp_ready),
    .io_out_resp_valid(xbar_1_io_out_resp_valid),
    .io_out_resp_bits_rdata(xbar_1_io_out_resp_bits_rdata)
  );
  assign auto_out_a_valid = xbar_auto_out_a_valid; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_out_a_bits_opcode = xbar_auto_out_a_bits_opcode; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_out_a_bits_param = xbar_auto_out_a_bits_param; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_out_a_bits_size = xbar_auto_out_a_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_out_a_bits_source = xbar_auto_out_a_bits_source; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_out_a_bits_address = xbar_auto_out_a_bits_address; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_out_a_bits_mask = xbar_auto_out_a_bits_mask; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_out_a_bits_data = xbar_auto_out_a_bits_data; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_out_b_ready = xbar_auto_out_b_ready; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_out_c_valid = xbar_auto_out_c_valid; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_out_c_bits_opcode = xbar_auto_out_c_bits_opcode; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_out_c_bits_param = xbar_auto_out_c_bits_param; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_out_c_bits_size = xbar_auto_out_c_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_out_c_bits_source = xbar_auto_out_c_bits_source; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_out_c_bits_address = xbar_auto_out_c_bits_address; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_out_c_bits_data = xbar_auto_out_c_bits_data; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_out_d_ready = xbar_auto_out_d_ready; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_out_e_valid = xbar_auto_out_e_valid; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_out_e_bits_sink = xbar_auto_out_e_bits_sink; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign icache_clock = clock;
  assign icache_reset = reset;
  assign icache_auto_out_a_ready = xbar_auto_in_0_a_ready; // @[LazyModule.scala 355:16]
  assign icache_auto_out_d_valid = xbar_auto_in_0_d_valid; // @[LazyModule.scala 355:16]
  assign icache_auto_out_d_bits_data = xbar_auto_in_0_d_bits_data; // @[LazyModule.scala 355:16]
  assign icache_io_cache_req_valid = core_io_imem_req_valid; // @[SoC.scala 46:30]
  assign icache_io_cache_req_bits_addr = core_io_imem_req_bits_addr; // @[SoC.scala 46:30]
  assign icache_io_cache_resp_ready = core_io_imem_resp_ready; // @[SoC.scala 46:30]
  assign icache_io_fence_i = core_io_fence_i; // @[SoC.scala 47:30]
  assign dcache_clock = clock;
  assign dcache_reset = reset;
  assign dcache_auto_out_a_ready = xbar_auto_in_2_a_ready; // @[LazyModule.scala 355:16]
  assign dcache_auto_out_b_valid = xbar_auto_in_2_b_valid; // @[LazyModule.scala 355:16]
  assign dcache_auto_out_b_bits_size = xbar_auto_in_2_b_bits_size; // @[LazyModule.scala 355:16]
  assign dcache_auto_out_b_bits_source = xbar_auto_in_2_b_bits_source; // @[LazyModule.scala 355:16]
  assign dcache_auto_out_b_bits_address = xbar_auto_in_2_b_bits_address; // @[LazyModule.scala 355:16]
  assign dcache_auto_out_c_ready = xbar_auto_in_2_c_ready; // @[LazyModule.scala 355:16]
  assign dcache_auto_out_d_valid = xbar_auto_in_2_d_valid; // @[LazyModule.scala 355:16]
  assign dcache_auto_out_d_bits_sink = xbar_auto_in_2_d_bits_sink; // @[LazyModule.scala 355:16]
  assign dcache_auto_out_d_bits_data = xbar_auto_in_2_d_bits_data; // @[LazyModule.scala 355:16]
  assign dcache_auto_out_e_ready = xbar_auto_in_2_e_ready; // @[LazyModule.scala 355:16]
  assign dcache_io_cache_req_valid = xbar_1_io_out_req_valid; // @[SoC.scala 54:28]
  assign dcache_io_cache_req_bits_addr = xbar_1_io_out_req_bits_addr; // @[SoC.scala 54:28]
  assign dcache_io_cache_req_bits_wdata = xbar_1_io_out_req_bits_wdata; // @[SoC.scala 54:28]
  assign dcache_io_cache_req_bits_wmask = xbar_1_io_out_req_bits_wmask; // @[SoC.scala 54:28]
  assign dcache_io_cache_req_bits_wen = xbar_1_io_out_req_bits_wen; // @[SoC.scala 54:28]
  assign dcache_io_cache_req_bits_len = xbar_1_io_out_req_bits_len; // @[SoC.scala 54:28]
  assign dcache_io_cache_req_bits_lrsc = xbar_1_io_out_req_bits_lrsc; // @[SoC.scala 54:28]
  assign dcache_io_cache_req_bits_amo = xbar_1_io_out_req_bits_amo; // @[SoC.scala 54:28]
  assign dcache_io_cache_resp_ready = xbar_1_io_out_resp_ready; // @[SoC.scala 54:28]
  assign uncache_clock = clock;
  assign uncache_reset = reset;
  assign uncache_auto_out_a_ready = widget_auto_in_a_ready; // @[LazyModule.scala 355:16]
  assign uncache_auto_out_d_valid = widget_auto_in_d_valid; // @[LazyModule.scala 355:16]
  assign uncache_auto_out_d_bits_data = widget_auto_in_d_bits_data; // @[LazyModule.scala 355:16]
  assign uncache_io_in_req_valid = core_io_uncache_req_valid; // @[SoC.scala 57:26]
  assign uncache_io_in_req_bits_addr = core_io_uncache_req_bits_addr; // @[SoC.scala 57:26]
  assign uncache_io_in_req_bits_wdata = core_io_uncache_req_bits_wdata; // @[SoC.scala 57:26]
  assign uncache_io_in_req_bits_wmask = core_io_uncache_req_bits_wmask; // @[SoC.scala 57:26]
  assign uncache_io_in_req_bits_wen = core_io_uncache_req_bits_wen; // @[SoC.scala 57:26]
  assign uncache_io_in_req_bits_len = core_io_uncache_req_bits_len; // @[SoC.scala 57:26]
  assign uncache_io_in_resp_ready = core_io_uncache_resp_ready; // @[SoC.scala 57:26]
  assign xbar_clock = clock;
  assign xbar_reset = reset;
  assign xbar_auto_in_2_a_valid = dcache_auto_out_a_valid; // @[LazyModule.scala 355:16]
  assign xbar_auto_in_2_a_bits_source = dcache_auto_out_a_bits_source; // @[LazyModule.scala 355:16]
  assign xbar_auto_in_2_a_bits_address = dcache_auto_out_a_bits_address; // @[LazyModule.scala 355:16]
  assign xbar_auto_in_2_b_ready = dcache_auto_out_b_ready; // @[LazyModule.scala 355:16]
  assign xbar_auto_in_2_c_valid = dcache_auto_out_c_valid; // @[LazyModule.scala 355:16]
  assign xbar_auto_in_2_c_bits_opcode = dcache_auto_out_c_bits_opcode; // @[LazyModule.scala 355:16]
  assign xbar_auto_in_2_c_bits_param = dcache_auto_out_c_bits_param; // @[LazyModule.scala 355:16]
  assign xbar_auto_in_2_c_bits_size = dcache_auto_out_c_bits_size; // @[LazyModule.scala 355:16]
  assign xbar_auto_in_2_c_bits_source = dcache_auto_out_c_bits_source; // @[LazyModule.scala 355:16]
  assign xbar_auto_in_2_c_bits_address = dcache_auto_out_c_bits_address; // @[LazyModule.scala 355:16]
  assign xbar_auto_in_2_c_bits_data = dcache_auto_out_c_bits_data; // @[LazyModule.scala 355:16]
  assign xbar_auto_in_2_d_ready = dcache_auto_out_d_ready; // @[LazyModule.scala 355:16]
  assign xbar_auto_in_2_e_valid = dcache_auto_out_e_valid; // @[LazyModule.scala 355:16]
  assign xbar_auto_in_2_e_bits_sink = dcache_auto_out_e_bits_sink; // @[LazyModule.scala 355:16]
  assign xbar_auto_in_1_a_valid = widget_auto_out_a_valid; // @[LazyModule.scala 353:16]
  assign xbar_auto_in_1_a_bits_opcode = widget_auto_out_a_bits_opcode; // @[LazyModule.scala 353:16]
  assign xbar_auto_in_1_a_bits_size = widget_auto_out_a_bits_size; // @[LazyModule.scala 353:16]
  assign xbar_auto_in_1_a_bits_source = widget_auto_out_a_bits_source; // @[LazyModule.scala 353:16]
  assign xbar_auto_in_1_a_bits_address = widget_auto_out_a_bits_address; // @[LazyModule.scala 353:16]
  assign xbar_auto_in_1_a_bits_mask = widget_auto_out_a_bits_mask; // @[LazyModule.scala 353:16]
  assign xbar_auto_in_1_a_bits_data = widget_auto_out_a_bits_data; // @[LazyModule.scala 353:16]
  assign xbar_auto_in_1_d_ready = widget_auto_out_d_ready; // @[LazyModule.scala 353:16]
  assign xbar_auto_in_0_a_valid = icache_auto_out_a_valid; // @[LazyModule.scala 355:16]
  assign xbar_auto_in_0_a_bits_source = icache_auto_out_a_bits_source; // @[LazyModule.scala 355:16]
  assign xbar_auto_in_0_a_bits_address = icache_auto_out_a_bits_address; // @[LazyModule.scala 355:16]
  assign xbar_auto_in_0_d_ready = icache_auto_out_d_ready; // @[LazyModule.scala 355:16]
  assign xbar_auto_out_a_ready = auto_out_a_ready; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign xbar_auto_out_b_valid = auto_out_b_valid; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign xbar_auto_out_b_bits_size = auto_out_b_bits_size; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign xbar_auto_out_b_bits_source = auto_out_b_bits_source; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign xbar_auto_out_b_bits_address = auto_out_b_bits_address; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign xbar_auto_out_c_ready = auto_out_c_ready; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign xbar_auto_out_d_valid = auto_out_d_valid; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign xbar_auto_out_d_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign xbar_auto_out_d_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign xbar_auto_out_d_bits_source = auto_out_d_bits_source; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign xbar_auto_out_d_bits_sink = auto_out_d_bits_sink; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign xbar_auto_out_d_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign xbar_auto_out_e_ready = auto_out_e_ready; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign widget_clock = clock;
  assign widget_reset = reset;
  assign widget_auto_in_a_valid = uncache_auto_out_a_valid; // @[LazyModule.scala 355:16]
  assign widget_auto_in_a_bits_opcode = uncache_auto_out_a_bits_opcode; // @[LazyModule.scala 355:16]
  assign widget_auto_in_a_bits_size = uncache_auto_out_a_bits_size; // @[LazyModule.scala 355:16]
  assign widget_auto_in_a_bits_source = uncache_auto_out_a_bits_source; // @[LazyModule.scala 355:16]
  assign widget_auto_in_a_bits_address = uncache_auto_out_a_bits_address; // @[LazyModule.scala 355:16]
  assign widget_auto_in_a_bits_mask = uncache_auto_out_a_bits_mask; // @[LazyModule.scala 355:16]
  assign widget_auto_in_a_bits_data = uncache_auto_out_a_bits_data; // @[LazyModule.scala 355:16]
  assign widget_auto_in_d_ready = uncache_auto_out_d_ready; // @[LazyModule.scala 355:16]
  assign widget_auto_out_a_ready = xbar_auto_in_1_a_ready; // @[LazyModule.scala 353:16]
  assign widget_auto_out_d_valid = xbar_auto_in_1_d_valid; // @[LazyModule.scala 353:16]
  assign widget_auto_out_d_bits_opcode = xbar_auto_in_1_d_bits_opcode; // @[LazyModule.scala 353:16]
  assign widget_auto_out_d_bits_size = xbar_auto_in_1_d_bits_size; // @[LazyModule.scala 353:16]
  assign widget_auto_out_d_bits_source = xbar_auto_in_1_d_bits_source; // @[LazyModule.scala 353:16]
  assign widget_auto_out_d_bits_data = xbar_auto_in_1_d_bits_data; // @[LazyModule.scala 353:16]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_imem_req_ready = icache_io_cache_req_ready; // @[SoC.scala 46:30]
  assign core_io_imem_resp_valid = icache_io_cache_resp_valid; // @[SoC.scala 46:30]
  assign core_io_imem_resp_bits_rdata = icache_io_cache_resp_bits_rdata; // @[SoC.scala 46:30]
  assign core_io_dmem_req_ready = xbar_1_io_in_0_req_ready; // @[SoC.scala 51:28]
  assign core_io_dmem_resp_valid = xbar_1_io_in_0_resp_valid; // @[SoC.scala 51:28]
  assign core_io_dmem_resp_bits_rdata = xbar_1_io_in_0_resp_bits_rdata; // @[SoC.scala 51:28]
  assign core_io_iptw_req_ready = xbar_1_io_in_1_req_ready; // @[SoC.scala 52:28]
  assign core_io_iptw_resp_valid = xbar_1_io_in_1_resp_valid; // @[SoC.scala 52:28]
  assign core_io_iptw_resp_bits_rdata = xbar_1_io_in_1_resp_bits_rdata; // @[SoC.scala 52:28]
  assign core_io_dptw_req_ready = xbar_1_io_in_2_req_ready; // @[SoC.scala 53:28]
  assign core_io_dptw_resp_valid = xbar_1_io_in_2_resp_valid; // @[SoC.scala 53:28]
  assign core_io_dptw_resp_bits_rdata = xbar_1_io_in_2_resp_bits_rdata; // @[SoC.scala 53:28]
  assign core_io_uncache_req_ready = uncache_io_in_req_ready; // @[SoC.scala 57:26]
  assign core_io_uncache_resp_valid = uncache_io_in_resp_valid; // @[SoC.scala 57:26]
  assign core_io_uncache_resp_bits_rdata = uncache_io_in_resp_bits_rdata; // @[SoC.scala 57:26]
  assign core_io_intr_mtip = io_intr_mtip; // @[SoC.scala 43:18]
  assign core_io_intr_msip = io_intr_msip; // @[SoC.scala 43:18]
  assign core_io_intr_meip = io_intr_meip; // @[SoC.scala 43:18]
  assign core_io_intr_seip = io_intr_seip; // @[SoC.scala 43:18]
  assign xbar_1_clock = clock;
  assign xbar_1_reset = reset;
  assign xbar_1_io_in_0_req_valid = core_io_dmem_req_valid; // @[SoC.scala 51:28]
  assign xbar_1_io_in_0_req_bits_addr = core_io_dmem_req_bits_addr; // @[SoC.scala 51:28]
  assign xbar_1_io_in_0_req_bits_wdata = core_io_dmem_req_bits_wdata; // @[SoC.scala 51:28]
  assign xbar_1_io_in_0_req_bits_wmask = core_io_dmem_req_bits_wmask; // @[SoC.scala 51:28]
  assign xbar_1_io_in_0_req_bits_wen = core_io_dmem_req_bits_wen; // @[SoC.scala 51:28]
  assign xbar_1_io_in_0_req_bits_len = core_io_dmem_req_bits_len; // @[SoC.scala 51:28]
  assign xbar_1_io_in_0_req_bits_lrsc = core_io_dmem_req_bits_lrsc; // @[SoC.scala 51:28]
  assign xbar_1_io_in_0_req_bits_amo = core_io_dmem_req_bits_amo; // @[SoC.scala 51:28]
  assign xbar_1_io_in_0_resp_ready = core_io_dmem_resp_ready; // @[SoC.scala 51:28]
  assign xbar_1_io_in_1_req_valid = core_io_iptw_req_valid; // @[SoC.scala 52:28]
  assign xbar_1_io_in_1_req_bits_addr = core_io_iptw_req_bits_addr; // @[SoC.scala 52:28]
  assign xbar_1_io_in_1_resp_ready = core_io_iptw_resp_ready; // @[SoC.scala 52:28]
  assign xbar_1_io_in_2_req_valid = core_io_dptw_req_valid; // @[SoC.scala 53:28]
  assign xbar_1_io_in_2_req_bits_addr = core_io_dptw_req_bits_addr; // @[SoC.scala 53:28]
  assign xbar_1_io_in_2_resp_ready = core_io_dptw_resp_ready; // @[SoC.scala 53:28]
  assign xbar_1_io_out_req_ready = dcache_io_cache_req_ready; // @[SoC.scala 54:28]
  assign xbar_1_io_out_resp_valid = dcache_io_cache_resp_valid; // @[SoC.scala 54:28]
  assign xbar_1_io_out_resp_bits_rdata = dcache_io_cache_resp_bits_rdata; // @[SoC.scala 54:28]
endmodule
module HellaPeekingArbiter(
  input          clock,
  input          reset,
  output         io_in_0_ready,
  input          io_in_0_valid,
  input  [31:0]  io_in_0_bits_union,
  output         io_in_1_ready,
  input          io_in_1_valid,
  input  [2:0]   io_in_1_bits_opcode,
  input  [2:0]   io_in_1_bits_param,
  input  [2:0]   io_in_1_bits_size,
  input  [3:0]   io_in_1_bits_source,
  input  [31:0]  io_in_1_bits_address,
  input  [255:0] io_in_1_bits_data,
  output         io_in_2_ready,
  input          io_in_2_valid,
  input  [2:0]   io_in_2_bits_opcode,
  input  [2:0]   io_in_2_bits_param,
  input  [2:0]   io_in_2_bits_size,
  input  [3:0]   io_in_2_bits_source,
  input  [31:0]  io_in_2_bits_address,
  input  [255:0] io_in_2_bits_data,
  input  [31:0]  io_in_2_bits_union,
  input          io_out_ready,
  output         io_out_valid,
  output [2:0]   io_out_bits_chanId,
  output [2:0]   io_out_bits_opcode,
  output [2:0]   io_out_bits_param,
  output [2:0]   io_out_bits_size,
  output [3:0]   io_out_bits_source,
  output [31:0]  io_out_bits_address,
  output [255:0] io_out_bits_data,
  output [31:0]  io_out_bits_union,
  output         io_out_bits_last
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] lockIdx; // @[Arbiters.scala 26:24]
  reg  locked; // @[Arbiters.scala 27:23]
  wire [1:0] _choice_T = io_in_1_valid ? 2'h1 : 2'h2; // @[Mux.scala 47:70]
  wire [1:0] choice = io_in_0_valid ? 2'h0 : _choice_T; // @[Mux.scala 47:70]
  wire [1:0] chosen = locked ? lockIdx : choice; // @[Arbiters.scala 37:19]
  wire  _GEN_1 = 2'h1 == chosen ? io_in_1_valid : io_in_0_valid; // @[Arbiters.scala 43:{16,16}]
  wire [2:0] _GEN_4 = 2'h1 == chosen ? 3'h2 : 3'h4; // @[Arbiters.scala 44:{15,15}]
  wire [2:0] _GEN_7 = 2'h1 == chosen ? io_in_1_bits_opcode : 3'h0; // @[Arbiters.scala 44:{15,15}]
  wire [2:0] _GEN_10 = 2'h1 == chosen ? io_in_1_bits_param : 3'h0; // @[Arbiters.scala 44:{15,15}]
  wire [2:0] _GEN_13 = 2'h1 == chosen ? io_in_1_bits_size : 3'h0; // @[Arbiters.scala 44:{15,15}]
  wire [3:0] _GEN_16 = 2'h1 == chosen ? io_in_1_bits_source : 4'h0; // @[Arbiters.scala 44:{15,15}]
  wire [31:0] _GEN_19 = 2'h1 == chosen ? io_in_1_bits_address : 32'h0; // @[Arbiters.scala 44:{15,15}]
  wire [255:0] _GEN_22 = 2'h1 == chosen ? io_in_1_bits_data : 256'h0; // @[Arbiters.scala 44:{15,15}]
  wire [31:0] _GEN_28 = 2'h1 == chosen ? 32'h0 : io_in_0_bits_union; // @[Arbiters.scala 44:{15,15}]
  wire  _T = io_out_ready & io_out_valid; // @[Decoupled.scala 51:35]
  wire  _GEN_34 = ~locked | locked; // @[Arbiters.scala 60:50 62:14 27:23]
  assign io_in_0_ready = io_out_ready & chosen == 2'h0; // @[Arbiters.scala 40:36]
  assign io_in_1_ready = io_out_ready & chosen == 2'h1; // @[Arbiters.scala 40:36]
  assign io_in_2_ready = io_out_ready & chosen == 2'h2; // @[Arbiters.scala 40:36]
  assign io_out_valid = 2'h2 == chosen ? io_in_2_valid : _GEN_1; // @[Arbiters.scala 43:{16,16}]
  assign io_out_bits_chanId = 2'h2 == chosen ? 3'h0 : _GEN_4; // @[Arbiters.scala 44:{15,15}]
  assign io_out_bits_opcode = 2'h2 == chosen ? io_in_2_bits_opcode : _GEN_7; // @[Arbiters.scala 44:{15,15}]
  assign io_out_bits_param = 2'h2 == chosen ? io_in_2_bits_param : _GEN_10; // @[Arbiters.scala 44:{15,15}]
  assign io_out_bits_size = 2'h2 == chosen ? io_in_2_bits_size : _GEN_13; // @[Arbiters.scala 44:{15,15}]
  assign io_out_bits_source = 2'h2 == chosen ? io_in_2_bits_source : _GEN_16; // @[Arbiters.scala 44:{15,15}]
  assign io_out_bits_address = 2'h2 == chosen ? io_in_2_bits_address : _GEN_19; // @[Arbiters.scala 44:{15,15}]
  assign io_out_bits_data = 2'h2 == chosen ? io_in_2_bits_data : _GEN_22; // @[Arbiters.scala 44:{15,15}]
  assign io_out_bits_union = 2'h2 == chosen ? io_in_2_bits_union : _GEN_28; // @[Arbiters.scala 44:{15,15}]
  assign io_out_bits_last = 1'h1; // @[Arbiters.scala 44:{15,15}]
  always @(posedge clock) begin
    if (reset) begin // @[Arbiters.scala 26:24]
      lockIdx <= 2'h0; // @[Arbiters.scala 26:24]
    end else if (_T) begin // @[Arbiters.scala 59:22]
      if (~locked) begin // @[Arbiters.scala 60:50]
        if (io_in_0_valid) begin // @[Mux.scala 47:70]
          lockIdx <= 2'h0;
        end else begin
          lockIdx <= _choice_T;
        end
      end
    end
    if (reset) begin // @[Arbiters.scala 27:23]
      locked <= 1'h0; // @[Arbiters.scala 27:23]
    end else if (_T) begin // @[Arbiters.scala 59:22]
      if (io_out_bits_last) begin // @[Arbiters.scala 65:35]
        locked <= 1'h0; // @[Arbiters.scala 66:14]
      end else begin
        locked <= _GEN_34;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lockIdx = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  locked = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module GenericSerializer(
  input          clock,
  input          reset,
  output         io_in_ready,
  input          io_in_valid,
  input  [2:0]   io_in_bits_chanId,
  input  [2:0]   io_in_bits_opcode,
  input  [2:0]   io_in_bits_param,
  input  [2:0]   io_in_bits_size,
  input  [3:0]   io_in_bits_source,
  input  [31:0]  io_in_bits_address,
  input  [255:0] io_in_bits_data,
  input  [31:0]  io_in_bits_union,
  input          io_out_ready,
  output         io_out_valid,
  output [7:0]   io_out_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [351:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [337:0] data; // @[Serdes.scala 173:22]
  reg  sending; // @[Serdes.scala 175:38]
  wire  _T = io_out_ready & io_out_valid; // @[Decoupled.scala 51:35]
  reg [5:0] sendCount; // @[Counter.scala 61:40]
  wire  wrap_wrap = sendCount == 6'h2a; // @[Counter.scala 73:24]
  wire [5:0] _wrap_value_T_1 = sendCount + 6'h1; // @[Counter.scala 77:24]
  wire  sendDone = _T & wrap_wrap; // @[Counter.scala 118:{16,23} 117:24]
  wire  _T_1 = io_in_ready & io_in_valid; // @[Decoupled.scala 51:35]
  wire [337:0] _data_T = {io_in_bits_chanId,io_in_bits_opcode,io_in_bits_param,io_in_bits_size,io_in_bits_source,
    io_in_bits_address,io_in_bits_data,1'h0,io_in_bits_union,1'h1}; // @[Serdes.scala 183:27]
  wire  _GEN_4 = _T_1 | sending; // @[Serdes.scala 182:20 184:13 175:38]
  wire [337:0] _data_T_1 = {{8'd0}, data[337:8]}; // @[Serdes.scala 187:36]
  assign io_in_ready = ~sending; // @[Serdes.scala 178:19]
  assign io_out_valid = sending; // @[Serdes.scala 179:16]
  assign io_out_bits = data[7:0]; // @[Serdes.scala 180:23]
  always @(posedge clock) begin
    if (_T) begin // @[Serdes.scala 187:21]
      data <= _data_T_1; // @[Serdes.scala 187:28]
    end else if (_T_1) begin // @[Serdes.scala 182:20]
      data <= _data_T; // @[Serdes.scala 183:13]
    end
    if (reset) begin // @[Serdes.scala 175:38]
      sending <= 1'h0; // @[Serdes.scala 175:38]
    end else if (sendDone) begin // @[Serdes.scala 189:18]
      sending <= 1'h0; // @[Serdes.scala 189:28]
    end else begin
      sending <= _GEN_4;
    end
    if (reset) begin // @[Counter.scala 61:40]
      sendCount <= 6'h0; // @[Counter.scala 61:40]
    end else if (_T) begin // @[Counter.scala 118:16]
      if (wrap_wrap) begin // @[Counter.scala 87:20]
        sendCount <= 6'h0; // @[Counter.scala 87:28]
      end else begin
        sendCount <= _wrap_value_T_1; // @[Counter.scala 77:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {11{`RANDOM}};
  data = _RAND_0[337:0];
  _RAND_1 = {1{`RANDOM}};
  sending = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  sendCount = _RAND_2[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module GenericDeserializer(
  input          clock,
  input          reset,
  output         io_in_ready,
  input          io_in_valid,
  input  [7:0]   io_in_bits,
  input          io_out_ready,
  output         io_out_valid,
  output [2:0]   io_out_bits_chanId,
  output [2:0]   io_out_bits_opcode,
  output [2:0]   io_out_bits_size,
  output [3:0]   io_out_bits_source,
  output [31:0]  io_out_bits_address,
  output [255:0] io_out_bits_data,
  output [31:0]  io_out_bits_union
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] data_0; // @[Serdes.scala 200:22]
  reg [7:0] data_1; // @[Serdes.scala 200:22]
  reg [7:0] data_2; // @[Serdes.scala 200:22]
  reg [7:0] data_3; // @[Serdes.scala 200:22]
  reg [7:0] data_4; // @[Serdes.scala 200:22]
  reg [7:0] data_5; // @[Serdes.scala 200:22]
  reg [7:0] data_6; // @[Serdes.scala 200:22]
  reg [7:0] data_7; // @[Serdes.scala 200:22]
  reg [7:0] data_8; // @[Serdes.scala 200:22]
  reg [7:0] data_9; // @[Serdes.scala 200:22]
  reg [7:0] data_10; // @[Serdes.scala 200:22]
  reg [7:0] data_11; // @[Serdes.scala 200:22]
  reg [7:0] data_12; // @[Serdes.scala 200:22]
  reg [7:0] data_13; // @[Serdes.scala 200:22]
  reg [7:0] data_14; // @[Serdes.scala 200:22]
  reg [7:0] data_15; // @[Serdes.scala 200:22]
  reg [7:0] data_16; // @[Serdes.scala 200:22]
  reg [7:0] data_17; // @[Serdes.scala 200:22]
  reg [7:0] data_18; // @[Serdes.scala 200:22]
  reg [7:0] data_19; // @[Serdes.scala 200:22]
  reg [7:0] data_20; // @[Serdes.scala 200:22]
  reg [7:0] data_21; // @[Serdes.scala 200:22]
  reg [7:0] data_22; // @[Serdes.scala 200:22]
  reg [7:0] data_23; // @[Serdes.scala 200:22]
  reg [7:0] data_24; // @[Serdes.scala 200:22]
  reg [7:0] data_25; // @[Serdes.scala 200:22]
  reg [7:0] data_26; // @[Serdes.scala 200:22]
  reg [7:0] data_27; // @[Serdes.scala 200:22]
  reg [7:0] data_28; // @[Serdes.scala 200:22]
  reg [7:0] data_29; // @[Serdes.scala 200:22]
  reg [7:0] data_30; // @[Serdes.scala 200:22]
  reg [7:0] data_31; // @[Serdes.scala 200:22]
  reg [7:0] data_32; // @[Serdes.scala 200:22]
  reg [7:0] data_33; // @[Serdes.scala 200:22]
  reg [7:0] data_34; // @[Serdes.scala 200:22]
  reg [7:0] data_35; // @[Serdes.scala 200:22]
  reg [7:0] data_36; // @[Serdes.scala 200:22]
  reg [7:0] data_37; // @[Serdes.scala 200:22]
  reg [7:0] data_38; // @[Serdes.scala 200:22]
  reg [7:0] data_39; // @[Serdes.scala 200:22]
  reg [7:0] data_40; // @[Serdes.scala 200:22]
  reg [7:0] data_41; // @[Serdes.scala 200:22]
  reg [7:0] data_42; // @[Serdes.scala 200:22]
  reg  receiving; // @[Serdes.scala 202:38]
  wire  _T = io_in_ready & io_in_valid; // @[Decoupled.scala 51:35]
  reg [5:0] recvCount; // @[Counter.scala 61:40]
  wire  wrap_wrap = recvCount == 6'h2a; // @[Counter.scala 73:24]
  wire [5:0] _wrap_value_T_1 = recvCount + 6'h1; // @[Counter.scala 77:24]
  wire  recvDone = _T & wrap_wrap; // @[Counter.scala 118:{16,23} 117:24]
  wire [79:0] io_out_bits_lo_lo = {data_9,data_8,data_7,data_6,data_5,data_4,data_3,data_2,data_1,data_0}; // @[Serdes.scala 207:24]
  wire [39:0] io_out_bits_lo_hi_lo = {data_14,data_13,data_12,data_11,data_10}; // @[Serdes.scala 207:24]
  wire [167:0] io_out_bits_lo = {data_20,data_19,data_18,data_17,data_16,data_15,io_out_bits_lo_hi_lo,io_out_bits_lo_lo}
    ; // @[Serdes.scala 207:24]
  wire [39:0] io_out_bits_hi_lo_lo = {data_25,data_24,data_23,data_22,data_21}; // @[Serdes.scala 207:24]
  wire [87:0] io_out_bits_hi_lo = {data_31,data_30,data_29,data_28,data_27,data_26,io_out_bits_hi_lo_lo}; // @[Serdes.scala 207:24]
  wire [39:0] io_out_bits_hi_hi_lo = {data_36,data_35,data_34,data_33,data_32}; // @[Serdes.scala 207:24]
  wire [343:0] _io_out_bits_T = {data_42,data_41,data_40,data_39,data_38,data_37,io_out_bits_hi_hi_lo,io_out_bits_hi_lo,
    io_out_bits_lo}; // @[Serdes.scala 207:24]
  wire  _GEN_89 = recvDone ? 1'h0 : receiving; // @[Serdes.scala 213:{18,30} 202:38]
  wire  _T_2 = io_out_ready & io_out_valid; // @[Decoupled.scala 51:35]
  wire  _GEN_90 = _T_2 | _GEN_89; // @[Serdes.scala 215:{21,33}]
  assign io_in_ready = receiving; // @[Serdes.scala 205:16]
  assign io_out_valid = ~receiving; // @[Serdes.scala 206:19]
  assign io_out_bits_chanId = _io_out_bits_T[337:335]; // @[Serdes.scala 207:39]
  assign io_out_bits_opcode = _io_out_bits_T[334:332]; // @[Serdes.scala 207:39]
  assign io_out_bits_size = _io_out_bits_T[328:326]; // @[Serdes.scala 207:39]
  assign io_out_bits_source = _io_out_bits_T[325:322]; // @[Serdes.scala 207:39]
  assign io_out_bits_address = _io_out_bits_T[321:290]; // @[Serdes.scala 207:39]
  assign io_out_bits_data = _io_out_bits_T[289:34]; // @[Serdes.scala 207:39]
  assign io_out_bits_union = _io_out_bits_T[32:1]; // @[Serdes.scala 207:39]
  always @(posedge clock) begin
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h0 == recvCount) begin // @[Serdes.scala 210:21]
        data_0 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h1 == recvCount) begin // @[Serdes.scala 210:21]
        data_1 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h2 == recvCount) begin // @[Serdes.scala 210:21]
        data_2 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h3 == recvCount) begin // @[Serdes.scala 210:21]
        data_3 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h4 == recvCount) begin // @[Serdes.scala 210:21]
        data_4 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h5 == recvCount) begin // @[Serdes.scala 210:21]
        data_5 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h6 == recvCount) begin // @[Serdes.scala 210:21]
        data_6 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h7 == recvCount) begin // @[Serdes.scala 210:21]
        data_7 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h8 == recvCount) begin // @[Serdes.scala 210:21]
        data_8 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h9 == recvCount) begin // @[Serdes.scala 210:21]
        data_9 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'ha == recvCount) begin // @[Serdes.scala 210:21]
        data_10 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'hb == recvCount) begin // @[Serdes.scala 210:21]
        data_11 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'hc == recvCount) begin // @[Serdes.scala 210:21]
        data_12 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'hd == recvCount) begin // @[Serdes.scala 210:21]
        data_13 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'he == recvCount) begin // @[Serdes.scala 210:21]
        data_14 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'hf == recvCount) begin // @[Serdes.scala 210:21]
        data_15 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h10 == recvCount) begin // @[Serdes.scala 210:21]
        data_16 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h11 == recvCount) begin // @[Serdes.scala 210:21]
        data_17 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h12 == recvCount) begin // @[Serdes.scala 210:21]
        data_18 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h13 == recvCount) begin // @[Serdes.scala 210:21]
        data_19 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h14 == recvCount) begin // @[Serdes.scala 210:21]
        data_20 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h15 == recvCount) begin // @[Serdes.scala 210:21]
        data_21 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h16 == recvCount) begin // @[Serdes.scala 210:21]
        data_22 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h17 == recvCount) begin // @[Serdes.scala 210:21]
        data_23 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h18 == recvCount) begin // @[Serdes.scala 210:21]
        data_24 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h19 == recvCount) begin // @[Serdes.scala 210:21]
        data_25 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h1a == recvCount) begin // @[Serdes.scala 210:21]
        data_26 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h1b == recvCount) begin // @[Serdes.scala 210:21]
        data_27 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h1c == recvCount) begin // @[Serdes.scala 210:21]
        data_28 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h1d == recvCount) begin // @[Serdes.scala 210:21]
        data_29 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h1e == recvCount) begin // @[Serdes.scala 210:21]
        data_30 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h1f == recvCount) begin // @[Serdes.scala 210:21]
        data_31 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h20 == recvCount) begin // @[Serdes.scala 210:21]
        data_32 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h21 == recvCount) begin // @[Serdes.scala 210:21]
        data_33 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h22 == recvCount) begin // @[Serdes.scala 210:21]
        data_34 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h23 == recvCount) begin // @[Serdes.scala 210:21]
        data_35 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h24 == recvCount) begin // @[Serdes.scala 210:21]
        data_36 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h25 == recvCount) begin // @[Serdes.scala 210:21]
        data_37 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h26 == recvCount) begin // @[Serdes.scala 210:21]
        data_38 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h27 == recvCount) begin // @[Serdes.scala 210:21]
        data_39 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h28 == recvCount) begin // @[Serdes.scala 210:21]
        data_40 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h29 == recvCount) begin // @[Serdes.scala 210:21]
        data_41 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h2a == recvCount) begin // @[Serdes.scala 210:21]
        data_42 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    receiving <= reset | _GEN_90; // @[Serdes.scala 202:{38,38}]
    if (reset) begin // @[Counter.scala 61:40]
      recvCount <= 6'h0; // @[Counter.scala 61:40]
    end else if (_T) begin // @[Counter.scala 118:16]
      if (wrap_wrap) begin // @[Counter.scala 87:20]
        recvCount <= 6'h0; // @[Counter.scala 87:28]
      end else begin
        recvCount <= _wrap_value_T_1; // @[Counter.scala 77:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  receiving = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  recvCount = _RAND_44[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLSerdes(
  input          clock,
  input          reset,
  output         auto_in_a_ready,
  input          auto_in_a_valid,
  input  [2:0]   auto_in_a_bits_opcode,
  input  [2:0]   auto_in_a_bits_param,
  input  [2:0]   auto_in_a_bits_size,
  input  [3:0]   auto_in_a_bits_source,
  input  [31:0]  auto_in_a_bits_address,
  input  [31:0]  auto_in_a_bits_mask,
  input  [255:0] auto_in_a_bits_data,
  input          auto_in_b_ready,
  output         auto_in_b_valid,
  output [2:0]   auto_in_b_bits_size,
  output [3:0]   auto_in_b_bits_source,
  output [31:0]  auto_in_b_bits_address,
  output         auto_in_c_ready,
  input          auto_in_c_valid,
  input  [2:0]   auto_in_c_bits_opcode,
  input  [2:0]   auto_in_c_bits_param,
  input  [2:0]   auto_in_c_bits_size,
  input  [3:0]   auto_in_c_bits_source,
  input  [31:0]  auto_in_c_bits_address,
  input  [255:0] auto_in_c_bits_data,
  input          auto_in_d_ready,
  output         auto_in_d_valid,
  output [2:0]   auto_in_d_bits_opcode,
  output [2:0]   auto_in_d_bits_size,
  output [3:0]   auto_in_d_bits_source,
  output [5:0]   auto_in_d_bits_sink,
  output [255:0] auto_in_d_bits_data,
  output         auto_in_e_ready,
  input          auto_in_e_valid,
  input  [5:0]   auto_in_e_bits_sink,
  output         io_ser_0_in_ready,
  input          io_ser_0_in_valid,
  input  [7:0]   io_ser_0_in_bits,
  input          io_ser_0_out_ready,
  output         io_ser_0_out_valid,
  output [7:0]   io_ser_0_out_bits
);
  wire  outArb_clock; // @[Serdes.scala 568:33]
  wire  outArb_reset; // @[Serdes.scala 568:33]
  wire  outArb_io_in_0_ready; // @[Serdes.scala 568:33]
  wire  outArb_io_in_0_valid; // @[Serdes.scala 568:33]
  wire [31:0] outArb_io_in_0_bits_union; // @[Serdes.scala 568:33]
  wire  outArb_io_in_1_ready; // @[Serdes.scala 568:33]
  wire  outArb_io_in_1_valid; // @[Serdes.scala 568:33]
  wire [2:0] outArb_io_in_1_bits_opcode; // @[Serdes.scala 568:33]
  wire [2:0] outArb_io_in_1_bits_param; // @[Serdes.scala 568:33]
  wire [2:0] outArb_io_in_1_bits_size; // @[Serdes.scala 568:33]
  wire [3:0] outArb_io_in_1_bits_source; // @[Serdes.scala 568:33]
  wire [31:0] outArb_io_in_1_bits_address; // @[Serdes.scala 568:33]
  wire [255:0] outArb_io_in_1_bits_data; // @[Serdes.scala 568:33]
  wire  outArb_io_in_2_ready; // @[Serdes.scala 568:33]
  wire  outArb_io_in_2_valid; // @[Serdes.scala 568:33]
  wire [2:0] outArb_io_in_2_bits_opcode; // @[Serdes.scala 568:33]
  wire [2:0] outArb_io_in_2_bits_param; // @[Serdes.scala 568:33]
  wire [2:0] outArb_io_in_2_bits_size; // @[Serdes.scala 568:33]
  wire [3:0] outArb_io_in_2_bits_source; // @[Serdes.scala 568:33]
  wire [31:0] outArb_io_in_2_bits_address; // @[Serdes.scala 568:33]
  wire [255:0] outArb_io_in_2_bits_data; // @[Serdes.scala 568:33]
  wire [31:0] outArb_io_in_2_bits_union; // @[Serdes.scala 568:33]
  wire  outArb_io_out_ready; // @[Serdes.scala 568:33]
  wire  outArb_io_out_valid; // @[Serdes.scala 568:33]
  wire [2:0] outArb_io_out_bits_chanId; // @[Serdes.scala 568:33]
  wire [2:0] outArb_io_out_bits_opcode; // @[Serdes.scala 568:33]
  wire [2:0] outArb_io_out_bits_param; // @[Serdes.scala 568:33]
  wire [2:0] outArb_io_out_bits_size; // @[Serdes.scala 568:33]
  wire [3:0] outArb_io_out_bits_source; // @[Serdes.scala 568:33]
  wire [31:0] outArb_io_out_bits_address; // @[Serdes.scala 568:33]
  wire [255:0] outArb_io_out_bits_data; // @[Serdes.scala 568:33]
  wire [31:0] outArb_io_out_bits_union; // @[Serdes.scala 568:33]
  wire  outArb_io_out_bits_last; // @[Serdes.scala 568:33]
  wire  outSer_clock; // @[Serdes.scala 569:33]
  wire  outSer_reset; // @[Serdes.scala 569:33]
  wire  outSer_io_in_ready; // @[Serdes.scala 569:33]
  wire  outSer_io_in_valid; // @[Serdes.scala 569:33]
  wire [2:0] outSer_io_in_bits_chanId; // @[Serdes.scala 569:33]
  wire [2:0] outSer_io_in_bits_opcode; // @[Serdes.scala 569:33]
  wire [2:0] outSer_io_in_bits_param; // @[Serdes.scala 569:33]
  wire [2:0] outSer_io_in_bits_size; // @[Serdes.scala 569:33]
  wire [3:0] outSer_io_in_bits_source; // @[Serdes.scala 569:33]
  wire [31:0] outSer_io_in_bits_address; // @[Serdes.scala 569:33]
  wire [255:0] outSer_io_in_bits_data; // @[Serdes.scala 569:33]
  wire [31:0] outSer_io_in_bits_union; // @[Serdes.scala 569:33]
  wire  outSer_io_out_ready; // @[Serdes.scala 569:33]
  wire  outSer_io_out_valid; // @[Serdes.scala 569:33]
  wire [7:0] outSer_io_out_bits; // @[Serdes.scala 569:33]
  wire  inDes_clock; // @[Serdes.scala 574:27]
  wire  inDes_reset; // @[Serdes.scala 574:27]
  wire  inDes_io_in_ready; // @[Serdes.scala 574:27]
  wire  inDes_io_in_valid; // @[Serdes.scala 574:27]
  wire [7:0] inDes_io_in_bits; // @[Serdes.scala 574:27]
  wire  inDes_io_out_ready; // @[Serdes.scala 574:27]
  wire  inDes_io_out_valid; // @[Serdes.scala 574:27]
  wire [2:0] inDes_io_out_bits_chanId; // @[Serdes.scala 574:27]
  wire [2:0] inDes_io_out_bits_opcode; // @[Serdes.scala 574:27]
  wire [2:0] inDes_io_out_bits_size; // @[Serdes.scala 574:27]
  wire [3:0] inDes_io_out_bits_source; // @[Serdes.scala 574:27]
  wire [31:0] inDes_io_out_bits_address; // @[Serdes.scala 574:27]
  wire [255:0] inDes_io_out_bits_data; // @[Serdes.scala 574:27]
  wire [31:0] inDes_io_out_bits_union; // @[Serdes.scala 574:27]
  wire [6:0] _outChannels_merged_bits_merged_union_T = {auto_in_e_bits_sink,1'h0}; // @[Cat.scala 33:92]
  wire  _bundleIn_0_b_valid_T = inDes_io_out_bits_chanId == 3'h1; // @[Serdes.scala 235:37]
  wire  _bundleIn_0_d_valid_T = inDes_io_out_bits_chanId == 3'h3; // @[Serdes.scala 237:37]
  wire [31:0] _bundleIn_0_d_bits_d_sink_T = {{1'd0}, inDes_io_out_bits_union[31:1]}; // @[Serdes.scala 486:31]
  HellaPeekingArbiter outArb ( // @[Serdes.scala 568:33]
    .clock(outArb_clock),
    .reset(outArb_reset),
    .io_in_0_ready(outArb_io_in_0_ready),
    .io_in_0_valid(outArb_io_in_0_valid),
    .io_in_0_bits_union(outArb_io_in_0_bits_union),
    .io_in_1_ready(outArb_io_in_1_ready),
    .io_in_1_valid(outArb_io_in_1_valid),
    .io_in_1_bits_opcode(outArb_io_in_1_bits_opcode),
    .io_in_1_bits_param(outArb_io_in_1_bits_param),
    .io_in_1_bits_size(outArb_io_in_1_bits_size),
    .io_in_1_bits_source(outArb_io_in_1_bits_source),
    .io_in_1_bits_address(outArb_io_in_1_bits_address),
    .io_in_1_bits_data(outArb_io_in_1_bits_data),
    .io_in_2_ready(outArb_io_in_2_ready),
    .io_in_2_valid(outArb_io_in_2_valid),
    .io_in_2_bits_opcode(outArb_io_in_2_bits_opcode),
    .io_in_2_bits_param(outArb_io_in_2_bits_param),
    .io_in_2_bits_size(outArb_io_in_2_bits_size),
    .io_in_2_bits_source(outArb_io_in_2_bits_source),
    .io_in_2_bits_address(outArb_io_in_2_bits_address),
    .io_in_2_bits_data(outArb_io_in_2_bits_data),
    .io_in_2_bits_union(outArb_io_in_2_bits_union),
    .io_out_ready(outArb_io_out_ready),
    .io_out_valid(outArb_io_out_valid),
    .io_out_bits_chanId(outArb_io_out_bits_chanId),
    .io_out_bits_opcode(outArb_io_out_bits_opcode),
    .io_out_bits_param(outArb_io_out_bits_param),
    .io_out_bits_size(outArb_io_out_bits_size),
    .io_out_bits_source(outArb_io_out_bits_source),
    .io_out_bits_address(outArb_io_out_bits_address),
    .io_out_bits_data(outArb_io_out_bits_data),
    .io_out_bits_union(outArb_io_out_bits_union),
    .io_out_bits_last(outArb_io_out_bits_last)
  );
  GenericSerializer outSer ( // @[Serdes.scala 569:33]
    .clock(outSer_clock),
    .reset(outSer_reset),
    .io_in_ready(outSer_io_in_ready),
    .io_in_valid(outSer_io_in_valid),
    .io_in_bits_chanId(outSer_io_in_bits_chanId),
    .io_in_bits_opcode(outSer_io_in_bits_opcode),
    .io_in_bits_param(outSer_io_in_bits_param),
    .io_in_bits_size(outSer_io_in_bits_size),
    .io_in_bits_source(outSer_io_in_bits_source),
    .io_in_bits_address(outSer_io_in_bits_address),
    .io_in_bits_data(outSer_io_in_bits_data),
    .io_in_bits_union(outSer_io_in_bits_union),
    .io_out_ready(outSer_io_out_ready),
    .io_out_valid(outSer_io_out_valid),
    .io_out_bits(outSer_io_out_bits)
  );
  GenericDeserializer inDes ( // @[Serdes.scala 574:27]
    .clock(inDes_clock),
    .reset(inDes_reset),
    .io_in_ready(inDes_io_in_ready),
    .io_in_valid(inDes_io_in_valid),
    .io_in_bits(inDes_io_in_bits),
    .io_out_ready(inDes_io_out_ready),
    .io_out_valid(inDes_io_out_valid),
    .io_out_bits_chanId(inDes_io_out_bits_chanId),
    .io_out_bits_opcode(inDes_io_out_bits_opcode),
    .io_out_bits_size(inDes_io_out_bits_size),
    .io_out_bits_source(inDes_io_out_bits_source),
    .io_out_bits_address(inDes_io_out_bits_address),
    .io_out_bits_data(inDes_io_out_bits_data),
    .io_out_bits_union(inDes_io_out_bits_union)
  );
  assign auto_in_a_ready = outArb_io_in_2_ready; // @[Serdes.scala 363:22 570:22]
  assign auto_in_b_valid = inDes_io_out_valid & _bundleIn_0_b_valid_T; // @[Serdes.scala 576:43]
  assign auto_in_b_bits_size = inDes_io_out_bits_size; // @[Serdes.scala 413:17 416:15]
  assign auto_in_b_bits_source = inDes_io_out_bits_source; // @[Serdes.scala 413:17 417:15]
  assign auto_in_b_bits_address = inDes_io_out_bits_address; // @[Serdes.scala 413:17 418:15]
  assign auto_in_c_ready = outArb_io_in_1_ready; // @[Serdes.scala 363:22 570:22]
  assign auto_in_d_valid = inDes_io_out_valid & _bundleIn_0_d_valid_T; // @[Serdes.scala 578:43]
  assign auto_in_d_bits_opcode = inDes_io_out_bits_opcode; // @[Serdes.scala 478:17 479:14]
  assign auto_in_d_bits_size = inDes_io_out_bits_size; // @[Serdes.scala 478:17 481:14]
  assign auto_in_d_bits_source = inDes_io_out_bits_source; // @[Serdes.scala 478:17 482:14]
  assign auto_in_d_bits_sink = _bundleIn_0_d_bits_d_sink_T[5:0]; // @[Serdes.scala 478:17 486:17]
  assign auto_in_d_bits_data = inDes_io_out_bits_data; // @[Serdes.scala 478:17 483:14]
  assign auto_in_e_ready = outArb_io_in_0_ready; // @[Serdes.scala 363:22 570:22]
  assign io_ser_0_in_ready = inDes_io_in_ready; // @[Serdes.scala 575:21]
  assign io_ser_0_out_valid = outSer_io_out_valid; // @[Serdes.scala 572:22]
  assign io_ser_0_out_bits = outSer_io_out_bits; // @[Serdes.scala 572:22]
  assign outArb_clock = clock;
  assign outArb_reset = reset;
  assign outArb_io_in_0_valid = auto_in_e_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign outArb_io_in_0_bits_union = {{25'd0}, _outChannels_merged_bits_merged_union_T}; // @[Serdes.scala 330:22 340:26]
  assign outArb_io_in_1_valid = auto_in_c_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign outArb_io_in_1_bits_opcode = auto_in_c_bits_opcode; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign outArb_io_in_1_bits_param = auto_in_c_bits_param; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign outArb_io_in_1_bits_size = auto_in_c_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign outArb_io_in_1_bits_source = auto_in_c_bits_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign outArb_io_in_1_bits_address = auto_in_c_bits_address; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign outArb_io_in_1_bits_data = auto_in_c_bits_data; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign outArb_io_in_2_valid = auto_in_a_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign outArb_io_in_2_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign outArb_io_in_2_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign outArb_io_in_2_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign outArb_io_in_2_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign outArb_io_in_2_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign outArb_io_in_2_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign outArb_io_in_2_bits_union = auto_in_a_bits_mask; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign outArb_io_out_ready = outSer_io_in_ready; // @[Serdes.scala 571:22]
  assign outSer_clock = clock;
  assign outSer_reset = reset;
  assign outSer_io_in_valid = outArb_io_out_valid; // @[Serdes.scala 571:22]
  assign outSer_io_in_bits_chanId = outArb_io_out_bits_chanId; // @[Serdes.scala 571:22]
  assign outSer_io_in_bits_opcode = outArb_io_out_bits_opcode; // @[Serdes.scala 571:22]
  assign outSer_io_in_bits_param = outArb_io_out_bits_param; // @[Serdes.scala 571:22]
  assign outSer_io_in_bits_size = outArb_io_out_bits_size; // @[Serdes.scala 571:22]
  assign outSer_io_in_bits_source = outArb_io_out_bits_source; // @[Serdes.scala 571:22]
  assign outSer_io_in_bits_address = outArb_io_out_bits_address; // @[Serdes.scala 571:22]
  assign outSer_io_in_bits_data = outArb_io_out_bits_data; // @[Serdes.scala 571:22]
  assign outSer_io_in_bits_union = outArb_io_out_bits_union; // @[Serdes.scala 571:22]
  assign outSer_io_out_ready = io_ser_0_out_ready; // @[Serdes.scala 572:22]
  assign inDes_clock = clock;
  assign inDes_reset = reset;
  assign inDes_io_in_valid = io_ser_0_in_valid; // @[Serdes.scala 575:21]
  assign inDes_io_in_bits = io_ser_0_in_bits; // @[Serdes.scala 575:21]
  assign inDes_io_out_ready = 3'h3 == inDes_io_out_bits_chanId ? auto_in_d_ready : 3'h1 == inDes_io_out_bits_chanId &
    auto_in_b_ready; // @[Mux.scala 81:58]
endmodule
module TLTraceBuffer(
  input          clock,
  input          reset,
  output         auto_in_a_ready,
  input          auto_in_a_valid,
  input  [2:0]   auto_in_a_bits_opcode,
  input  [2:0]   auto_in_a_bits_param,
  input  [2:0]   auto_in_a_bits_size,
  input  [3:0]   auto_in_a_bits_source,
  input  [31:0]  auto_in_a_bits_address,
  input  [31:0]  auto_in_a_bits_mask,
  input  [255:0] auto_in_a_bits_data,
  input          auto_in_b_ready,
  output         auto_in_b_valid,
  output [2:0]   auto_in_b_bits_size,
  output [3:0]   auto_in_b_bits_source,
  output [31:0]  auto_in_b_bits_address,
  output         auto_in_c_ready,
  input          auto_in_c_valid,
  input  [2:0]   auto_in_c_bits_opcode,
  input  [2:0]   auto_in_c_bits_param,
  input  [2:0]   auto_in_c_bits_size,
  input  [3:0]   auto_in_c_bits_source,
  input  [31:0]  auto_in_c_bits_address,
  input  [255:0] auto_in_c_bits_data,
  input          auto_in_d_ready,
  output         auto_in_d_valid,
  output [2:0]   auto_in_d_bits_opcode,
  output [2:0]   auto_in_d_bits_size,
  output [3:0]   auto_in_d_bits_source,
  output [5:0]   auto_in_d_bits_sink,
  output [255:0] auto_in_d_bits_data,
  output         auto_in_e_ready,
  input          auto_in_e_valid,
  input  [5:0]   auto_in_e_bits_sink,
  input          auto_out_a_ready,
  output         auto_out_a_valid,
  output [2:0]   auto_out_a_bits_opcode,
  output [2:0]   auto_out_a_bits_param,
  output [2:0]   auto_out_a_bits_size,
  output [3:0]   auto_out_a_bits_source,
  output [31:0]  auto_out_a_bits_address,
  output [31:0]  auto_out_a_bits_mask,
  output [255:0] auto_out_a_bits_data,
  output         auto_out_b_ready,
  input          auto_out_b_valid,
  input  [2:0]   auto_out_b_bits_size,
  input  [3:0]   auto_out_b_bits_source,
  input  [31:0]  auto_out_b_bits_address,
  input          auto_out_c_ready,
  output         auto_out_c_valid,
  output [2:0]   auto_out_c_bits_opcode,
  output [2:0]   auto_out_c_bits_param,
  output [2:0]   auto_out_c_bits_size,
  output [3:0]   auto_out_c_bits_source,
  output [31:0]  auto_out_c_bits_address,
  output [255:0] auto_out_c_bits_data,
  output         auto_out_d_ready,
  input          auto_out_d_valid,
  input  [2:0]   auto_out_d_bits_opcode,
  input  [2:0]   auto_out_d_bits_size,
  input  [3:0]   auto_out_d_bits_source,
  input  [5:0]   auto_out_d_bits_sink,
  input  [255:0] auto_out_d_bits_data,
  input          auto_out_e_ready,
  output         auto_out_e_valid,
  output [5:0]   auto_out_e_bits_sink
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [255:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [255:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [255:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
`endif // RANDOMIZE_REG_INIT
  reg  in_a_scan_valid; // @[Utils.scala 36:20]
  wire  _x1_a_ready_T_1 = auto_out_a_ready & in_a_scan_valid; // @[Decoupled.scala 51:35]
  wire  tl_in_a_ready = ~in_a_scan_valid | _x1_a_ready_T_1; // @[TLTraceBuffer.scala 30:38]
  wire  _in_a_scan_bits_T = tl_in_a_ready & auto_in_a_valid; // @[Decoupled.scala 51:35]
  reg [2:0] in_a_scan_bits_opcode; // @[Reg.scala 35:20]
  reg [2:0] in_a_scan_bits_param; // @[Reg.scala 35:20]
  reg [2:0] in_a_scan_bits_size; // @[Reg.scala 35:20]
  reg [3:0] in_a_scan_bits_source; // @[Reg.scala 35:20]
  reg [31:0] in_a_scan_bits_address; // @[Reg.scala 35:20]
  reg [31:0] in_a_scan_bits_mask; // @[Reg.scala 35:20]
  reg [255:0] in_a_scan_bits_data; // @[Reg.scala 35:20]
  wire  _GEN_8 = _x1_a_ready_T_1 ? 1'h0 : in_a_scan_valid; // @[Utils.scala 38:18 36:20 38:22]
  wire  _GEN_9 = _in_a_scan_bits_T | _GEN_8; // @[Utils.scala 39:{19,23}]
  reg  out_b_scan_valid; // @[Utils.scala 36:20]
  wire  _x1_b_ready_T_1 = auto_in_b_ready & out_b_scan_valid; // @[Decoupled.scala 51:35]
  wire  tl_out_b_ready = ~out_b_scan_valid | _x1_b_ready_T_1; // @[TLTraceBuffer.scala 33:39]
  wire  _out_b_scan_bits_T = tl_out_b_ready & auto_out_b_valid; // @[Decoupled.scala 51:35]
  reg [2:0] out_b_scan_bits_size; // @[Reg.scala 35:20]
  reg [3:0] out_b_scan_bits_source; // @[Reg.scala 35:20]
  reg [31:0] out_b_scan_bits_address; // @[Reg.scala 35:20]
  wire  _GEN_18 = _x1_b_ready_T_1 ? 1'h0 : out_b_scan_valid; // @[Utils.scala 38:18 36:20 38:22]
  wire  _GEN_19 = _out_b_scan_bits_T | _GEN_18; // @[Utils.scala 39:{19,23}]
  reg  in_c_scan_valid; // @[Utils.scala 36:20]
  wire  _x1_c_ready_T_1 = auto_out_c_ready & in_c_scan_valid; // @[Decoupled.scala 51:35]
  wire  tl_in_c_ready = ~in_c_scan_valid | _x1_c_ready_T_1; // @[TLTraceBuffer.scala 36:38]
  wire  _in_c_scan_bits_T = tl_in_c_ready & auto_in_c_valid; // @[Decoupled.scala 51:35]
  reg [2:0] in_c_scan_bits_opcode; // @[Reg.scala 35:20]
  reg [2:0] in_c_scan_bits_param; // @[Reg.scala 35:20]
  reg [2:0] in_c_scan_bits_size; // @[Reg.scala 35:20]
  reg [3:0] in_c_scan_bits_source; // @[Reg.scala 35:20]
  reg [31:0] in_c_scan_bits_address; // @[Reg.scala 35:20]
  reg [255:0] in_c_scan_bits_data; // @[Reg.scala 35:20]
  wire  _GEN_27 = _x1_c_ready_T_1 ? 1'h0 : in_c_scan_valid; // @[Utils.scala 38:18 36:20 38:22]
  wire  _GEN_28 = _in_c_scan_bits_T | _GEN_27; // @[Utils.scala 39:{19,23}]
  reg  out_d_scan_valid; // @[Utils.scala 36:20]
  wire  _x1_d_ready_T_1 = auto_in_d_ready & out_d_scan_valid; // @[Decoupled.scala 51:35]
  wire  tl_out_d_ready = ~out_d_scan_valid | _x1_d_ready_T_1; // @[TLTraceBuffer.scala 39:39]
  wire  _out_d_scan_bits_T = tl_out_d_ready & auto_out_d_valid; // @[Decoupled.scala 51:35]
  reg [2:0] out_d_scan_bits_opcode; // @[Reg.scala 35:20]
  reg [2:0] out_d_scan_bits_size; // @[Reg.scala 35:20]
  reg [3:0] out_d_scan_bits_source; // @[Reg.scala 35:20]
  reg [5:0] out_d_scan_bits_sink; // @[Reg.scala 35:20]
  reg [255:0] out_d_scan_bits_data; // @[Reg.scala 35:20]
  wire  _GEN_37 = _x1_d_ready_T_1 ? 1'h0 : out_d_scan_valid; // @[Utils.scala 38:18 36:20 38:22]
  wire  _GEN_38 = _out_d_scan_bits_T | _GEN_37; // @[Utils.scala 39:{19,23}]
  reg  in_e_scan_valid; // @[Utils.scala 36:20]
  wire  _x1_e_ready_T_1 = auto_out_e_ready & in_e_scan_valid; // @[Decoupled.scala 51:35]
  wire  tl_in_e_ready = ~in_e_scan_valid | _x1_e_ready_T_1; // @[TLTraceBuffer.scala 42:38]
  wire  _in_e_scan_bits_T = tl_in_e_ready & auto_in_e_valid; // @[Decoupled.scala 51:35]
  reg [5:0] in_e_scan_bits_sink; // @[Reg.scala 35:20]
  wire  _GEN_40 = _x1_e_ready_T_1 ? 1'h0 : in_e_scan_valid; // @[Utils.scala 38:18 36:20 38:22]
  wire  _GEN_41 = _in_e_scan_bits_T | _GEN_40; // @[Utils.scala 39:{19,23}]
  assign auto_in_a_ready = ~in_a_scan_valid | _x1_a_ready_T_1; // @[TLTraceBuffer.scala 30:38]
  assign auto_in_b_valid = out_b_scan_valid; // @[Nodes.scala 1215:84 TLTraceBuffer.scala 31:18]
  assign auto_in_b_bits_size = out_b_scan_bits_size; // @[Nodes.scala 1215:84 TLTraceBuffer.scala 32:18]
  assign auto_in_b_bits_source = out_b_scan_bits_source; // @[Nodes.scala 1215:84 TLTraceBuffer.scala 32:18]
  assign auto_in_b_bits_address = out_b_scan_bits_address; // @[Nodes.scala 1215:84 TLTraceBuffer.scala 32:18]
  assign auto_in_c_ready = ~in_c_scan_valid | _x1_c_ready_T_1; // @[TLTraceBuffer.scala 36:38]
  assign auto_in_d_valid = out_d_scan_valid; // @[Nodes.scala 1215:84 TLTraceBuffer.scala 37:18]
  assign auto_in_d_bits_opcode = out_d_scan_bits_opcode; // @[Nodes.scala 1215:84 TLTraceBuffer.scala 38:18]
  assign auto_in_d_bits_size = out_d_scan_bits_size; // @[Nodes.scala 1215:84 TLTraceBuffer.scala 38:18]
  assign auto_in_d_bits_source = out_d_scan_bits_source; // @[Nodes.scala 1215:84 TLTraceBuffer.scala 38:18]
  assign auto_in_d_bits_sink = out_d_scan_bits_sink; // @[Nodes.scala 1215:84 TLTraceBuffer.scala 38:18]
  assign auto_in_d_bits_data = out_d_scan_bits_data; // @[Nodes.scala 1215:84 TLTraceBuffer.scala 38:18]
  assign auto_in_e_ready = ~in_e_scan_valid | _x1_e_ready_T_1; // @[TLTraceBuffer.scala 42:38]
  assign auto_out_a_valid = in_a_scan_valid; // @[Nodes.scala 1212:84 TLTraceBuffer.scala 28:18]
  assign auto_out_a_bits_opcode = in_a_scan_bits_opcode; // @[Nodes.scala 1212:84 TLTraceBuffer.scala 29:18]
  assign auto_out_a_bits_param = in_a_scan_bits_param; // @[Nodes.scala 1212:84 TLTraceBuffer.scala 29:18]
  assign auto_out_a_bits_size = in_a_scan_bits_size; // @[Nodes.scala 1212:84 TLTraceBuffer.scala 29:18]
  assign auto_out_a_bits_source = in_a_scan_bits_source; // @[Nodes.scala 1212:84 TLTraceBuffer.scala 29:18]
  assign auto_out_a_bits_address = in_a_scan_bits_address; // @[Nodes.scala 1212:84 TLTraceBuffer.scala 29:18]
  assign auto_out_a_bits_mask = in_a_scan_bits_mask; // @[Nodes.scala 1212:84 TLTraceBuffer.scala 29:18]
  assign auto_out_a_bits_data = in_a_scan_bits_data; // @[Nodes.scala 1212:84 TLTraceBuffer.scala 29:18]
  assign auto_out_b_ready = ~out_b_scan_valid | _x1_b_ready_T_1; // @[TLTraceBuffer.scala 33:39]
  assign auto_out_c_valid = in_c_scan_valid; // @[Nodes.scala 1212:84 TLTraceBuffer.scala 34:18]
  assign auto_out_c_bits_opcode = in_c_scan_bits_opcode; // @[Nodes.scala 1212:84 TLTraceBuffer.scala 35:18]
  assign auto_out_c_bits_param = in_c_scan_bits_param; // @[Nodes.scala 1212:84 TLTraceBuffer.scala 35:18]
  assign auto_out_c_bits_size = in_c_scan_bits_size; // @[Nodes.scala 1212:84 TLTraceBuffer.scala 35:18]
  assign auto_out_c_bits_source = in_c_scan_bits_source; // @[Nodes.scala 1212:84 TLTraceBuffer.scala 35:18]
  assign auto_out_c_bits_address = in_c_scan_bits_address; // @[Nodes.scala 1212:84 TLTraceBuffer.scala 35:18]
  assign auto_out_c_bits_data = in_c_scan_bits_data; // @[Nodes.scala 1212:84 TLTraceBuffer.scala 35:18]
  assign auto_out_d_ready = ~out_d_scan_valid | _x1_d_ready_T_1; // @[TLTraceBuffer.scala 39:39]
  assign auto_out_e_valid = in_e_scan_valid; // @[Nodes.scala 1212:84 TLTraceBuffer.scala 40:18]
  assign auto_out_e_bits_sink = in_e_scan_bits_sink; // @[Nodes.scala 1212:84 TLTraceBuffer.scala 41:18]
  always @(posedge clock) begin
    if (reset) begin // @[Utils.scala 36:20]
      in_a_scan_valid <= 1'h0; // @[Utils.scala 36:20]
    end else begin
      in_a_scan_valid <= _GEN_9;
    end
    if (reset) begin // @[Reg.scala 35:20]
      in_a_scan_bits_opcode <= 3'h0; // @[Reg.scala 35:20]
    end else if (_in_a_scan_bits_T) begin // @[Reg.scala 36:18]
      in_a_scan_bits_opcode <= auto_in_a_bits_opcode; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      in_a_scan_bits_param <= 3'h0; // @[Reg.scala 35:20]
    end else if (_in_a_scan_bits_T) begin // @[Reg.scala 36:18]
      in_a_scan_bits_param <= auto_in_a_bits_param; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      in_a_scan_bits_size <= 3'h0; // @[Reg.scala 35:20]
    end else if (_in_a_scan_bits_T) begin // @[Reg.scala 36:18]
      in_a_scan_bits_size <= auto_in_a_bits_size; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      in_a_scan_bits_source <= 4'h0; // @[Reg.scala 35:20]
    end else if (_in_a_scan_bits_T) begin // @[Reg.scala 36:18]
      in_a_scan_bits_source <= auto_in_a_bits_source; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      in_a_scan_bits_address <= 32'h0; // @[Reg.scala 35:20]
    end else if (_in_a_scan_bits_T) begin // @[Reg.scala 36:18]
      in_a_scan_bits_address <= auto_in_a_bits_address; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      in_a_scan_bits_mask <= 32'h0; // @[Reg.scala 35:20]
    end else if (_in_a_scan_bits_T) begin // @[Reg.scala 36:18]
      in_a_scan_bits_mask <= auto_in_a_bits_mask; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      in_a_scan_bits_data <= 256'h0; // @[Reg.scala 35:20]
    end else if (_in_a_scan_bits_T) begin // @[Reg.scala 36:18]
      in_a_scan_bits_data <= auto_in_a_bits_data; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Utils.scala 36:20]
      out_b_scan_valid <= 1'h0; // @[Utils.scala 36:20]
    end else begin
      out_b_scan_valid <= _GEN_19;
    end
    if (reset) begin // @[Reg.scala 35:20]
      out_b_scan_bits_size <= 3'h0; // @[Reg.scala 35:20]
    end else if (_out_b_scan_bits_T) begin // @[Reg.scala 36:18]
      out_b_scan_bits_size <= auto_out_b_bits_size; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      out_b_scan_bits_source <= 4'h0; // @[Reg.scala 35:20]
    end else if (_out_b_scan_bits_T) begin // @[Reg.scala 36:18]
      out_b_scan_bits_source <= auto_out_b_bits_source; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      out_b_scan_bits_address <= 32'h0; // @[Reg.scala 35:20]
    end else if (_out_b_scan_bits_T) begin // @[Reg.scala 36:18]
      out_b_scan_bits_address <= auto_out_b_bits_address; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Utils.scala 36:20]
      in_c_scan_valid <= 1'h0; // @[Utils.scala 36:20]
    end else begin
      in_c_scan_valid <= _GEN_28;
    end
    if (reset) begin // @[Reg.scala 35:20]
      in_c_scan_bits_opcode <= 3'h0; // @[Reg.scala 35:20]
    end else if (_in_c_scan_bits_T) begin // @[Reg.scala 36:18]
      in_c_scan_bits_opcode <= auto_in_c_bits_opcode; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      in_c_scan_bits_param <= 3'h0; // @[Reg.scala 35:20]
    end else if (_in_c_scan_bits_T) begin // @[Reg.scala 36:18]
      in_c_scan_bits_param <= auto_in_c_bits_param; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      in_c_scan_bits_size <= 3'h0; // @[Reg.scala 35:20]
    end else if (_in_c_scan_bits_T) begin // @[Reg.scala 36:18]
      in_c_scan_bits_size <= auto_in_c_bits_size; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      in_c_scan_bits_source <= 4'h0; // @[Reg.scala 35:20]
    end else if (_in_c_scan_bits_T) begin // @[Reg.scala 36:18]
      in_c_scan_bits_source <= auto_in_c_bits_source; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      in_c_scan_bits_address <= 32'h0; // @[Reg.scala 35:20]
    end else if (_in_c_scan_bits_T) begin // @[Reg.scala 36:18]
      in_c_scan_bits_address <= auto_in_c_bits_address; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      in_c_scan_bits_data <= 256'h0; // @[Reg.scala 35:20]
    end else if (_in_c_scan_bits_T) begin // @[Reg.scala 36:18]
      in_c_scan_bits_data <= auto_in_c_bits_data; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Utils.scala 36:20]
      out_d_scan_valid <= 1'h0; // @[Utils.scala 36:20]
    end else begin
      out_d_scan_valid <= _GEN_38;
    end
    if (reset) begin // @[Reg.scala 35:20]
      out_d_scan_bits_opcode <= 3'h0; // @[Reg.scala 35:20]
    end else if (_out_d_scan_bits_T) begin // @[Reg.scala 36:18]
      out_d_scan_bits_opcode <= auto_out_d_bits_opcode; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      out_d_scan_bits_size <= 3'h0; // @[Reg.scala 35:20]
    end else if (_out_d_scan_bits_T) begin // @[Reg.scala 36:18]
      out_d_scan_bits_size <= auto_out_d_bits_size; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      out_d_scan_bits_source <= 4'h0; // @[Reg.scala 35:20]
    end else if (_out_d_scan_bits_T) begin // @[Reg.scala 36:18]
      out_d_scan_bits_source <= auto_out_d_bits_source; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      out_d_scan_bits_sink <= 6'h0; // @[Reg.scala 35:20]
    end else if (_out_d_scan_bits_T) begin // @[Reg.scala 36:18]
      out_d_scan_bits_sink <= auto_out_d_bits_sink; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      out_d_scan_bits_data <= 256'h0; // @[Reg.scala 35:20]
    end else if (_out_d_scan_bits_T) begin // @[Reg.scala 36:18]
      out_d_scan_bits_data <= auto_out_d_bits_data; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Utils.scala 36:20]
      in_e_scan_valid <= 1'h0; // @[Utils.scala 36:20]
    end else begin
      in_e_scan_valid <= _GEN_41;
    end
    if (reset) begin // @[Reg.scala 35:20]
      in_e_scan_bits_sink <= 6'h0; // @[Reg.scala 35:20]
    end else if (_in_e_scan_bits_T) begin // @[Reg.scala 36:18]
      in_e_scan_bits_sink <= auto_in_e_bits_sink; // @[Reg.scala 36:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  in_a_scan_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  in_a_scan_bits_opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  in_a_scan_bits_param = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  in_a_scan_bits_size = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  in_a_scan_bits_source = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  in_a_scan_bits_address = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  in_a_scan_bits_mask = _RAND_6[31:0];
  _RAND_7 = {8{`RANDOM}};
  in_a_scan_bits_data = _RAND_7[255:0];
  _RAND_8 = {1{`RANDOM}};
  out_b_scan_valid = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  out_b_scan_bits_size = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  out_b_scan_bits_source = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  out_b_scan_bits_address = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  in_c_scan_valid = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  in_c_scan_bits_opcode = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  in_c_scan_bits_param = _RAND_14[2:0];
  _RAND_15 = {1{`RANDOM}};
  in_c_scan_bits_size = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  in_c_scan_bits_source = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
  in_c_scan_bits_address = _RAND_17[31:0];
  _RAND_18 = {8{`RANDOM}};
  in_c_scan_bits_data = _RAND_18[255:0];
  _RAND_19 = {1{`RANDOM}};
  out_d_scan_valid = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  out_d_scan_bits_opcode = _RAND_20[2:0];
  _RAND_21 = {1{`RANDOM}};
  out_d_scan_bits_size = _RAND_21[2:0];
  _RAND_22 = {1{`RANDOM}};
  out_d_scan_bits_source = _RAND_22[3:0];
  _RAND_23 = {1{`RANDOM}};
  out_d_scan_bits_sink = _RAND_23[5:0];
  _RAND_24 = {8{`RANDOM}};
  out_d_scan_bits_data = _RAND_24[255:0];
  _RAND_25 = {1{`RANDOM}};
  in_e_scan_valid = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  in_e_scan_bits_sink = _RAND_26[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AsyncResetSynchronizerPrimitiveShiftReg_d3_i0(
  input   clock,
  input   reset,
  input   io_d,
  output  io_q
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg  sync_0; // @[SynchronizerReg.scala 51:87]
  reg  sync_1; // @[SynchronizerReg.scala 51:87]
  reg  sync_2; // @[SynchronizerReg.scala 51:87]
  assign io_q = sync_0; // @[SynchronizerReg.scala 59:8]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SynchronizerReg.scala 51:87]
      sync_0 <= 1'h0; // @[SynchronizerReg.scala 51:87]
    end else begin
      sync_0 <= sync_1; // @[SynchronizerReg.scala 57:10]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SynchronizerReg.scala 51:87]
      sync_1 <= 1'h0; // @[SynchronizerReg.scala 51:87]
    end else begin
      sync_1 <= sync_2; // @[SynchronizerReg.scala 57:10]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SynchronizerReg.scala 54:22]
      sync_2 <= 1'h0;
    end else begin
      sync_2 <= io_d;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sync_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  sync_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  sync_2 = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    sync_0 = 1'h0;
  end
  if (reset) begin
    sync_1 = 1'h0;
  end
  if (reset) begin
    sync_2 = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AsyncResetSynchronizerShiftReg_w4_d3_i0(
  input        clock,
  input        reset,
  input  [3:0] io_d,
  output [3:0] io_q
);
  wire  output_chain_clock; // @[ShiftReg.scala 45:23]
  wire  output_chain_reset; // @[ShiftReg.scala 45:23]
  wire  output_chain_io_d; // @[ShiftReg.scala 45:23]
  wire  output_chain_io_q; // @[ShiftReg.scala 45:23]
  wire  output_chain_1_clock; // @[ShiftReg.scala 45:23]
  wire  output_chain_1_reset; // @[ShiftReg.scala 45:23]
  wire  output_chain_1_io_d; // @[ShiftReg.scala 45:23]
  wire  output_chain_1_io_q; // @[ShiftReg.scala 45:23]
  wire  output_chain_2_clock; // @[ShiftReg.scala 45:23]
  wire  output_chain_2_reset; // @[ShiftReg.scala 45:23]
  wire  output_chain_2_io_d; // @[ShiftReg.scala 45:23]
  wire  output_chain_2_io_q; // @[ShiftReg.scala 45:23]
  wire  output_chain_3_clock; // @[ShiftReg.scala 45:23]
  wire  output_chain_3_reset; // @[ShiftReg.scala 45:23]
  wire  output_chain_3_io_d; // @[ShiftReg.scala 45:23]
  wire  output_chain_3_io_q; // @[ShiftReg.scala 45:23]
  wire  output_1 = output_chain_1_io_q; // @[ShiftReg.scala 48:{24,24}]
  wire  output_0 = output_chain_io_q; // @[ShiftReg.scala 48:{24,24}]
  wire [1:0] io_q_lo = {output_1,output_0}; // @[Cat.scala 33:92]
  wire  output_3 = output_chain_3_io_q; // @[ShiftReg.scala 48:{24,24}]
  wire  output_2 = output_chain_2_io_q; // @[ShiftReg.scala 48:{24,24}]
  wire [1:0] io_q_hi = {output_3,output_2}; // @[Cat.scala 33:92]
  AsyncResetSynchronizerPrimitiveShiftReg_d3_i0 output_chain ( // @[ShiftReg.scala 45:23]
    .clock(output_chain_clock),
    .reset(output_chain_reset),
    .io_d(output_chain_io_d),
    .io_q(output_chain_io_q)
  );
  AsyncResetSynchronizerPrimitiveShiftReg_d3_i0 output_chain_1 ( // @[ShiftReg.scala 45:23]
    .clock(output_chain_1_clock),
    .reset(output_chain_1_reset),
    .io_d(output_chain_1_io_d),
    .io_q(output_chain_1_io_q)
  );
  AsyncResetSynchronizerPrimitiveShiftReg_d3_i0 output_chain_2 ( // @[ShiftReg.scala 45:23]
    .clock(output_chain_2_clock),
    .reset(output_chain_2_reset),
    .io_d(output_chain_2_io_d),
    .io_q(output_chain_2_io_q)
  );
  AsyncResetSynchronizerPrimitiveShiftReg_d3_i0 output_chain_3 ( // @[ShiftReg.scala 45:23]
    .clock(output_chain_3_clock),
    .reset(output_chain_3_reset),
    .io_d(output_chain_3_io_d),
    .io_q(output_chain_3_io_q)
  );
  assign io_q = {io_q_hi,io_q_lo}; // @[Cat.scala 33:92]
  assign output_chain_clock = clock;
  assign output_chain_reset = reset; // @[SynchronizerReg.scala 86:21]
  assign output_chain_io_d = io_d[0]; // @[SynchronizerReg.scala 87:41]
  assign output_chain_1_clock = clock;
  assign output_chain_1_reset = reset; // @[SynchronizerReg.scala 86:21]
  assign output_chain_1_io_d = io_d[1]; // @[SynchronizerReg.scala 87:41]
  assign output_chain_2_clock = clock;
  assign output_chain_2_reset = reset; // @[SynchronizerReg.scala 86:21]
  assign output_chain_2_io_d = io_d[2]; // @[SynchronizerReg.scala 87:41]
  assign output_chain_3_clock = clock;
  assign output_chain_3_reset = reset; // @[SynchronizerReg.scala 86:21]
  assign output_chain_3_io_d = io_d[3]; // @[SynchronizerReg.scala 87:41]
endmodule
module AsyncResetSynchronizerShiftReg_w1_d3_i0(
  input   clock,
  input   reset,
  input   io_d,
  output  io_q
);
  wire  output_chain_clock; // @[ShiftReg.scala 45:23]
  wire  output_chain_reset; // @[ShiftReg.scala 45:23]
  wire  output_chain_io_d; // @[ShiftReg.scala 45:23]
  wire  output_chain_io_q; // @[ShiftReg.scala 45:23]
  AsyncResetSynchronizerPrimitiveShiftReg_d3_i0 output_chain ( // @[ShiftReg.scala 45:23]
    .clock(output_chain_clock),
    .reset(output_chain_reset),
    .io_d(output_chain_io_d),
    .io_q(output_chain_io_q)
  );
  assign io_q = output_chain_io_q; // @[ShiftReg.scala 48:{24,24}]
  assign output_chain_clock = clock;
  assign output_chain_reset = reset; // @[SynchronizerReg.scala 86:21]
  assign output_chain_io_d = io_d; // @[SynchronizerReg.scala 87:41]
endmodule
module AsyncValidSync(
  input   io_in,
  output  io_out,
  input   clock,
  input   reset
);
  wire  io_out_source_valid_0_clock; // @[ShiftReg.scala 45:23]
  wire  io_out_source_valid_0_reset; // @[ShiftReg.scala 45:23]
  wire  io_out_source_valid_0_io_d; // @[ShiftReg.scala 45:23]
  wire  io_out_source_valid_0_io_q; // @[ShiftReg.scala 45:23]
  AsyncResetSynchronizerShiftReg_w1_d3_i0 io_out_source_valid_0 ( // @[ShiftReg.scala 45:23]
    .clock(io_out_source_valid_0_clock),
    .reset(io_out_source_valid_0_reset),
    .io_d(io_out_source_valid_0_io_d),
    .io_q(io_out_source_valid_0_io_q)
  );
  assign io_out = io_out_source_valid_0_io_q; // @[ShiftReg.scala 48:{24,24}]
  assign io_out_source_valid_0_clock = clock;
  assign io_out_source_valid_0_reset = reset;
  assign io_out_source_valid_0_io_d = io_in; // @[ShiftReg.scala 47:16]
endmodule
module AsyncQueueSource(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [7:0] io_enq_bits,
  output [7:0] io_async_mem_0,
  output [7:0] io_async_mem_1,
  output [7:0] io_async_mem_2,
  output [7:0] io_async_mem_3,
  output [7:0] io_async_mem_4,
  output [7:0] io_async_mem_5,
  output [7:0] io_async_mem_6,
  output [7:0] io_async_mem_7,
  input  [3:0] io_async_ridx,
  output [3:0] io_async_widx,
  input        io_async_safe_ridx_valid,
  output       io_async_safe_widx_valid,
  output       io_async_safe_source_reset_n,
  input        io_async_safe_sink_reset_n
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire  ridx_ridx_gray_clock; // @[ShiftReg.scala 45:23]
  wire  ridx_ridx_gray_reset; // @[ShiftReg.scala 45:23]
  wire [3:0] ridx_ridx_gray_io_d; // @[ShiftReg.scala 45:23]
  wire [3:0] ridx_ridx_gray_io_q; // @[ShiftReg.scala 45:23]
  wire  source_valid_0_io_in; // @[AsyncQueue.scala 100:32]
  wire  source_valid_0_io_out; // @[AsyncQueue.scala 100:32]
  wire  source_valid_0_clock; // @[AsyncQueue.scala 100:32]
  wire  source_valid_0_reset; // @[AsyncQueue.scala 100:32]
  wire  source_valid_1_io_in; // @[AsyncQueue.scala 101:32]
  wire  source_valid_1_io_out; // @[AsyncQueue.scala 101:32]
  wire  source_valid_1_clock; // @[AsyncQueue.scala 101:32]
  wire  source_valid_1_reset; // @[AsyncQueue.scala 101:32]
  wire  sink_extend_io_in; // @[AsyncQueue.scala 103:30]
  wire  sink_extend_io_out; // @[AsyncQueue.scala 103:30]
  wire  sink_extend_clock; // @[AsyncQueue.scala 103:30]
  wire  sink_extend_reset; // @[AsyncQueue.scala 103:30]
  wire  sink_valid_io_in; // @[AsyncQueue.scala 104:30]
  wire  sink_valid_io_out; // @[AsyncQueue.scala 104:30]
  wire  sink_valid_clock; // @[AsyncQueue.scala 104:30]
  wire  sink_valid_reset; // @[AsyncQueue.scala 104:30]
  reg [7:0] mem_0; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7; // @[AsyncQueue.scala 80:16]
  wire  _widx_T_1 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  sink_ready = sink_valid_io_out; // @[AsyncQueue.scala 120:16 79:28]
  wire  _widx_T_2 = ~sink_ready; // @[AsyncQueue.scala 81:79]
  reg [3:0] widx_widx_bin; // @[AsyncQueue.scala 52:25]
  wire [3:0] _GEN_16 = {{3'd0}, _widx_T_1}; // @[AsyncQueue.scala 53:43]
  wire [3:0] _widx_incremented_T_1 = widx_widx_bin + _GEN_16; // @[AsyncQueue.scala 53:43]
  wire [3:0] widx_incremented = _widx_T_2 ? 4'h0 : _widx_incremented_T_1; // @[AsyncQueue.scala 53:23]
  wire [3:0] _GEN_17 = {{1'd0}, widx_incremented[3:1]}; // @[AsyncQueue.scala 54:17]
  wire [3:0] widx = widx_incremented ^ _GEN_17; // @[AsyncQueue.scala 54:17]
  wire [3:0] ridx = ridx_ridx_gray_io_q; // @[ShiftReg.scala 48:{24,24}]
  wire [3:0] _ready_T = ridx ^ 4'hc; // @[AsyncQueue.scala 83:44]
  wire [2:0] _index_T_2 = {io_async_widx[3], 2'h0}; // @[AsyncQueue.scala 85:93]
  wire [2:0] index = io_async_widx[2:0] ^ _index_T_2; // @[AsyncQueue.scala 85:64]
  reg  ready_reg; // @[AsyncQueue.scala 88:56]
  reg [3:0] widx_gray; // @[AsyncQueue.scala 91:55]
  AsyncResetSynchronizerShiftReg_w4_d3_i0 ridx_ridx_gray ( // @[ShiftReg.scala 45:23]
    .clock(ridx_ridx_gray_clock),
    .reset(ridx_ridx_gray_reset),
    .io_d(ridx_ridx_gray_io_d),
    .io_q(ridx_ridx_gray_io_q)
  );
  AsyncValidSync source_valid_0 ( // @[AsyncQueue.scala 100:32]
    .io_in(source_valid_0_io_in),
    .io_out(source_valid_0_io_out),
    .clock(source_valid_0_clock),
    .reset(source_valid_0_reset)
  );
  AsyncValidSync source_valid_1 ( // @[AsyncQueue.scala 101:32]
    .io_in(source_valid_1_io_in),
    .io_out(source_valid_1_io_out),
    .clock(source_valid_1_clock),
    .reset(source_valid_1_reset)
  );
  AsyncValidSync sink_extend ( // @[AsyncQueue.scala 103:30]
    .io_in(sink_extend_io_in),
    .io_out(sink_extend_io_out),
    .clock(sink_extend_clock),
    .reset(sink_extend_reset)
  );
  AsyncValidSync sink_valid ( // @[AsyncQueue.scala 104:30]
    .io_in(sink_valid_io_in),
    .io_out(sink_valid_io_out),
    .clock(sink_valid_clock),
    .reset(sink_valid_reset)
  );
  assign io_enq_ready = ready_reg & sink_ready; // @[AsyncQueue.scala 89:29]
  assign io_async_mem_0 = mem_0; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1 = mem_1; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2 = mem_2; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3 = mem_3; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4 = mem_4; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5 = mem_5; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6 = mem_6; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7 = mem_7; // @[AsyncQueue.scala 96:31]
  assign io_async_widx = widx_gray; // @[AsyncQueue.scala 92:17]
  assign io_async_safe_widx_valid = source_valid_1_io_out; // @[AsyncQueue.scala 117:20]
  assign io_async_safe_source_reset_n = ~reset; // @[AsyncQueue.scala 121:27]
  assign ridx_ridx_gray_clock = clock;
  assign ridx_ridx_gray_reset = reset;
  assign ridx_ridx_gray_io_d = io_async_ridx; // @[ShiftReg.scala 47:16]
  assign source_valid_0_io_in = 1'h1; // @[AsyncQueue.scala 115:26]
  assign source_valid_0_clock = clock; // @[AsyncQueue.scala 110:26]
  assign source_valid_0_reset = reset | ~io_async_safe_sink_reset_n; // @[AsyncQueue.scala 105:65]
  assign source_valid_1_io_in = source_valid_0_io_out; // @[AsyncQueue.scala 116:26]
  assign source_valid_1_clock = clock; // @[AsyncQueue.scala 111:26]
  assign source_valid_1_reset = reset | ~io_async_safe_sink_reset_n; // @[AsyncQueue.scala 106:65]
  assign sink_extend_io_in = io_async_safe_ridx_valid; // @[AsyncQueue.scala 118:23]
  assign sink_extend_clock = clock; // @[AsyncQueue.scala 112:26]
  assign sink_extend_reset = reset | ~io_async_safe_sink_reset_n; // @[AsyncQueue.scala 107:65]
  assign sink_valid_io_in = sink_extend_io_out; // @[AsyncQueue.scala 119:22]
  assign sink_valid_clock = clock; // @[AsyncQueue.scala 113:26]
  assign sink_valid_reset = reset; // @[AsyncQueue.scala 108:35]
  always @(posedge clock) begin
    if (_widx_T_1) begin // @[AsyncQueue.scala 86:24]
      if (3'h0 == index) begin // @[AsyncQueue.scala 86:37]
        mem_0 <= io_enq_bits; // @[AsyncQueue.scala 86:37]
      end
    end
    if (_widx_T_1) begin // @[AsyncQueue.scala 86:24]
      if (3'h1 == index) begin // @[AsyncQueue.scala 86:37]
        mem_1 <= io_enq_bits; // @[AsyncQueue.scala 86:37]
      end
    end
    if (_widx_T_1) begin // @[AsyncQueue.scala 86:24]
      if (3'h2 == index) begin // @[AsyncQueue.scala 86:37]
        mem_2 <= io_enq_bits; // @[AsyncQueue.scala 86:37]
      end
    end
    if (_widx_T_1) begin // @[AsyncQueue.scala 86:24]
      if (3'h3 == index) begin // @[AsyncQueue.scala 86:37]
        mem_3 <= io_enq_bits; // @[AsyncQueue.scala 86:37]
      end
    end
    if (_widx_T_1) begin // @[AsyncQueue.scala 86:24]
      if (3'h4 == index) begin // @[AsyncQueue.scala 86:37]
        mem_4 <= io_enq_bits; // @[AsyncQueue.scala 86:37]
      end
    end
    if (_widx_T_1) begin // @[AsyncQueue.scala 86:24]
      if (3'h5 == index) begin // @[AsyncQueue.scala 86:37]
        mem_5 <= io_enq_bits; // @[AsyncQueue.scala 86:37]
      end
    end
    if (_widx_T_1) begin // @[AsyncQueue.scala 86:24]
      if (3'h6 == index) begin // @[AsyncQueue.scala 86:37]
        mem_6 <= io_enq_bits; // @[AsyncQueue.scala 86:37]
      end
    end
    if (_widx_T_1) begin // @[AsyncQueue.scala 86:24]
      if (3'h7 == index) begin // @[AsyncQueue.scala 86:37]
        mem_7 <= io_enq_bits; // @[AsyncQueue.scala 86:37]
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsyncQueue.scala 53:23]
      widx_widx_bin <= 4'h0;
    end else if (_widx_T_2) begin
      widx_widx_bin <= 4'h0;
    end else begin
      widx_widx_bin <= _widx_incremented_T_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsyncQueue.scala 83:26]
      ready_reg <= 1'h0;
    end else begin
      ready_reg <= sink_ready & widx != _ready_T;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsyncQueue.scala 54:17]
      widx_gray <= 4'h0;
    end else begin
      widx_gray <= widx_incremented ^ _GEN_17;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mem_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  mem_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  mem_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  mem_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  mem_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  mem_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  mem_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  mem_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  widx_widx_bin = _RAND_8[3:0];
  _RAND_9 = {1{`RANDOM}};
  ready_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  widx_gray = _RAND_10[3:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    widx_widx_bin = 4'h0;
  end
  if (reset) begin
    ready_reg = 1'h0;
  end
  if (reset) begin
    widx_gray = 4'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ClockCrossingReg_w8(
  input        clock,
  input  [7:0] io_d,
  output [7:0] io_q,
  input        io_en
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] cdc_reg; // @[Reg.scala 19:16]
  assign io_q = cdc_reg; // @[SynchronizerReg.scala 202:8]
  always @(posedge clock) begin
    if (io_en) begin // @[Reg.scala 20:18]
      cdc_reg <= io_d; // @[Reg.scala 20:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cdc_reg = _RAND_0[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AsyncQueueSink(
  input        clock,
  input        reset,
  input        io_deq_ready,
  output       io_deq_valid,
  output [7:0] io_deq_bits,
  input  [7:0] io_async_mem_0,
  input  [7:0] io_async_mem_1,
  input  [7:0] io_async_mem_2,
  input  [7:0] io_async_mem_3,
  input  [7:0] io_async_mem_4,
  input  [7:0] io_async_mem_5,
  input  [7:0] io_async_mem_6,
  input  [7:0] io_async_mem_7,
  output [3:0] io_async_ridx,
  input  [3:0] io_async_widx,
  output       io_async_safe_ridx_valid,
  input        io_async_safe_widx_valid,
  input        io_async_safe_source_reset_n,
  output       io_async_safe_sink_reset_n
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  widx_widx_gray_clock; // @[ShiftReg.scala 45:23]
  wire  widx_widx_gray_reset; // @[ShiftReg.scala 45:23]
  wire [3:0] widx_widx_gray_io_d; // @[ShiftReg.scala 45:23]
  wire [3:0] widx_widx_gray_io_q; // @[ShiftReg.scala 45:23]
  wire  io_deq_bits_deq_bits_reg_clock; // @[SynchronizerReg.scala 207:25]
  wire [7:0] io_deq_bits_deq_bits_reg_io_d; // @[SynchronizerReg.scala 207:25]
  wire [7:0] io_deq_bits_deq_bits_reg_io_q; // @[SynchronizerReg.scala 207:25]
  wire  io_deq_bits_deq_bits_reg_io_en; // @[SynchronizerReg.scala 207:25]
  wire  sink_valid_0_io_in; // @[AsyncQueue.scala 168:33]
  wire  sink_valid_0_io_out; // @[AsyncQueue.scala 168:33]
  wire  sink_valid_0_clock; // @[AsyncQueue.scala 168:33]
  wire  sink_valid_0_reset; // @[AsyncQueue.scala 168:33]
  wire  sink_valid_1_io_in; // @[AsyncQueue.scala 169:33]
  wire  sink_valid_1_io_out; // @[AsyncQueue.scala 169:33]
  wire  sink_valid_1_clock; // @[AsyncQueue.scala 169:33]
  wire  sink_valid_1_reset; // @[AsyncQueue.scala 169:33]
  wire  source_extend_io_in; // @[AsyncQueue.scala 171:31]
  wire  source_extend_io_out; // @[AsyncQueue.scala 171:31]
  wire  source_extend_clock; // @[AsyncQueue.scala 171:31]
  wire  source_extend_reset; // @[AsyncQueue.scala 171:31]
  wire  source_valid_io_in; // @[AsyncQueue.scala 172:31]
  wire  source_valid_io_out; // @[AsyncQueue.scala 172:31]
  wire  source_valid_clock; // @[AsyncQueue.scala 172:31]
  wire  source_valid_reset; // @[AsyncQueue.scala 172:31]
  wire  _ridx_T_1 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  wire  source_ready = source_valid_io_out; // @[AsyncQueue.scala 143:30 188:18]
  wire  _ridx_T_2 = ~source_ready; // @[AsyncQueue.scala 144:79]
  reg [3:0] ridx_ridx_bin; // @[AsyncQueue.scala 52:25]
  wire [3:0] _GEN_8 = {{3'd0}, _ridx_T_1}; // @[AsyncQueue.scala 53:43]
  wire [3:0] _ridx_incremented_T_1 = ridx_ridx_bin + _GEN_8; // @[AsyncQueue.scala 53:43]
  wire [3:0] ridx_incremented = _ridx_T_2 ? 4'h0 : _ridx_incremented_T_1; // @[AsyncQueue.scala 53:23]
  wire [3:0] _GEN_9 = {{1'd0}, ridx_incremented[3:1]}; // @[AsyncQueue.scala 54:17]
  wire [3:0] ridx = ridx_incremented ^ _GEN_9; // @[AsyncQueue.scala 54:17]
  wire [3:0] widx = widx_widx_gray_io_q; // @[ShiftReg.scala 48:{24,24}]
  wire [2:0] _index_T_2 = {ridx[3], 2'h0}; // @[AsyncQueue.scala 152:75]
  wire [2:0] index = ridx[2:0] ^ _index_T_2; // @[AsyncQueue.scala 152:55]
  wire [7:0] _GEN_1 = 3'h1 == index ? io_async_mem_1 : io_async_mem_0; // @[SynchronizerReg.scala 209:{18,18}]
  wire [7:0] _GEN_2 = 3'h2 == index ? io_async_mem_2 : _GEN_1; // @[SynchronizerReg.scala 209:{18,18}]
  wire [7:0] _GEN_3 = 3'h3 == index ? io_async_mem_3 : _GEN_2; // @[SynchronizerReg.scala 209:{18,18}]
  wire [7:0] _GEN_4 = 3'h4 == index ? io_async_mem_4 : _GEN_3; // @[SynchronizerReg.scala 209:{18,18}]
  wire [7:0] _GEN_5 = 3'h5 == index ? io_async_mem_5 : _GEN_4; // @[SynchronizerReg.scala 209:{18,18}]
  wire [7:0] _GEN_6 = 3'h6 == index ? io_async_mem_6 : _GEN_5; // @[SynchronizerReg.scala 209:{18,18}]
  reg  valid_reg; // @[AsyncQueue.scala 161:56]
  reg [3:0] ridx_gray; // @[AsyncQueue.scala 164:55]
  AsyncResetSynchronizerShiftReg_w4_d3_i0 widx_widx_gray ( // @[ShiftReg.scala 45:23]
    .clock(widx_widx_gray_clock),
    .reset(widx_widx_gray_reset),
    .io_d(widx_widx_gray_io_d),
    .io_q(widx_widx_gray_io_q)
  );
  ClockCrossingReg_w8 io_deq_bits_deq_bits_reg ( // @[SynchronizerReg.scala 207:25]
    .clock(io_deq_bits_deq_bits_reg_clock),
    .io_d(io_deq_bits_deq_bits_reg_io_d),
    .io_q(io_deq_bits_deq_bits_reg_io_q),
    .io_en(io_deq_bits_deq_bits_reg_io_en)
  );
  AsyncValidSync sink_valid_0 ( // @[AsyncQueue.scala 168:33]
    .io_in(sink_valid_0_io_in),
    .io_out(sink_valid_0_io_out),
    .clock(sink_valid_0_clock),
    .reset(sink_valid_0_reset)
  );
  AsyncValidSync sink_valid_1 ( // @[AsyncQueue.scala 169:33]
    .io_in(sink_valid_1_io_in),
    .io_out(sink_valid_1_io_out),
    .clock(sink_valid_1_clock),
    .reset(sink_valid_1_reset)
  );
  AsyncValidSync source_extend ( // @[AsyncQueue.scala 171:31]
    .io_in(source_extend_io_in),
    .io_out(source_extend_io_out),
    .clock(source_extend_clock),
    .reset(source_extend_reset)
  );
  AsyncValidSync source_valid ( // @[AsyncQueue.scala 172:31]
    .io_in(source_valid_io_in),
    .io_out(source_valid_io_out),
    .clock(source_valid_clock),
    .reset(source_valid_reset)
  );
  assign io_deq_valid = valid_reg & source_ready; // @[AsyncQueue.scala 162:29]
  assign io_deq_bits = io_deq_bits_deq_bits_reg_io_q; // @[SynchronizerReg.scala 211:{26,26}]
  assign io_async_ridx = ridx_gray; // @[AsyncQueue.scala 165:17]
  assign io_async_safe_ridx_valid = sink_valid_1_io_out; // @[AsyncQueue.scala 185:20]
  assign io_async_safe_sink_reset_n = ~reset; // @[AsyncQueue.scala 189:25]
  assign widx_widx_gray_clock = clock;
  assign widx_widx_gray_reset = reset;
  assign widx_widx_gray_io_d = io_async_widx; // @[ShiftReg.scala 47:16]
  assign io_deq_bits_deq_bits_reg_clock = clock;
  assign io_deq_bits_deq_bits_reg_io_d = 3'h7 == index ? io_async_mem_7 : _GEN_6; // @[SynchronizerReg.scala 209:{18,18}]
  assign io_deq_bits_deq_bits_reg_io_en = source_ready & ridx != widx; // @[AsyncQueue.scala 146:28]
  assign sink_valid_0_io_in = 1'h1; // @[AsyncQueue.scala 183:24]
  assign sink_valid_0_clock = clock; // @[AsyncQueue.scala 178:25]
  assign sink_valid_0_reset = reset | ~io_async_safe_source_reset_n; // @[AsyncQueue.scala 173:66]
  assign sink_valid_1_io_in = sink_valid_0_io_out; // @[AsyncQueue.scala 184:24]
  assign sink_valid_1_clock = clock; // @[AsyncQueue.scala 179:25]
  assign sink_valid_1_reset = reset | ~io_async_safe_source_reset_n; // @[AsyncQueue.scala 174:66]
  assign source_extend_io_in = io_async_safe_widx_valid; // @[AsyncQueue.scala 186:25]
  assign source_extend_clock = clock; // @[AsyncQueue.scala 180:25]
  assign source_extend_reset = reset | ~io_async_safe_source_reset_n; // @[AsyncQueue.scala 175:66]
  assign source_valid_io_in = source_extend_io_out; // @[AsyncQueue.scala 187:24]
  assign source_valid_clock = clock; // @[AsyncQueue.scala 181:25]
  assign source_valid_reset = reset; // @[AsyncQueue.scala 176:34]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsyncQueue.scala 53:23]
      ridx_ridx_bin <= 4'h0;
    end else if (_ridx_T_2) begin
      ridx_ridx_bin <= 4'h0;
    end else begin
      ridx_ridx_bin <= _ridx_incremented_T_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsyncQueue.scala 146:28]
      valid_reg <= 1'h0;
    end else begin
      valid_reg <= source_ready & ridx != widx;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsyncQueue.scala 54:17]
      ridx_gray <= 4'h0;
    end else begin
      ridx_gray <= ridx_incremented ^ _GEN_9;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ridx_ridx_bin = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  ridx_gray = _RAND_2[3:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    ridx_ridx_bin = 4'h0;
  end
  if (reset) begin
    valid_reg = 1'h0;
  end
  if (reset) begin
    ridx_gray = 4'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AsyncQueue(
  input        io_enq_clock,
  input        io_enq_reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [7:0] io_enq_bits,
  input        io_deq_clock,
  input        io_deq_reset,
  input        io_deq_ready,
  output       io_deq_valid,
  output [7:0] io_deq_bits
);
  wire  source_clock; // @[AsyncQueue.scala 224:22]
  wire  source_reset; // @[AsyncQueue.scala 224:22]
  wire  source_io_enq_ready; // @[AsyncQueue.scala 224:22]
  wire  source_io_enq_valid; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7; // @[AsyncQueue.scala 224:22]
  wire [3:0] source_io_async_ridx; // @[AsyncQueue.scala 224:22]
  wire [3:0] source_io_async_widx; // @[AsyncQueue.scala 224:22]
  wire  source_io_async_safe_ridx_valid; // @[AsyncQueue.scala 224:22]
  wire  source_io_async_safe_widx_valid; // @[AsyncQueue.scala 224:22]
  wire  source_io_async_safe_source_reset_n; // @[AsyncQueue.scala 224:22]
  wire  source_io_async_safe_sink_reset_n; // @[AsyncQueue.scala 224:22]
  wire  sink_clock; // @[AsyncQueue.scala 225:22]
  wire  sink_reset; // @[AsyncQueue.scala 225:22]
  wire  sink_io_deq_ready; // @[AsyncQueue.scala 225:22]
  wire  sink_io_deq_valid; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7; // @[AsyncQueue.scala 225:22]
  wire [3:0] sink_io_async_ridx; // @[AsyncQueue.scala 225:22]
  wire [3:0] sink_io_async_widx; // @[AsyncQueue.scala 225:22]
  wire  sink_io_async_safe_ridx_valid; // @[AsyncQueue.scala 225:22]
  wire  sink_io_async_safe_widx_valid; // @[AsyncQueue.scala 225:22]
  wire  sink_io_async_safe_source_reset_n; // @[AsyncQueue.scala 225:22]
  wire  sink_io_async_safe_sink_reset_n; // @[AsyncQueue.scala 225:22]
  AsyncQueueSource source ( // @[AsyncQueue.scala 224:22]
    .clock(source_clock),
    .reset(source_reset),
    .io_enq_ready(source_io_enq_ready),
    .io_enq_valid(source_io_enq_valid),
    .io_enq_bits(source_io_enq_bits),
    .io_async_mem_0(source_io_async_mem_0),
    .io_async_mem_1(source_io_async_mem_1),
    .io_async_mem_2(source_io_async_mem_2),
    .io_async_mem_3(source_io_async_mem_3),
    .io_async_mem_4(source_io_async_mem_4),
    .io_async_mem_5(source_io_async_mem_5),
    .io_async_mem_6(source_io_async_mem_6),
    .io_async_mem_7(source_io_async_mem_7),
    .io_async_ridx(source_io_async_ridx),
    .io_async_widx(source_io_async_widx),
    .io_async_safe_ridx_valid(source_io_async_safe_ridx_valid),
    .io_async_safe_widx_valid(source_io_async_safe_widx_valid),
    .io_async_safe_source_reset_n(source_io_async_safe_source_reset_n),
    .io_async_safe_sink_reset_n(source_io_async_safe_sink_reset_n)
  );
  AsyncQueueSink sink ( // @[AsyncQueue.scala 225:22]
    .clock(sink_clock),
    .reset(sink_reset),
    .io_deq_ready(sink_io_deq_ready),
    .io_deq_valid(sink_io_deq_valid),
    .io_deq_bits(sink_io_deq_bits),
    .io_async_mem_0(sink_io_async_mem_0),
    .io_async_mem_1(sink_io_async_mem_1),
    .io_async_mem_2(sink_io_async_mem_2),
    .io_async_mem_3(sink_io_async_mem_3),
    .io_async_mem_4(sink_io_async_mem_4),
    .io_async_mem_5(sink_io_async_mem_5),
    .io_async_mem_6(sink_io_async_mem_6),
    .io_async_mem_7(sink_io_async_mem_7),
    .io_async_ridx(sink_io_async_ridx),
    .io_async_widx(sink_io_async_widx),
    .io_async_safe_ridx_valid(sink_io_async_safe_ridx_valid),
    .io_async_safe_widx_valid(sink_io_async_safe_widx_valid),
    .io_async_safe_source_reset_n(sink_io_async_safe_source_reset_n),
    .io_async_safe_sink_reset_n(sink_io_async_safe_sink_reset_n)
  );
  assign io_enq_ready = source_io_enq_ready; // @[AsyncQueue.scala 232:17]
  assign io_deq_valid = sink_io_deq_valid; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits = sink_io_deq_bits; // @[AsyncQueue.scala 233:10]
  assign source_clock = io_enq_clock; // @[AsyncQueue.scala 227:16]
  assign source_reset = io_enq_reset; // @[AsyncQueue.scala 228:16]
  assign source_io_enq_valid = io_enq_valid; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits = io_enq_bits; // @[AsyncQueue.scala 232:17]
  assign source_io_async_ridx = sink_io_async_ridx; // @[AsyncQueue.scala 234:17]
  assign source_io_async_safe_ridx_valid = sink_io_async_safe_ridx_valid; // @[AsyncQueue.scala 234:17]
  assign source_io_async_safe_sink_reset_n = sink_io_async_safe_sink_reset_n; // @[AsyncQueue.scala 234:17]
  assign sink_clock = io_deq_clock; // @[AsyncQueue.scala 229:14]
  assign sink_reset = io_deq_reset; // @[AsyncQueue.scala 230:14]
  assign sink_io_deq_ready = io_deq_ready; // @[AsyncQueue.scala 233:10]
  assign sink_io_async_mem_0 = source_io_async_mem_0; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1 = source_io_async_mem_1; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2 = source_io_async_mem_2; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3 = source_io_async_mem_3; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4 = source_io_async_mem_4; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5 = source_io_async_mem_5; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6 = source_io_async_mem_6; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7 = source_io_async_mem_7; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_widx = source_io_async_widx; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_safe_widx_valid = source_io_async_safe_widx_valid; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_safe_source_reset_n = source_io_async_safe_source_reset_n; // @[AsyncQueue.scala 234:17]
endmodule
module SoC(
  input        clock,
  input        reset,
  output       io_in_ready,
  input        io_in_valid,
  input  [7:0] io_in_bits,
  input        io_out_ready,
  output       io_out_valid,
  output [7:0] io_out_bits,
  input        io_io_clock,
  input        io_io_reset,
  input        io_intr_mtip,
  input        io_intr_msip,
  input        io_intr_meip,
  input        io_intr_seip
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  wire  soc_imp_clock; // @[SoC.scala 81:27]
  wire  soc_imp_reset; // @[SoC.scala 81:27]
  wire  soc_imp_auto_out_a_ready; // @[SoC.scala 81:27]
  wire  soc_imp_auto_out_a_valid; // @[SoC.scala 81:27]
  wire [2:0] soc_imp_auto_out_a_bits_opcode; // @[SoC.scala 81:27]
  wire [2:0] soc_imp_auto_out_a_bits_param; // @[SoC.scala 81:27]
  wire [2:0] soc_imp_auto_out_a_bits_size; // @[SoC.scala 81:27]
  wire [3:0] soc_imp_auto_out_a_bits_source; // @[SoC.scala 81:27]
  wire [31:0] soc_imp_auto_out_a_bits_address; // @[SoC.scala 81:27]
  wire [31:0] soc_imp_auto_out_a_bits_mask; // @[SoC.scala 81:27]
  wire [255:0] soc_imp_auto_out_a_bits_data; // @[SoC.scala 81:27]
  wire  soc_imp_auto_out_b_ready; // @[SoC.scala 81:27]
  wire  soc_imp_auto_out_b_valid; // @[SoC.scala 81:27]
  wire [2:0] soc_imp_auto_out_b_bits_size; // @[SoC.scala 81:27]
  wire [3:0] soc_imp_auto_out_b_bits_source; // @[SoC.scala 81:27]
  wire [31:0] soc_imp_auto_out_b_bits_address; // @[SoC.scala 81:27]
  wire  soc_imp_auto_out_c_ready; // @[SoC.scala 81:27]
  wire  soc_imp_auto_out_c_valid; // @[SoC.scala 81:27]
  wire [2:0] soc_imp_auto_out_c_bits_opcode; // @[SoC.scala 81:27]
  wire [2:0] soc_imp_auto_out_c_bits_param; // @[SoC.scala 81:27]
  wire [2:0] soc_imp_auto_out_c_bits_size; // @[SoC.scala 81:27]
  wire [3:0] soc_imp_auto_out_c_bits_source; // @[SoC.scala 81:27]
  wire [31:0] soc_imp_auto_out_c_bits_address; // @[SoC.scala 81:27]
  wire [255:0] soc_imp_auto_out_c_bits_data; // @[SoC.scala 81:27]
  wire  soc_imp_auto_out_d_ready; // @[SoC.scala 81:27]
  wire  soc_imp_auto_out_d_valid; // @[SoC.scala 81:27]
  wire [2:0] soc_imp_auto_out_d_bits_opcode; // @[SoC.scala 81:27]
  wire [2:0] soc_imp_auto_out_d_bits_size; // @[SoC.scala 81:27]
  wire [3:0] soc_imp_auto_out_d_bits_source; // @[SoC.scala 81:27]
  wire [5:0] soc_imp_auto_out_d_bits_sink; // @[SoC.scala 81:27]
  wire [255:0] soc_imp_auto_out_d_bits_data; // @[SoC.scala 81:27]
  wire  soc_imp_auto_out_e_ready; // @[SoC.scala 81:27]
  wire  soc_imp_auto_out_e_valid; // @[SoC.scala 81:27]
  wire [5:0] soc_imp_auto_out_e_bits_sink; // @[SoC.scala 81:27]
  wire  soc_imp_io_intr_mtip; // @[SoC.scala 81:27]
  wire  soc_imp_io_intr_msip; // @[SoC.scala 81:27]
  wire  soc_imp_io_intr_meip; // @[SoC.scala 81:27]
  wire  soc_imp_io_intr_seip; // @[SoC.scala 81:27]
  wire  serdes_clock; // @[SoC.scala 87:26]
  wire  serdes_reset; // @[SoC.scala 87:26]
  wire  serdes_auto_in_a_ready; // @[SoC.scala 87:26]
  wire  serdes_auto_in_a_valid; // @[SoC.scala 87:26]
  wire [2:0] serdes_auto_in_a_bits_opcode; // @[SoC.scala 87:26]
  wire [2:0] serdes_auto_in_a_bits_param; // @[SoC.scala 87:26]
  wire [2:0] serdes_auto_in_a_bits_size; // @[SoC.scala 87:26]
  wire [3:0] serdes_auto_in_a_bits_source; // @[SoC.scala 87:26]
  wire [31:0] serdes_auto_in_a_bits_address; // @[SoC.scala 87:26]
  wire [31:0] serdes_auto_in_a_bits_mask; // @[SoC.scala 87:26]
  wire [255:0] serdes_auto_in_a_bits_data; // @[SoC.scala 87:26]
  wire  serdes_auto_in_b_ready; // @[SoC.scala 87:26]
  wire  serdes_auto_in_b_valid; // @[SoC.scala 87:26]
  wire [2:0] serdes_auto_in_b_bits_size; // @[SoC.scala 87:26]
  wire [3:0] serdes_auto_in_b_bits_source; // @[SoC.scala 87:26]
  wire [31:0] serdes_auto_in_b_bits_address; // @[SoC.scala 87:26]
  wire  serdes_auto_in_c_ready; // @[SoC.scala 87:26]
  wire  serdes_auto_in_c_valid; // @[SoC.scala 87:26]
  wire [2:0] serdes_auto_in_c_bits_opcode; // @[SoC.scala 87:26]
  wire [2:0] serdes_auto_in_c_bits_param; // @[SoC.scala 87:26]
  wire [2:0] serdes_auto_in_c_bits_size; // @[SoC.scala 87:26]
  wire [3:0] serdes_auto_in_c_bits_source; // @[SoC.scala 87:26]
  wire [31:0] serdes_auto_in_c_bits_address; // @[SoC.scala 87:26]
  wire [255:0] serdes_auto_in_c_bits_data; // @[SoC.scala 87:26]
  wire  serdes_auto_in_d_ready; // @[SoC.scala 87:26]
  wire  serdes_auto_in_d_valid; // @[SoC.scala 87:26]
  wire [2:0] serdes_auto_in_d_bits_opcode; // @[SoC.scala 87:26]
  wire [2:0] serdes_auto_in_d_bits_size; // @[SoC.scala 87:26]
  wire [3:0] serdes_auto_in_d_bits_source; // @[SoC.scala 87:26]
  wire [5:0] serdes_auto_in_d_bits_sink; // @[SoC.scala 87:26]
  wire [255:0] serdes_auto_in_d_bits_data; // @[SoC.scala 87:26]
  wire  serdes_auto_in_e_ready; // @[SoC.scala 87:26]
  wire  serdes_auto_in_e_valid; // @[SoC.scala 87:26]
  wire [5:0] serdes_auto_in_e_bits_sink; // @[SoC.scala 87:26]
  wire  serdes_io_ser_0_in_ready; // @[SoC.scala 87:26]
  wire  serdes_io_ser_0_in_valid; // @[SoC.scala 87:26]
  wire [7:0] serdes_io_ser_0_in_bits; // @[SoC.scala 87:26]
  wire  serdes_io_ser_0_out_ready; // @[SoC.scala 87:26]
  wire  serdes_io_ser_0_out_valid; // @[SoC.scala 87:26]
  wire [7:0] serdes_io_ser_0_out_bits; // @[SoC.scala 87:26]
  wire  trace_buffer_clock; // @[TLTraceBuffer.scala 47:34]
  wire  trace_buffer_reset; // @[TLTraceBuffer.scala 47:34]
  wire  trace_buffer_auto_in_a_ready; // @[TLTraceBuffer.scala 47:34]
  wire  trace_buffer_auto_in_a_valid; // @[TLTraceBuffer.scala 47:34]
  wire [2:0] trace_buffer_auto_in_a_bits_opcode; // @[TLTraceBuffer.scala 47:34]
  wire [2:0] trace_buffer_auto_in_a_bits_param; // @[TLTraceBuffer.scala 47:34]
  wire [2:0] trace_buffer_auto_in_a_bits_size; // @[TLTraceBuffer.scala 47:34]
  wire [3:0] trace_buffer_auto_in_a_bits_source; // @[TLTraceBuffer.scala 47:34]
  wire [31:0] trace_buffer_auto_in_a_bits_address; // @[TLTraceBuffer.scala 47:34]
  wire [31:0] trace_buffer_auto_in_a_bits_mask; // @[TLTraceBuffer.scala 47:34]
  wire [255:0] trace_buffer_auto_in_a_bits_data; // @[TLTraceBuffer.scala 47:34]
  wire  trace_buffer_auto_in_b_ready; // @[TLTraceBuffer.scala 47:34]
  wire  trace_buffer_auto_in_b_valid; // @[TLTraceBuffer.scala 47:34]
  wire [2:0] trace_buffer_auto_in_b_bits_size; // @[TLTraceBuffer.scala 47:34]
  wire [3:0] trace_buffer_auto_in_b_bits_source; // @[TLTraceBuffer.scala 47:34]
  wire [31:0] trace_buffer_auto_in_b_bits_address; // @[TLTraceBuffer.scala 47:34]
  wire  trace_buffer_auto_in_c_ready; // @[TLTraceBuffer.scala 47:34]
  wire  trace_buffer_auto_in_c_valid; // @[TLTraceBuffer.scala 47:34]
  wire [2:0] trace_buffer_auto_in_c_bits_opcode; // @[TLTraceBuffer.scala 47:34]
  wire [2:0] trace_buffer_auto_in_c_bits_param; // @[TLTraceBuffer.scala 47:34]
  wire [2:0] trace_buffer_auto_in_c_bits_size; // @[TLTraceBuffer.scala 47:34]
  wire [3:0] trace_buffer_auto_in_c_bits_source; // @[TLTraceBuffer.scala 47:34]
  wire [31:0] trace_buffer_auto_in_c_bits_address; // @[TLTraceBuffer.scala 47:34]
  wire [255:0] trace_buffer_auto_in_c_bits_data; // @[TLTraceBuffer.scala 47:34]
  wire  trace_buffer_auto_in_d_ready; // @[TLTraceBuffer.scala 47:34]
  wire  trace_buffer_auto_in_d_valid; // @[TLTraceBuffer.scala 47:34]
  wire [2:0] trace_buffer_auto_in_d_bits_opcode; // @[TLTraceBuffer.scala 47:34]
  wire [2:0] trace_buffer_auto_in_d_bits_size; // @[TLTraceBuffer.scala 47:34]
  wire [3:0] trace_buffer_auto_in_d_bits_source; // @[TLTraceBuffer.scala 47:34]
  wire [5:0] trace_buffer_auto_in_d_bits_sink; // @[TLTraceBuffer.scala 47:34]
  wire [255:0] trace_buffer_auto_in_d_bits_data; // @[TLTraceBuffer.scala 47:34]
  wire  trace_buffer_auto_in_e_ready; // @[TLTraceBuffer.scala 47:34]
  wire  trace_buffer_auto_in_e_valid; // @[TLTraceBuffer.scala 47:34]
  wire [5:0] trace_buffer_auto_in_e_bits_sink; // @[TLTraceBuffer.scala 47:34]
  wire  trace_buffer_auto_out_a_ready; // @[TLTraceBuffer.scala 47:34]
  wire  trace_buffer_auto_out_a_valid; // @[TLTraceBuffer.scala 47:34]
  wire [2:0] trace_buffer_auto_out_a_bits_opcode; // @[TLTraceBuffer.scala 47:34]
  wire [2:0] trace_buffer_auto_out_a_bits_param; // @[TLTraceBuffer.scala 47:34]
  wire [2:0] trace_buffer_auto_out_a_bits_size; // @[TLTraceBuffer.scala 47:34]
  wire [3:0] trace_buffer_auto_out_a_bits_source; // @[TLTraceBuffer.scala 47:34]
  wire [31:0] trace_buffer_auto_out_a_bits_address; // @[TLTraceBuffer.scala 47:34]
  wire [31:0] trace_buffer_auto_out_a_bits_mask; // @[TLTraceBuffer.scala 47:34]
  wire [255:0] trace_buffer_auto_out_a_bits_data; // @[TLTraceBuffer.scala 47:34]
  wire  trace_buffer_auto_out_b_ready; // @[TLTraceBuffer.scala 47:34]
  wire  trace_buffer_auto_out_b_valid; // @[TLTraceBuffer.scala 47:34]
  wire [2:0] trace_buffer_auto_out_b_bits_size; // @[TLTraceBuffer.scala 47:34]
  wire [3:0] trace_buffer_auto_out_b_bits_source; // @[TLTraceBuffer.scala 47:34]
  wire [31:0] trace_buffer_auto_out_b_bits_address; // @[TLTraceBuffer.scala 47:34]
  wire  trace_buffer_auto_out_c_ready; // @[TLTraceBuffer.scala 47:34]
  wire  trace_buffer_auto_out_c_valid; // @[TLTraceBuffer.scala 47:34]
  wire [2:0] trace_buffer_auto_out_c_bits_opcode; // @[TLTraceBuffer.scala 47:34]
  wire [2:0] trace_buffer_auto_out_c_bits_param; // @[TLTraceBuffer.scala 47:34]
  wire [2:0] trace_buffer_auto_out_c_bits_size; // @[TLTraceBuffer.scala 47:34]
  wire [3:0] trace_buffer_auto_out_c_bits_source; // @[TLTraceBuffer.scala 47:34]
  wire [31:0] trace_buffer_auto_out_c_bits_address; // @[TLTraceBuffer.scala 47:34]
  wire [255:0] trace_buffer_auto_out_c_bits_data; // @[TLTraceBuffer.scala 47:34]
  wire  trace_buffer_auto_out_d_ready; // @[TLTraceBuffer.scala 47:34]
  wire  trace_buffer_auto_out_d_valid; // @[TLTraceBuffer.scala 47:34]
  wire [2:0] trace_buffer_auto_out_d_bits_opcode; // @[TLTraceBuffer.scala 47:34]
  wire [2:0] trace_buffer_auto_out_d_bits_size; // @[TLTraceBuffer.scala 47:34]
  wire [3:0] trace_buffer_auto_out_d_bits_source; // @[TLTraceBuffer.scala 47:34]
  wire [5:0] trace_buffer_auto_out_d_bits_sink; // @[TLTraceBuffer.scala 47:34]
  wire [255:0] trace_buffer_auto_out_d_bits_data; // @[TLTraceBuffer.scala 47:34]
  wire  trace_buffer_auto_out_e_ready; // @[TLTraceBuffer.scala 47:34]
  wire  trace_buffer_auto_out_e_valid; // @[TLTraceBuffer.scala 47:34]
  wire [5:0] trace_buffer_auto_out_e_bits_sink; // @[TLTraceBuffer.scala 47:34]
  wire  in_fifo_io_enq_clock; // @[SoC.scala 111:26]
  wire  in_fifo_io_enq_reset; // @[SoC.scala 111:26]
  wire  in_fifo_io_enq_ready; // @[SoC.scala 111:26]
  wire  in_fifo_io_enq_valid; // @[SoC.scala 111:26]
  wire [7:0] in_fifo_io_enq_bits; // @[SoC.scala 111:26]
  wire  in_fifo_io_deq_clock; // @[SoC.scala 111:26]
  wire  in_fifo_io_deq_reset; // @[SoC.scala 111:26]
  wire  in_fifo_io_deq_ready; // @[SoC.scala 111:26]
  wire  in_fifo_io_deq_valid; // @[SoC.scala 111:26]
  wire [7:0] in_fifo_io_deq_bits; // @[SoC.scala 111:26]
  wire  out_fifo_io_enq_clock; // @[SoC.scala 112:26]
  wire  out_fifo_io_enq_reset; // @[SoC.scala 112:26]
  wire  out_fifo_io_enq_ready; // @[SoC.scala 112:26]
  wire  out_fifo_io_enq_valid; // @[SoC.scala 112:26]
  wire [7:0] out_fifo_io_enq_bits; // @[SoC.scala 112:26]
  wire  out_fifo_io_deq_clock; // @[SoC.scala 112:26]
  wire  out_fifo_io_deq_reset; // @[SoC.scala 112:26]
  wire  out_fifo_io_deq_ready; // @[SoC.scala 112:26]
  wire  out_fifo_io_deq_valid; // @[SoC.scala 112:26]
  wire [7:0] out_fifo_io_deq_bits; // @[SoC.scala 112:26]
  reg  sync_dff_0_mtip; // @[SoC.scala 127:27]
  reg  sync_dff_0_msip; // @[SoC.scala 127:27]
  reg  sync_dff_0_meip; // @[SoC.scala 127:27]
  reg  sync_dff_0_seip; // @[SoC.scala 127:27]
  reg  sync_dff_1_mtip; // @[SoC.scala 127:27]
  reg  sync_dff_1_msip; // @[SoC.scala 127:27]
  reg  sync_dff_1_meip; // @[SoC.scala 127:27]
  reg  sync_dff_1_seip; // @[SoC.scala 127:27]
  reg  sync_dff_2_mtip; // @[SoC.scala 127:27]
  reg  sync_dff_2_msip; // @[SoC.scala 127:27]
  reg  sync_dff_2_meip; // @[SoC.scala 127:27]
  reg  sync_dff_2_seip; // @[SoC.scala 127:27]
  SoCImp soc_imp ( // @[SoC.scala 81:27]
    .clock(soc_imp_clock),
    .reset(soc_imp_reset),
    .auto_out_a_ready(soc_imp_auto_out_a_ready),
    .auto_out_a_valid(soc_imp_auto_out_a_valid),
    .auto_out_a_bits_opcode(soc_imp_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(soc_imp_auto_out_a_bits_param),
    .auto_out_a_bits_size(soc_imp_auto_out_a_bits_size),
    .auto_out_a_bits_source(soc_imp_auto_out_a_bits_source),
    .auto_out_a_bits_address(soc_imp_auto_out_a_bits_address),
    .auto_out_a_bits_mask(soc_imp_auto_out_a_bits_mask),
    .auto_out_a_bits_data(soc_imp_auto_out_a_bits_data),
    .auto_out_b_ready(soc_imp_auto_out_b_ready),
    .auto_out_b_valid(soc_imp_auto_out_b_valid),
    .auto_out_b_bits_size(soc_imp_auto_out_b_bits_size),
    .auto_out_b_bits_source(soc_imp_auto_out_b_bits_source),
    .auto_out_b_bits_address(soc_imp_auto_out_b_bits_address),
    .auto_out_c_ready(soc_imp_auto_out_c_ready),
    .auto_out_c_valid(soc_imp_auto_out_c_valid),
    .auto_out_c_bits_opcode(soc_imp_auto_out_c_bits_opcode),
    .auto_out_c_bits_param(soc_imp_auto_out_c_bits_param),
    .auto_out_c_bits_size(soc_imp_auto_out_c_bits_size),
    .auto_out_c_bits_source(soc_imp_auto_out_c_bits_source),
    .auto_out_c_bits_address(soc_imp_auto_out_c_bits_address),
    .auto_out_c_bits_data(soc_imp_auto_out_c_bits_data),
    .auto_out_d_ready(soc_imp_auto_out_d_ready),
    .auto_out_d_valid(soc_imp_auto_out_d_valid),
    .auto_out_d_bits_opcode(soc_imp_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(soc_imp_auto_out_d_bits_size),
    .auto_out_d_bits_source(soc_imp_auto_out_d_bits_source),
    .auto_out_d_bits_sink(soc_imp_auto_out_d_bits_sink),
    .auto_out_d_bits_data(soc_imp_auto_out_d_bits_data),
    .auto_out_e_ready(soc_imp_auto_out_e_ready),
    .auto_out_e_valid(soc_imp_auto_out_e_valid),
    .auto_out_e_bits_sink(soc_imp_auto_out_e_bits_sink),
    .io_intr_mtip(soc_imp_io_intr_mtip),
    .io_intr_msip(soc_imp_io_intr_msip),
    .io_intr_meip(soc_imp_io_intr_meip),
    .io_intr_seip(soc_imp_io_intr_seip)
  );
  TLSerdes serdes ( // @[SoC.scala 87:26]
    .clock(serdes_clock),
    .reset(serdes_reset),
    .auto_in_a_ready(serdes_auto_in_a_ready),
    .auto_in_a_valid(serdes_auto_in_a_valid),
    .auto_in_a_bits_opcode(serdes_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(serdes_auto_in_a_bits_param),
    .auto_in_a_bits_size(serdes_auto_in_a_bits_size),
    .auto_in_a_bits_source(serdes_auto_in_a_bits_source),
    .auto_in_a_bits_address(serdes_auto_in_a_bits_address),
    .auto_in_a_bits_mask(serdes_auto_in_a_bits_mask),
    .auto_in_a_bits_data(serdes_auto_in_a_bits_data),
    .auto_in_b_ready(serdes_auto_in_b_ready),
    .auto_in_b_valid(serdes_auto_in_b_valid),
    .auto_in_b_bits_size(serdes_auto_in_b_bits_size),
    .auto_in_b_bits_source(serdes_auto_in_b_bits_source),
    .auto_in_b_bits_address(serdes_auto_in_b_bits_address),
    .auto_in_c_ready(serdes_auto_in_c_ready),
    .auto_in_c_valid(serdes_auto_in_c_valid),
    .auto_in_c_bits_opcode(serdes_auto_in_c_bits_opcode),
    .auto_in_c_bits_param(serdes_auto_in_c_bits_param),
    .auto_in_c_bits_size(serdes_auto_in_c_bits_size),
    .auto_in_c_bits_source(serdes_auto_in_c_bits_source),
    .auto_in_c_bits_address(serdes_auto_in_c_bits_address),
    .auto_in_c_bits_data(serdes_auto_in_c_bits_data),
    .auto_in_d_ready(serdes_auto_in_d_ready),
    .auto_in_d_valid(serdes_auto_in_d_valid),
    .auto_in_d_bits_opcode(serdes_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(serdes_auto_in_d_bits_size),
    .auto_in_d_bits_source(serdes_auto_in_d_bits_source),
    .auto_in_d_bits_sink(serdes_auto_in_d_bits_sink),
    .auto_in_d_bits_data(serdes_auto_in_d_bits_data),
    .auto_in_e_ready(serdes_auto_in_e_ready),
    .auto_in_e_valid(serdes_auto_in_e_valid),
    .auto_in_e_bits_sink(serdes_auto_in_e_bits_sink),
    .io_ser_0_in_ready(serdes_io_ser_0_in_ready),
    .io_ser_0_in_valid(serdes_io_ser_0_in_valid),
    .io_ser_0_in_bits(serdes_io_ser_0_in_bits),
    .io_ser_0_out_ready(serdes_io_ser_0_out_ready),
    .io_ser_0_out_valid(serdes_io_ser_0_out_valid),
    .io_ser_0_out_bits(serdes_io_ser_0_out_bits)
  );
  TLTraceBuffer trace_buffer ( // @[TLTraceBuffer.scala 47:34]
    .clock(trace_buffer_clock),
    .reset(trace_buffer_reset),
    .auto_in_a_ready(trace_buffer_auto_in_a_ready),
    .auto_in_a_valid(trace_buffer_auto_in_a_valid),
    .auto_in_a_bits_opcode(trace_buffer_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(trace_buffer_auto_in_a_bits_param),
    .auto_in_a_bits_size(trace_buffer_auto_in_a_bits_size),
    .auto_in_a_bits_source(trace_buffer_auto_in_a_bits_source),
    .auto_in_a_bits_address(trace_buffer_auto_in_a_bits_address),
    .auto_in_a_bits_mask(trace_buffer_auto_in_a_bits_mask),
    .auto_in_a_bits_data(trace_buffer_auto_in_a_bits_data),
    .auto_in_b_ready(trace_buffer_auto_in_b_ready),
    .auto_in_b_valid(trace_buffer_auto_in_b_valid),
    .auto_in_b_bits_size(trace_buffer_auto_in_b_bits_size),
    .auto_in_b_bits_source(trace_buffer_auto_in_b_bits_source),
    .auto_in_b_bits_address(trace_buffer_auto_in_b_bits_address),
    .auto_in_c_ready(trace_buffer_auto_in_c_ready),
    .auto_in_c_valid(trace_buffer_auto_in_c_valid),
    .auto_in_c_bits_opcode(trace_buffer_auto_in_c_bits_opcode),
    .auto_in_c_bits_param(trace_buffer_auto_in_c_bits_param),
    .auto_in_c_bits_size(trace_buffer_auto_in_c_bits_size),
    .auto_in_c_bits_source(trace_buffer_auto_in_c_bits_source),
    .auto_in_c_bits_address(trace_buffer_auto_in_c_bits_address),
    .auto_in_c_bits_data(trace_buffer_auto_in_c_bits_data),
    .auto_in_d_ready(trace_buffer_auto_in_d_ready),
    .auto_in_d_valid(trace_buffer_auto_in_d_valid),
    .auto_in_d_bits_opcode(trace_buffer_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(trace_buffer_auto_in_d_bits_size),
    .auto_in_d_bits_source(trace_buffer_auto_in_d_bits_source),
    .auto_in_d_bits_sink(trace_buffer_auto_in_d_bits_sink),
    .auto_in_d_bits_data(trace_buffer_auto_in_d_bits_data),
    .auto_in_e_ready(trace_buffer_auto_in_e_ready),
    .auto_in_e_valid(trace_buffer_auto_in_e_valid),
    .auto_in_e_bits_sink(trace_buffer_auto_in_e_bits_sink),
    .auto_out_a_ready(trace_buffer_auto_out_a_ready),
    .auto_out_a_valid(trace_buffer_auto_out_a_valid),
    .auto_out_a_bits_opcode(trace_buffer_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(trace_buffer_auto_out_a_bits_param),
    .auto_out_a_bits_size(trace_buffer_auto_out_a_bits_size),
    .auto_out_a_bits_source(trace_buffer_auto_out_a_bits_source),
    .auto_out_a_bits_address(trace_buffer_auto_out_a_bits_address),
    .auto_out_a_bits_mask(trace_buffer_auto_out_a_bits_mask),
    .auto_out_a_bits_data(trace_buffer_auto_out_a_bits_data),
    .auto_out_b_ready(trace_buffer_auto_out_b_ready),
    .auto_out_b_valid(trace_buffer_auto_out_b_valid),
    .auto_out_b_bits_size(trace_buffer_auto_out_b_bits_size),
    .auto_out_b_bits_source(trace_buffer_auto_out_b_bits_source),
    .auto_out_b_bits_address(trace_buffer_auto_out_b_bits_address),
    .auto_out_c_ready(trace_buffer_auto_out_c_ready),
    .auto_out_c_valid(trace_buffer_auto_out_c_valid),
    .auto_out_c_bits_opcode(trace_buffer_auto_out_c_bits_opcode),
    .auto_out_c_bits_param(trace_buffer_auto_out_c_bits_param),
    .auto_out_c_bits_size(trace_buffer_auto_out_c_bits_size),
    .auto_out_c_bits_source(trace_buffer_auto_out_c_bits_source),
    .auto_out_c_bits_address(trace_buffer_auto_out_c_bits_address),
    .auto_out_c_bits_data(trace_buffer_auto_out_c_bits_data),
    .auto_out_d_ready(trace_buffer_auto_out_d_ready),
    .auto_out_d_valid(trace_buffer_auto_out_d_valid),
    .auto_out_d_bits_opcode(trace_buffer_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(trace_buffer_auto_out_d_bits_size),
    .auto_out_d_bits_source(trace_buffer_auto_out_d_bits_source),
    .auto_out_d_bits_sink(trace_buffer_auto_out_d_bits_sink),
    .auto_out_d_bits_data(trace_buffer_auto_out_d_bits_data),
    .auto_out_e_ready(trace_buffer_auto_out_e_ready),
    .auto_out_e_valid(trace_buffer_auto_out_e_valid),
    .auto_out_e_bits_sink(trace_buffer_auto_out_e_bits_sink)
  );
  AsyncQueue in_fifo ( // @[SoC.scala 111:26]
    .io_enq_clock(in_fifo_io_enq_clock),
    .io_enq_reset(in_fifo_io_enq_reset),
    .io_enq_ready(in_fifo_io_enq_ready),
    .io_enq_valid(in_fifo_io_enq_valid),
    .io_enq_bits(in_fifo_io_enq_bits),
    .io_deq_clock(in_fifo_io_deq_clock),
    .io_deq_reset(in_fifo_io_deq_reset),
    .io_deq_ready(in_fifo_io_deq_ready),
    .io_deq_valid(in_fifo_io_deq_valid),
    .io_deq_bits(in_fifo_io_deq_bits)
  );
  AsyncQueue out_fifo ( // @[SoC.scala 112:26]
    .io_enq_clock(out_fifo_io_enq_clock),
    .io_enq_reset(out_fifo_io_enq_reset),
    .io_enq_ready(out_fifo_io_enq_ready),
    .io_enq_valid(out_fifo_io_enq_valid),
    .io_enq_bits(out_fifo_io_enq_bits),
    .io_deq_clock(out_fifo_io_deq_clock),
    .io_deq_reset(out_fifo_io_deq_reset),
    .io_deq_ready(out_fifo_io_deq_ready),
    .io_deq_valid(out_fifo_io_deq_valid),
    .io_deq_bits(out_fifo_io_deq_bits)
  );
  assign io_in_ready = in_fifo_io_enq_ready; // @[SoC.scala 113:27]
  assign io_out_valid = out_fifo_io_deq_valid; // @[SoC.scala 122:27]
  assign io_out_bits = out_fifo_io_deq_bits; // @[SoC.scala 122:27]
  assign soc_imp_clock = clock;
  assign soc_imp_reset = reset;
  assign soc_imp_auto_out_a_ready = trace_buffer_auto_in_a_ready; // @[LazyModule.scala 355:16]
  assign soc_imp_auto_out_b_valid = trace_buffer_auto_in_b_valid; // @[LazyModule.scala 355:16]
  assign soc_imp_auto_out_b_bits_size = trace_buffer_auto_in_b_bits_size; // @[LazyModule.scala 355:16]
  assign soc_imp_auto_out_b_bits_source = trace_buffer_auto_in_b_bits_source; // @[LazyModule.scala 355:16]
  assign soc_imp_auto_out_b_bits_address = trace_buffer_auto_in_b_bits_address; // @[LazyModule.scala 355:16]
  assign soc_imp_auto_out_c_ready = trace_buffer_auto_in_c_ready; // @[LazyModule.scala 355:16]
  assign soc_imp_auto_out_d_valid = trace_buffer_auto_in_d_valid; // @[LazyModule.scala 355:16]
  assign soc_imp_auto_out_d_bits_opcode = trace_buffer_auto_in_d_bits_opcode; // @[LazyModule.scala 355:16]
  assign soc_imp_auto_out_d_bits_size = trace_buffer_auto_in_d_bits_size; // @[LazyModule.scala 355:16]
  assign soc_imp_auto_out_d_bits_source = trace_buffer_auto_in_d_bits_source; // @[LazyModule.scala 355:16]
  assign soc_imp_auto_out_d_bits_sink = trace_buffer_auto_in_d_bits_sink; // @[LazyModule.scala 355:16]
  assign soc_imp_auto_out_d_bits_data = trace_buffer_auto_in_d_bits_data; // @[LazyModule.scala 355:16]
  assign soc_imp_auto_out_e_ready = trace_buffer_auto_in_e_ready; // @[LazyModule.scala 355:16]
  assign soc_imp_io_intr_mtip = sync_dff_2_mtip; // @[SoC.scala 131:28]
  assign soc_imp_io_intr_msip = sync_dff_2_msip; // @[SoC.scala 131:28]
  assign soc_imp_io_intr_meip = sync_dff_2_meip; // @[SoC.scala 131:28]
  assign soc_imp_io_intr_seip = sync_dff_2_seip; // @[SoC.scala 131:28]
  assign serdes_clock = clock;
  assign serdes_reset = reset;
  assign serdes_auto_in_a_valid = trace_buffer_auto_out_a_valid; // @[LazyModule.scala 353:16]
  assign serdes_auto_in_a_bits_opcode = trace_buffer_auto_out_a_bits_opcode; // @[LazyModule.scala 353:16]
  assign serdes_auto_in_a_bits_param = trace_buffer_auto_out_a_bits_param; // @[LazyModule.scala 353:16]
  assign serdes_auto_in_a_bits_size = trace_buffer_auto_out_a_bits_size; // @[LazyModule.scala 353:16]
  assign serdes_auto_in_a_bits_source = trace_buffer_auto_out_a_bits_source; // @[LazyModule.scala 353:16]
  assign serdes_auto_in_a_bits_address = trace_buffer_auto_out_a_bits_address; // @[LazyModule.scala 353:16]
  assign serdes_auto_in_a_bits_mask = trace_buffer_auto_out_a_bits_mask; // @[LazyModule.scala 353:16]
  assign serdes_auto_in_a_bits_data = trace_buffer_auto_out_a_bits_data; // @[LazyModule.scala 353:16]
  assign serdes_auto_in_b_ready = trace_buffer_auto_out_b_ready; // @[LazyModule.scala 353:16]
  assign serdes_auto_in_c_valid = trace_buffer_auto_out_c_valid; // @[LazyModule.scala 353:16]
  assign serdes_auto_in_c_bits_opcode = trace_buffer_auto_out_c_bits_opcode; // @[LazyModule.scala 353:16]
  assign serdes_auto_in_c_bits_param = trace_buffer_auto_out_c_bits_param; // @[LazyModule.scala 353:16]
  assign serdes_auto_in_c_bits_size = trace_buffer_auto_out_c_bits_size; // @[LazyModule.scala 353:16]
  assign serdes_auto_in_c_bits_source = trace_buffer_auto_out_c_bits_source; // @[LazyModule.scala 353:16]
  assign serdes_auto_in_c_bits_address = trace_buffer_auto_out_c_bits_address; // @[LazyModule.scala 353:16]
  assign serdes_auto_in_c_bits_data = trace_buffer_auto_out_c_bits_data; // @[LazyModule.scala 353:16]
  assign serdes_auto_in_d_ready = trace_buffer_auto_out_d_ready; // @[LazyModule.scala 353:16]
  assign serdes_auto_in_e_valid = trace_buffer_auto_out_e_valid; // @[LazyModule.scala 353:16]
  assign serdes_auto_in_e_bits_sink = trace_buffer_auto_out_e_bits_sink; // @[LazyModule.scala 353:16]
  assign serdes_io_ser_0_in_valid = in_fifo_io_deq_valid; // @[SoC.scala 116:27]
  assign serdes_io_ser_0_in_bits = in_fifo_io_deq_bits; // @[SoC.scala 116:27]
  assign serdes_io_ser_0_out_ready = out_fifo_io_enq_ready; // @[SoC.scala 119:27]
  assign trace_buffer_clock = clock;
  assign trace_buffer_reset = reset;
  assign trace_buffer_auto_in_a_valid = soc_imp_auto_out_a_valid; // @[LazyModule.scala 355:16]
  assign trace_buffer_auto_in_a_bits_opcode = soc_imp_auto_out_a_bits_opcode; // @[LazyModule.scala 355:16]
  assign trace_buffer_auto_in_a_bits_param = soc_imp_auto_out_a_bits_param; // @[LazyModule.scala 355:16]
  assign trace_buffer_auto_in_a_bits_size = soc_imp_auto_out_a_bits_size; // @[LazyModule.scala 355:16]
  assign trace_buffer_auto_in_a_bits_source = soc_imp_auto_out_a_bits_source; // @[LazyModule.scala 355:16]
  assign trace_buffer_auto_in_a_bits_address = soc_imp_auto_out_a_bits_address; // @[LazyModule.scala 355:16]
  assign trace_buffer_auto_in_a_bits_mask = soc_imp_auto_out_a_bits_mask; // @[LazyModule.scala 355:16]
  assign trace_buffer_auto_in_a_bits_data = soc_imp_auto_out_a_bits_data; // @[LazyModule.scala 355:16]
  assign trace_buffer_auto_in_b_ready = soc_imp_auto_out_b_ready; // @[LazyModule.scala 355:16]
  assign trace_buffer_auto_in_c_valid = soc_imp_auto_out_c_valid; // @[LazyModule.scala 355:16]
  assign trace_buffer_auto_in_c_bits_opcode = soc_imp_auto_out_c_bits_opcode; // @[LazyModule.scala 355:16]
  assign trace_buffer_auto_in_c_bits_param = soc_imp_auto_out_c_bits_param; // @[LazyModule.scala 355:16]
  assign trace_buffer_auto_in_c_bits_size = soc_imp_auto_out_c_bits_size; // @[LazyModule.scala 355:16]
  assign trace_buffer_auto_in_c_bits_source = soc_imp_auto_out_c_bits_source; // @[LazyModule.scala 355:16]
  assign trace_buffer_auto_in_c_bits_address = soc_imp_auto_out_c_bits_address; // @[LazyModule.scala 355:16]
  assign trace_buffer_auto_in_c_bits_data = soc_imp_auto_out_c_bits_data; // @[LazyModule.scala 355:16]
  assign trace_buffer_auto_in_d_ready = soc_imp_auto_out_d_ready; // @[LazyModule.scala 355:16]
  assign trace_buffer_auto_in_e_valid = soc_imp_auto_out_e_valid; // @[LazyModule.scala 355:16]
  assign trace_buffer_auto_in_e_bits_sink = soc_imp_auto_out_e_bits_sink; // @[LazyModule.scala 355:16]
  assign trace_buffer_auto_out_a_ready = serdes_auto_in_a_ready; // @[LazyModule.scala 353:16]
  assign trace_buffer_auto_out_b_valid = serdes_auto_in_b_valid; // @[LazyModule.scala 353:16]
  assign trace_buffer_auto_out_b_bits_size = serdes_auto_in_b_bits_size; // @[LazyModule.scala 353:16]
  assign trace_buffer_auto_out_b_bits_source = serdes_auto_in_b_bits_source; // @[LazyModule.scala 353:16]
  assign trace_buffer_auto_out_b_bits_address = serdes_auto_in_b_bits_address; // @[LazyModule.scala 353:16]
  assign trace_buffer_auto_out_c_ready = serdes_auto_in_c_ready; // @[LazyModule.scala 353:16]
  assign trace_buffer_auto_out_d_valid = serdes_auto_in_d_valid; // @[LazyModule.scala 353:16]
  assign trace_buffer_auto_out_d_bits_opcode = serdes_auto_in_d_bits_opcode; // @[LazyModule.scala 353:16]
  assign trace_buffer_auto_out_d_bits_size = serdes_auto_in_d_bits_size; // @[LazyModule.scala 353:16]
  assign trace_buffer_auto_out_d_bits_source = serdes_auto_in_d_bits_source; // @[LazyModule.scala 353:16]
  assign trace_buffer_auto_out_d_bits_sink = serdes_auto_in_d_bits_sink; // @[LazyModule.scala 353:16]
  assign trace_buffer_auto_out_d_bits_data = serdes_auto_in_d_bits_data; // @[LazyModule.scala 353:16]
  assign trace_buffer_auto_out_e_ready = serdes_auto_in_e_ready; // @[LazyModule.scala 353:16]
  assign in_fifo_io_enq_clock = io_io_clock; // @[SoC.scala 114:27]
  assign in_fifo_io_enq_reset = io_io_reset; // @[SoC.scala 115:27]
  assign in_fifo_io_enq_valid = io_in_valid; // @[SoC.scala 113:27]
  assign in_fifo_io_enq_bits = io_in_bits; // @[SoC.scala 113:27]
  assign in_fifo_io_deq_clock = clock; // @[SoC.scala 117:27]
  assign in_fifo_io_deq_reset = reset; // @[SoC.scala 118:27]
  assign in_fifo_io_deq_ready = serdes_io_ser_0_in_ready; // @[SoC.scala 116:27]
  assign out_fifo_io_enq_clock = clock; // @[SoC.scala 120:27]
  assign out_fifo_io_enq_reset = reset; // @[SoC.scala 121:27]
  assign out_fifo_io_enq_valid = serdes_io_ser_0_out_valid; // @[SoC.scala 119:27]
  assign out_fifo_io_enq_bits = serdes_io_ser_0_out_bits; // @[SoC.scala 119:27]
  assign out_fifo_io_deq_clock = io_io_clock; // @[SoC.scala 123:27]
  assign out_fifo_io_deq_reset = io_io_reset; // @[SoC.scala 124:27]
  assign out_fifo_io_deq_ready = io_out_ready; // @[SoC.scala 122:27]
  always @(posedge clock) begin
    if (reset) begin // @[SoC.scala 127:27]
      sync_dff_0_mtip <= 1'h0; // @[SoC.scala 127:27]
    end else begin
      sync_dff_0_mtip <= io_intr_mtip; // @[SoC.scala 128:28]
    end
    if (reset) begin // @[SoC.scala 127:27]
      sync_dff_0_msip <= 1'h0; // @[SoC.scala 127:27]
    end else begin
      sync_dff_0_msip <= io_intr_msip; // @[SoC.scala 128:28]
    end
    if (reset) begin // @[SoC.scala 127:27]
      sync_dff_0_meip <= 1'h0; // @[SoC.scala 127:27]
    end else begin
      sync_dff_0_meip <= io_intr_meip; // @[SoC.scala 128:28]
    end
    if (reset) begin // @[SoC.scala 127:27]
      sync_dff_0_seip <= 1'h0; // @[SoC.scala 127:27]
    end else begin
      sync_dff_0_seip <= io_intr_seip; // @[SoC.scala 128:28]
    end
    if (reset) begin // @[SoC.scala 127:27]
      sync_dff_1_mtip <= 1'h0; // @[SoC.scala 127:27]
    end else begin
      sync_dff_1_mtip <= sync_dff_0_mtip; // @[SoC.scala 129:28]
    end
    if (reset) begin // @[SoC.scala 127:27]
      sync_dff_1_msip <= 1'h0; // @[SoC.scala 127:27]
    end else begin
      sync_dff_1_msip <= sync_dff_0_msip; // @[SoC.scala 129:28]
    end
    if (reset) begin // @[SoC.scala 127:27]
      sync_dff_1_meip <= 1'h0; // @[SoC.scala 127:27]
    end else begin
      sync_dff_1_meip <= sync_dff_0_meip; // @[SoC.scala 129:28]
    end
    if (reset) begin // @[SoC.scala 127:27]
      sync_dff_1_seip <= 1'h0; // @[SoC.scala 127:27]
    end else begin
      sync_dff_1_seip <= sync_dff_0_seip; // @[SoC.scala 129:28]
    end
    if (reset) begin // @[SoC.scala 127:27]
      sync_dff_2_mtip <= 1'h0; // @[SoC.scala 127:27]
    end else begin
      sync_dff_2_mtip <= sync_dff_1_mtip; // @[SoC.scala 130:28]
    end
    if (reset) begin // @[SoC.scala 127:27]
      sync_dff_2_msip <= 1'h0; // @[SoC.scala 127:27]
    end else begin
      sync_dff_2_msip <= sync_dff_1_msip; // @[SoC.scala 130:28]
    end
    if (reset) begin // @[SoC.scala 127:27]
      sync_dff_2_meip <= 1'h0; // @[SoC.scala 127:27]
    end else begin
      sync_dff_2_meip <= sync_dff_1_meip; // @[SoC.scala 130:28]
    end
    if (reset) begin // @[SoC.scala 127:27]
      sync_dff_2_seip <= 1'h0; // @[SoC.scala 127:27]
    end else begin
      sync_dff_2_seip <= sync_dff_1_seip; // @[SoC.scala 130:28]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sync_dff_0_mtip = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  sync_dff_0_msip = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  sync_dff_0_meip = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  sync_dff_0_seip = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  sync_dff_1_mtip = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  sync_dff_1_msip = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  sync_dff_1_meip = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  sync_dff_1_seip = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  sync_dff_2_mtip = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  sync_dff_2_msip = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  sync_dff_2_meip = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  sync_dff_2_seip = _RAND_11[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
