module SRAM(
  input          clock,
  input          io_en,
  input  [9:0]   io_addr,
  input  [272:0] io_wdata,
  input          io_wen,
  output [272:0] io_rdata
);
`ifdef RANDOMIZE_MEM_INIT
  reg [287:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [272:0] array [0:1023]; // @[SRAM.scala 13:26]
  wire  array_io_rdata_MPORT_en; // @[SRAM.scala 13:26]
  wire [9:0] array_io_rdata_MPORT_addr; // @[SRAM.scala 13:26]
  wire [272:0] array_io_rdata_MPORT_data; // @[SRAM.scala 13:26]
  wire [272:0] array_MPORT_data; // @[SRAM.scala 13:26]
  wire [9:0] array_MPORT_addr; // @[SRAM.scala 13:26]
  wire  array_MPORT_mask; // @[SRAM.scala 13:26]
  wire  array_MPORT_en; // @[SRAM.scala 13:26]
  reg  array_io_rdata_MPORT_en_pipe_0;
  reg [9:0] array_io_rdata_MPORT_addr_pipe_0;
  reg  io_rdata_REG; // @[SRAM.scala 15:26]
  assign array_io_rdata_MPORT_en = array_io_rdata_MPORT_en_pipe_0;
  assign array_io_rdata_MPORT_addr = array_io_rdata_MPORT_addr_pipe_0;
  assign array_io_rdata_MPORT_data = array[array_io_rdata_MPORT_addr]; // @[SRAM.scala 13:26]
  assign array_MPORT_data = io_wdata;
  assign array_MPORT_addr = io_addr;
  assign array_MPORT_mask = 1'h1;
  assign array_MPORT_en = io_en & io_wen;
  assign io_rdata = io_rdata_REG ? array_io_rdata_MPORT_data : 273'h0; // @[SRAM.scala 15:18]
  always @(posedge clock) begin
    if (array_MPORT_en & array_MPORT_mask) begin
      array[array_MPORT_addr] <= array_MPORT_data; // @[SRAM.scala 13:26]
    end
    array_io_rdata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      array_io_rdata_MPORT_addr_pipe_0 <= io_addr;
    end
    io_rdata_REG <= io_en; // @[SRAM.scala 15:26]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {9{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    array[initvar] = _RAND_0[272:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  array_io_rdata_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  array_io_rdata_MPORT_addr_pipe_0 = _RAND_2[9:0];
  _RAND_3 = {1{`RANDOM}};
  io_rdata_REG = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ICache(
  input          clock,
  input          reset,
  input          auto_out_a_ready,
  output         auto_out_a_valid,
  output [1:0]   auto_out_a_bits_source,
  output [31:0]  auto_out_a_bits_address,
  output         auto_out_d_ready,
  input          auto_out_d_valid,
  input  [255:0] auto_out_d_bits_data,
  output         io_cache_req_ready,
  input          io_cache_req_valid,
  input  [38:0]  io_cache_req_bits_addr,
  input          io_cache_resp_ready,
  output         io_cache_resp_valid,
  output [63:0]  io_cache_resp_bits_rdata,
  input          io_fence_i
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [287:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [63:0] _RAND_1029;
  reg [255:0] _RAND_1030;
  reg [31:0] _RAND_1031;
`endif // RANDOMIZE_REG_INIT
  wire  array_clock; // @[ICache.scala 50:21]
  wire  array_io_en; // @[ICache.scala 50:21]
  wire [9:0] array_io_addr; // @[ICache.scala 50:21]
  wire [272:0] array_io_wdata; // @[ICache.scala 50:21]
  wire  array_io_wen; // @[ICache.scala 50:21]
  wire [272:0] array_io_rdata; // @[ICache.scala 50:21]
  reg [38:0] req_r_addr; // @[ICache.scala 48:22]
  reg  valid_0; // @[ICache.scala 51:22]
  reg  valid_1; // @[ICache.scala 51:22]
  reg  valid_2; // @[ICache.scala 51:22]
  reg  valid_3; // @[ICache.scala 51:22]
  reg  valid_4; // @[ICache.scala 51:22]
  reg  valid_5; // @[ICache.scala 51:22]
  reg  valid_6; // @[ICache.scala 51:22]
  reg  valid_7; // @[ICache.scala 51:22]
  reg  valid_8; // @[ICache.scala 51:22]
  reg  valid_9; // @[ICache.scala 51:22]
  reg  valid_10; // @[ICache.scala 51:22]
  reg  valid_11; // @[ICache.scala 51:22]
  reg  valid_12; // @[ICache.scala 51:22]
  reg  valid_13; // @[ICache.scala 51:22]
  reg  valid_14; // @[ICache.scala 51:22]
  reg  valid_15; // @[ICache.scala 51:22]
  reg  valid_16; // @[ICache.scala 51:22]
  reg  valid_17; // @[ICache.scala 51:22]
  reg  valid_18; // @[ICache.scala 51:22]
  reg  valid_19; // @[ICache.scala 51:22]
  reg  valid_20; // @[ICache.scala 51:22]
  reg  valid_21; // @[ICache.scala 51:22]
  reg  valid_22; // @[ICache.scala 51:22]
  reg  valid_23; // @[ICache.scala 51:22]
  reg  valid_24; // @[ICache.scala 51:22]
  reg  valid_25; // @[ICache.scala 51:22]
  reg  valid_26; // @[ICache.scala 51:22]
  reg  valid_27; // @[ICache.scala 51:22]
  reg  valid_28; // @[ICache.scala 51:22]
  reg  valid_29; // @[ICache.scala 51:22]
  reg  valid_30; // @[ICache.scala 51:22]
  reg  valid_31; // @[ICache.scala 51:22]
  reg  valid_32; // @[ICache.scala 51:22]
  reg  valid_33; // @[ICache.scala 51:22]
  reg  valid_34; // @[ICache.scala 51:22]
  reg  valid_35; // @[ICache.scala 51:22]
  reg  valid_36; // @[ICache.scala 51:22]
  reg  valid_37; // @[ICache.scala 51:22]
  reg  valid_38; // @[ICache.scala 51:22]
  reg  valid_39; // @[ICache.scala 51:22]
  reg  valid_40; // @[ICache.scala 51:22]
  reg  valid_41; // @[ICache.scala 51:22]
  reg  valid_42; // @[ICache.scala 51:22]
  reg  valid_43; // @[ICache.scala 51:22]
  reg  valid_44; // @[ICache.scala 51:22]
  reg  valid_45; // @[ICache.scala 51:22]
  reg  valid_46; // @[ICache.scala 51:22]
  reg  valid_47; // @[ICache.scala 51:22]
  reg  valid_48; // @[ICache.scala 51:22]
  reg  valid_49; // @[ICache.scala 51:22]
  reg  valid_50; // @[ICache.scala 51:22]
  reg  valid_51; // @[ICache.scala 51:22]
  reg  valid_52; // @[ICache.scala 51:22]
  reg  valid_53; // @[ICache.scala 51:22]
  reg  valid_54; // @[ICache.scala 51:22]
  reg  valid_55; // @[ICache.scala 51:22]
  reg  valid_56; // @[ICache.scala 51:22]
  reg  valid_57; // @[ICache.scala 51:22]
  reg  valid_58; // @[ICache.scala 51:22]
  reg  valid_59; // @[ICache.scala 51:22]
  reg  valid_60; // @[ICache.scala 51:22]
  reg  valid_61; // @[ICache.scala 51:22]
  reg  valid_62; // @[ICache.scala 51:22]
  reg  valid_63; // @[ICache.scala 51:22]
  reg  valid_64; // @[ICache.scala 51:22]
  reg  valid_65; // @[ICache.scala 51:22]
  reg  valid_66; // @[ICache.scala 51:22]
  reg  valid_67; // @[ICache.scala 51:22]
  reg  valid_68; // @[ICache.scala 51:22]
  reg  valid_69; // @[ICache.scala 51:22]
  reg  valid_70; // @[ICache.scala 51:22]
  reg  valid_71; // @[ICache.scala 51:22]
  reg  valid_72; // @[ICache.scala 51:22]
  reg  valid_73; // @[ICache.scala 51:22]
  reg  valid_74; // @[ICache.scala 51:22]
  reg  valid_75; // @[ICache.scala 51:22]
  reg  valid_76; // @[ICache.scala 51:22]
  reg  valid_77; // @[ICache.scala 51:22]
  reg  valid_78; // @[ICache.scala 51:22]
  reg  valid_79; // @[ICache.scala 51:22]
  reg  valid_80; // @[ICache.scala 51:22]
  reg  valid_81; // @[ICache.scala 51:22]
  reg  valid_82; // @[ICache.scala 51:22]
  reg  valid_83; // @[ICache.scala 51:22]
  reg  valid_84; // @[ICache.scala 51:22]
  reg  valid_85; // @[ICache.scala 51:22]
  reg  valid_86; // @[ICache.scala 51:22]
  reg  valid_87; // @[ICache.scala 51:22]
  reg  valid_88; // @[ICache.scala 51:22]
  reg  valid_89; // @[ICache.scala 51:22]
  reg  valid_90; // @[ICache.scala 51:22]
  reg  valid_91; // @[ICache.scala 51:22]
  reg  valid_92; // @[ICache.scala 51:22]
  reg  valid_93; // @[ICache.scala 51:22]
  reg  valid_94; // @[ICache.scala 51:22]
  reg  valid_95; // @[ICache.scala 51:22]
  reg  valid_96; // @[ICache.scala 51:22]
  reg  valid_97; // @[ICache.scala 51:22]
  reg  valid_98; // @[ICache.scala 51:22]
  reg  valid_99; // @[ICache.scala 51:22]
  reg  valid_100; // @[ICache.scala 51:22]
  reg  valid_101; // @[ICache.scala 51:22]
  reg  valid_102; // @[ICache.scala 51:22]
  reg  valid_103; // @[ICache.scala 51:22]
  reg  valid_104; // @[ICache.scala 51:22]
  reg  valid_105; // @[ICache.scala 51:22]
  reg  valid_106; // @[ICache.scala 51:22]
  reg  valid_107; // @[ICache.scala 51:22]
  reg  valid_108; // @[ICache.scala 51:22]
  reg  valid_109; // @[ICache.scala 51:22]
  reg  valid_110; // @[ICache.scala 51:22]
  reg  valid_111; // @[ICache.scala 51:22]
  reg  valid_112; // @[ICache.scala 51:22]
  reg  valid_113; // @[ICache.scala 51:22]
  reg  valid_114; // @[ICache.scala 51:22]
  reg  valid_115; // @[ICache.scala 51:22]
  reg  valid_116; // @[ICache.scala 51:22]
  reg  valid_117; // @[ICache.scala 51:22]
  reg  valid_118; // @[ICache.scala 51:22]
  reg  valid_119; // @[ICache.scala 51:22]
  reg  valid_120; // @[ICache.scala 51:22]
  reg  valid_121; // @[ICache.scala 51:22]
  reg  valid_122; // @[ICache.scala 51:22]
  reg  valid_123; // @[ICache.scala 51:22]
  reg  valid_124; // @[ICache.scala 51:22]
  reg  valid_125; // @[ICache.scala 51:22]
  reg  valid_126; // @[ICache.scala 51:22]
  reg  valid_127; // @[ICache.scala 51:22]
  reg  valid_128; // @[ICache.scala 51:22]
  reg  valid_129; // @[ICache.scala 51:22]
  reg  valid_130; // @[ICache.scala 51:22]
  reg  valid_131; // @[ICache.scala 51:22]
  reg  valid_132; // @[ICache.scala 51:22]
  reg  valid_133; // @[ICache.scala 51:22]
  reg  valid_134; // @[ICache.scala 51:22]
  reg  valid_135; // @[ICache.scala 51:22]
  reg  valid_136; // @[ICache.scala 51:22]
  reg  valid_137; // @[ICache.scala 51:22]
  reg  valid_138; // @[ICache.scala 51:22]
  reg  valid_139; // @[ICache.scala 51:22]
  reg  valid_140; // @[ICache.scala 51:22]
  reg  valid_141; // @[ICache.scala 51:22]
  reg  valid_142; // @[ICache.scala 51:22]
  reg  valid_143; // @[ICache.scala 51:22]
  reg  valid_144; // @[ICache.scala 51:22]
  reg  valid_145; // @[ICache.scala 51:22]
  reg  valid_146; // @[ICache.scala 51:22]
  reg  valid_147; // @[ICache.scala 51:22]
  reg  valid_148; // @[ICache.scala 51:22]
  reg  valid_149; // @[ICache.scala 51:22]
  reg  valid_150; // @[ICache.scala 51:22]
  reg  valid_151; // @[ICache.scala 51:22]
  reg  valid_152; // @[ICache.scala 51:22]
  reg  valid_153; // @[ICache.scala 51:22]
  reg  valid_154; // @[ICache.scala 51:22]
  reg  valid_155; // @[ICache.scala 51:22]
  reg  valid_156; // @[ICache.scala 51:22]
  reg  valid_157; // @[ICache.scala 51:22]
  reg  valid_158; // @[ICache.scala 51:22]
  reg  valid_159; // @[ICache.scala 51:22]
  reg  valid_160; // @[ICache.scala 51:22]
  reg  valid_161; // @[ICache.scala 51:22]
  reg  valid_162; // @[ICache.scala 51:22]
  reg  valid_163; // @[ICache.scala 51:22]
  reg  valid_164; // @[ICache.scala 51:22]
  reg  valid_165; // @[ICache.scala 51:22]
  reg  valid_166; // @[ICache.scala 51:22]
  reg  valid_167; // @[ICache.scala 51:22]
  reg  valid_168; // @[ICache.scala 51:22]
  reg  valid_169; // @[ICache.scala 51:22]
  reg  valid_170; // @[ICache.scala 51:22]
  reg  valid_171; // @[ICache.scala 51:22]
  reg  valid_172; // @[ICache.scala 51:22]
  reg  valid_173; // @[ICache.scala 51:22]
  reg  valid_174; // @[ICache.scala 51:22]
  reg  valid_175; // @[ICache.scala 51:22]
  reg  valid_176; // @[ICache.scala 51:22]
  reg  valid_177; // @[ICache.scala 51:22]
  reg  valid_178; // @[ICache.scala 51:22]
  reg  valid_179; // @[ICache.scala 51:22]
  reg  valid_180; // @[ICache.scala 51:22]
  reg  valid_181; // @[ICache.scala 51:22]
  reg  valid_182; // @[ICache.scala 51:22]
  reg  valid_183; // @[ICache.scala 51:22]
  reg  valid_184; // @[ICache.scala 51:22]
  reg  valid_185; // @[ICache.scala 51:22]
  reg  valid_186; // @[ICache.scala 51:22]
  reg  valid_187; // @[ICache.scala 51:22]
  reg  valid_188; // @[ICache.scala 51:22]
  reg  valid_189; // @[ICache.scala 51:22]
  reg  valid_190; // @[ICache.scala 51:22]
  reg  valid_191; // @[ICache.scala 51:22]
  reg  valid_192; // @[ICache.scala 51:22]
  reg  valid_193; // @[ICache.scala 51:22]
  reg  valid_194; // @[ICache.scala 51:22]
  reg  valid_195; // @[ICache.scala 51:22]
  reg  valid_196; // @[ICache.scala 51:22]
  reg  valid_197; // @[ICache.scala 51:22]
  reg  valid_198; // @[ICache.scala 51:22]
  reg  valid_199; // @[ICache.scala 51:22]
  reg  valid_200; // @[ICache.scala 51:22]
  reg  valid_201; // @[ICache.scala 51:22]
  reg  valid_202; // @[ICache.scala 51:22]
  reg  valid_203; // @[ICache.scala 51:22]
  reg  valid_204; // @[ICache.scala 51:22]
  reg  valid_205; // @[ICache.scala 51:22]
  reg  valid_206; // @[ICache.scala 51:22]
  reg  valid_207; // @[ICache.scala 51:22]
  reg  valid_208; // @[ICache.scala 51:22]
  reg  valid_209; // @[ICache.scala 51:22]
  reg  valid_210; // @[ICache.scala 51:22]
  reg  valid_211; // @[ICache.scala 51:22]
  reg  valid_212; // @[ICache.scala 51:22]
  reg  valid_213; // @[ICache.scala 51:22]
  reg  valid_214; // @[ICache.scala 51:22]
  reg  valid_215; // @[ICache.scala 51:22]
  reg  valid_216; // @[ICache.scala 51:22]
  reg  valid_217; // @[ICache.scala 51:22]
  reg  valid_218; // @[ICache.scala 51:22]
  reg  valid_219; // @[ICache.scala 51:22]
  reg  valid_220; // @[ICache.scala 51:22]
  reg  valid_221; // @[ICache.scala 51:22]
  reg  valid_222; // @[ICache.scala 51:22]
  reg  valid_223; // @[ICache.scala 51:22]
  reg  valid_224; // @[ICache.scala 51:22]
  reg  valid_225; // @[ICache.scala 51:22]
  reg  valid_226; // @[ICache.scala 51:22]
  reg  valid_227; // @[ICache.scala 51:22]
  reg  valid_228; // @[ICache.scala 51:22]
  reg  valid_229; // @[ICache.scala 51:22]
  reg  valid_230; // @[ICache.scala 51:22]
  reg  valid_231; // @[ICache.scala 51:22]
  reg  valid_232; // @[ICache.scala 51:22]
  reg  valid_233; // @[ICache.scala 51:22]
  reg  valid_234; // @[ICache.scala 51:22]
  reg  valid_235; // @[ICache.scala 51:22]
  reg  valid_236; // @[ICache.scala 51:22]
  reg  valid_237; // @[ICache.scala 51:22]
  reg  valid_238; // @[ICache.scala 51:22]
  reg  valid_239; // @[ICache.scala 51:22]
  reg  valid_240; // @[ICache.scala 51:22]
  reg  valid_241; // @[ICache.scala 51:22]
  reg  valid_242; // @[ICache.scala 51:22]
  reg  valid_243; // @[ICache.scala 51:22]
  reg  valid_244; // @[ICache.scala 51:22]
  reg  valid_245; // @[ICache.scala 51:22]
  reg  valid_246; // @[ICache.scala 51:22]
  reg  valid_247; // @[ICache.scala 51:22]
  reg  valid_248; // @[ICache.scala 51:22]
  reg  valid_249; // @[ICache.scala 51:22]
  reg  valid_250; // @[ICache.scala 51:22]
  reg  valid_251; // @[ICache.scala 51:22]
  reg  valid_252; // @[ICache.scala 51:22]
  reg  valid_253; // @[ICache.scala 51:22]
  reg  valid_254; // @[ICache.scala 51:22]
  reg  valid_255; // @[ICache.scala 51:22]
  reg  valid_256; // @[ICache.scala 51:22]
  reg  valid_257; // @[ICache.scala 51:22]
  reg  valid_258; // @[ICache.scala 51:22]
  reg  valid_259; // @[ICache.scala 51:22]
  reg  valid_260; // @[ICache.scala 51:22]
  reg  valid_261; // @[ICache.scala 51:22]
  reg  valid_262; // @[ICache.scala 51:22]
  reg  valid_263; // @[ICache.scala 51:22]
  reg  valid_264; // @[ICache.scala 51:22]
  reg  valid_265; // @[ICache.scala 51:22]
  reg  valid_266; // @[ICache.scala 51:22]
  reg  valid_267; // @[ICache.scala 51:22]
  reg  valid_268; // @[ICache.scala 51:22]
  reg  valid_269; // @[ICache.scala 51:22]
  reg  valid_270; // @[ICache.scala 51:22]
  reg  valid_271; // @[ICache.scala 51:22]
  reg  valid_272; // @[ICache.scala 51:22]
  reg  valid_273; // @[ICache.scala 51:22]
  reg  valid_274; // @[ICache.scala 51:22]
  reg  valid_275; // @[ICache.scala 51:22]
  reg  valid_276; // @[ICache.scala 51:22]
  reg  valid_277; // @[ICache.scala 51:22]
  reg  valid_278; // @[ICache.scala 51:22]
  reg  valid_279; // @[ICache.scala 51:22]
  reg  valid_280; // @[ICache.scala 51:22]
  reg  valid_281; // @[ICache.scala 51:22]
  reg  valid_282; // @[ICache.scala 51:22]
  reg  valid_283; // @[ICache.scala 51:22]
  reg  valid_284; // @[ICache.scala 51:22]
  reg  valid_285; // @[ICache.scala 51:22]
  reg  valid_286; // @[ICache.scala 51:22]
  reg  valid_287; // @[ICache.scala 51:22]
  reg  valid_288; // @[ICache.scala 51:22]
  reg  valid_289; // @[ICache.scala 51:22]
  reg  valid_290; // @[ICache.scala 51:22]
  reg  valid_291; // @[ICache.scala 51:22]
  reg  valid_292; // @[ICache.scala 51:22]
  reg  valid_293; // @[ICache.scala 51:22]
  reg  valid_294; // @[ICache.scala 51:22]
  reg  valid_295; // @[ICache.scala 51:22]
  reg  valid_296; // @[ICache.scala 51:22]
  reg  valid_297; // @[ICache.scala 51:22]
  reg  valid_298; // @[ICache.scala 51:22]
  reg  valid_299; // @[ICache.scala 51:22]
  reg  valid_300; // @[ICache.scala 51:22]
  reg  valid_301; // @[ICache.scala 51:22]
  reg  valid_302; // @[ICache.scala 51:22]
  reg  valid_303; // @[ICache.scala 51:22]
  reg  valid_304; // @[ICache.scala 51:22]
  reg  valid_305; // @[ICache.scala 51:22]
  reg  valid_306; // @[ICache.scala 51:22]
  reg  valid_307; // @[ICache.scala 51:22]
  reg  valid_308; // @[ICache.scala 51:22]
  reg  valid_309; // @[ICache.scala 51:22]
  reg  valid_310; // @[ICache.scala 51:22]
  reg  valid_311; // @[ICache.scala 51:22]
  reg  valid_312; // @[ICache.scala 51:22]
  reg  valid_313; // @[ICache.scala 51:22]
  reg  valid_314; // @[ICache.scala 51:22]
  reg  valid_315; // @[ICache.scala 51:22]
  reg  valid_316; // @[ICache.scala 51:22]
  reg  valid_317; // @[ICache.scala 51:22]
  reg  valid_318; // @[ICache.scala 51:22]
  reg  valid_319; // @[ICache.scala 51:22]
  reg  valid_320; // @[ICache.scala 51:22]
  reg  valid_321; // @[ICache.scala 51:22]
  reg  valid_322; // @[ICache.scala 51:22]
  reg  valid_323; // @[ICache.scala 51:22]
  reg  valid_324; // @[ICache.scala 51:22]
  reg  valid_325; // @[ICache.scala 51:22]
  reg  valid_326; // @[ICache.scala 51:22]
  reg  valid_327; // @[ICache.scala 51:22]
  reg  valid_328; // @[ICache.scala 51:22]
  reg  valid_329; // @[ICache.scala 51:22]
  reg  valid_330; // @[ICache.scala 51:22]
  reg  valid_331; // @[ICache.scala 51:22]
  reg  valid_332; // @[ICache.scala 51:22]
  reg  valid_333; // @[ICache.scala 51:22]
  reg  valid_334; // @[ICache.scala 51:22]
  reg  valid_335; // @[ICache.scala 51:22]
  reg  valid_336; // @[ICache.scala 51:22]
  reg  valid_337; // @[ICache.scala 51:22]
  reg  valid_338; // @[ICache.scala 51:22]
  reg  valid_339; // @[ICache.scala 51:22]
  reg  valid_340; // @[ICache.scala 51:22]
  reg  valid_341; // @[ICache.scala 51:22]
  reg  valid_342; // @[ICache.scala 51:22]
  reg  valid_343; // @[ICache.scala 51:22]
  reg  valid_344; // @[ICache.scala 51:22]
  reg  valid_345; // @[ICache.scala 51:22]
  reg  valid_346; // @[ICache.scala 51:22]
  reg  valid_347; // @[ICache.scala 51:22]
  reg  valid_348; // @[ICache.scala 51:22]
  reg  valid_349; // @[ICache.scala 51:22]
  reg  valid_350; // @[ICache.scala 51:22]
  reg  valid_351; // @[ICache.scala 51:22]
  reg  valid_352; // @[ICache.scala 51:22]
  reg  valid_353; // @[ICache.scala 51:22]
  reg  valid_354; // @[ICache.scala 51:22]
  reg  valid_355; // @[ICache.scala 51:22]
  reg  valid_356; // @[ICache.scala 51:22]
  reg  valid_357; // @[ICache.scala 51:22]
  reg  valid_358; // @[ICache.scala 51:22]
  reg  valid_359; // @[ICache.scala 51:22]
  reg  valid_360; // @[ICache.scala 51:22]
  reg  valid_361; // @[ICache.scala 51:22]
  reg  valid_362; // @[ICache.scala 51:22]
  reg  valid_363; // @[ICache.scala 51:22]
  reg  valid_364; // @[ICache.scala 51:22]
  reg  valid_365; // @[ICache.scala 51:22]
  reg  valid_366; // @[ICache.scala 51:22]
  reg  valid_367; // @[ICache.scala 51:22]
  reg  valid_368; // @[ICache.scala 51:22]
  reg  valid_369; // @[ICache.scala 51:22]
  reg  valid_370; // @[ICache.scala 51:22]
  reg  valid_371; // @[ICache.scala 51:22]
  reg  valid_372; // @[ICache.scala 51:22]
  reg  valid_373; // @[ICache.scala 51:22]
  reg  valid_374; // @[ICache.scala 51:22]
  reg  valid_375; // @[ICache.scala 51:22]
  reg  valid_376; // @[ICache.scala 51:22]
  reg  valid_377; // @[ICache.scala 51:22]
  reg  valid_378; // @[ICache.scala 51:22]
  reg  valid_379; // @[ICache.scala 51:22]
  reg  valid_380; // @[ICache.scala 51:22]
  reg  valid_381; // @[ICache.scala 51:22]
  reg  valid_382; // @[ICache.scala 51:22]
  reg  valid_383; // @[ICache.scala 51:22]
  reg  valid_384; // @[ICache.scala 51:22]
  reg  valid_385; // @[ICache.scala 51:22]
  reg  valid_386; // @[ICache.scala 51:22]
  reg  valid_387; // @[ICache.scala 51:22]
  reg  valid_388; // @[ICache.scala 51:22]
  reg  valid_389; // @[ICache.scala 51:22]
  reg  valid_390; // @[ICache.scala 51:22]
  reg  valid_391; // @[ICache.scala 51:22]
  reg  valid_392; // @[ICache.scala 51:22]
  reg  valid_393; // @[ICache.scala 51:22]
  reg  valid_394; // @[ICache.scala 51:22]
  reg  valid_395; // @[ICache.scala 51:22]
  reg  valid_396; // @[ICache.scala 51:22]
  reg  valid_397; // @[ICache.scala 51:22]
  reg  valid_398; // @[ICache.scala 51:22]
  reg  valid_399; // @[ICache.scala 51:22]
  reg  valid_400; // @[ICache.scala 51:22]
  reg  valid_401; // @[ICache.scala 51:22]
  reg  valid_402; // @[ICache.scala 51:22]
  reg  valid_403; // @[ICache.scala 51:22]
  reg  valid_404; // @[ICache.scala 51:22]
  reg  valid_405; // @[ICache.scala 51:22]
  reg  valid_406; // @[ICache.scala 51:22]
  reg  valid_407; // @[ICache.scala 51:22]
  reg  valid_408; // @[ICache.scala 51:22]
  reg  valid_409; // @[ICache.scala 51:22]
  reg  valid_410; // @[ICache.scala 51:22]
  reg  valid_411; // @[ICache.scala 51:22]
  reg  valid_412; // @[ICache.scala 51:22]
  reg  valid_413; // @[ICache.scala 51:22]
  reg  valid_414; // @[ICache.scala 51:22]
  reg  valid_415; // @[ICache.scala 51:22]
  reg  valid_416; // @[ICache.scala 51:22]
  reg  valid_417; // @[ICache.scala 51:22]
  reg  valid_418; // @[ICache.scala 51:22]
  reg  valid_419; // @[ICache.scala 51:22]
  reg  valid_420; // @[ICache.scala 51:22]
  reg  valid_421; // @[ICache.scala 51:22]
  reg  valid_422; // @[ICache.scala 51:22]
  reg  valid_423; // @[ICache.scala 51:22]
  reg  valid_424; // @[ICache.scala 51:22]
  reg  valid_425; // @[ICache.scala 51:22]
  reg  valid_426; // @[ICache.scala 51:22]
  reg  valid_427; // @[ICache.scala 51:22]
  reg  valid_428; // @[ICache.scala 51:22]
  reg  valid_429; // @[ICache.scala 51:22]
  reg  valid_430; // @[ICache.scala 51:22]
  reg  valid_431; // @[ICache.scala 51:22]
  reg  valid_432; // @[ICache.scala 51:22]
  reg  valid_433; // @[ICache.scala 51:22]
  reg  valid_434; // @[ICache.scala 51:22]
  reg  valid_435; // @[ICache.scala 51:22]
  reg  valid_436; // @[ICache.scala 51:22]
  reg  valid_437; // @[ICache.scala 51:22]
  reg  valid_438; // @[ICache.scala 51:22]
  reg  valid_439; // @[ICache.scala 51:22]
  reg  valid_440; // @[ICache.scala 51:22]
  reg  valid_441; // @[ICache.scala 51:22]
  reg  valid_442; // @[ICache.scala 51:22]
  reg  valid_443; // @[ICache.scala 51:22]
  reg  valid_444; // @[ICache.scala 51:22]
  reg  valid_445; // @[ICache.scala 51:22]
  reg  valid_446; // @[ICache.scala 51:22]
  reg  valid_447; // @[ICache.scala 51:22]
  reg  valid_448; // @[ICache.scala 51:22]
  reg  valid_449; // @[ICache.scala 51:22]
  reg  valid_450; // @[ICache.scala 51:22]
  reg  valid_451; // @[ICache.scala 51:22]
  reg  valid_452; // @[ICache.scala 51:22]
  reg  valid_453; // @[ICache.scala 51:22]
  reg  valid_454; // @[ICache.scala 51:22]
  reg  valid_455; // @[ICache.scala 51:22]
  reg  valid_456; // @[ICache.scala 51:22]
  reg  valid_457; // @[ICache.scala 51:22]
  reg  valid_458; // @[ICache.scala 51:22]
  reg  valid_459; // @[ICache.scala 51:22]
  reg  valid_460; // @[ICache.scala 51:22]
  reg  valid_461; // @[ICache.scala 51:22]
  reg  valid_462; // @[ICache.scala 51:22]
  reg  valid_463; // @[ICache.scala 51:22]
  reg  valid_464; // @[ICache.scala 51:22]
  reg  valid_465; // @[ICache.scala 51:22]
  reg  valid_466; // @[ICache.scala 51:22]
  reg  valid_467; // @[ICache.scala 51:22]
  reg  valid_468; // @[ICache.scala 51:22]
  reg  valid_469; // @[ICache.scala 51:22]
  reg  valid_470; // @[ICache.scala 51:22]
  reg  valid_471; // @[ICache.scala 51:22]
  reg  valid_472; // @[ICache.scala 51:22]
  reg  valid_473; // @[ICache.scala 51:22]
  reg  valid_474; // @[ICache.scala 51:22]
  reg  valid_475; // @[ICache.scala 51:22]
  reg  valid_476; // @[ICache.scala 51:22]
  reg  valid_477; // @[ICache.scala 51:22]
  reg  valid_478; // @[ICache.scala 51:22]
  reg  valid_479; // @[ICache.scala 51:22]
  reg  valid_480; // @[ICache.scala 51:22]
  reg  valid_481; // @[ICache.scala 51:22]
  reg  valid_482; // @[ICache.scala 51:22]
  reg  valid_483; // @[ICache.scala 51:22]
  reg  valid_484; // @[ICache.scala 51:22]
  reg  valid_485; // @[ICache.scala 51:22]
  reg  valid_486; // @[ICache.scala 51:22]
  reg  valid_487; // @[ICache.scala 51:22]
  reg  valid_488; // @[ICache.scala 51:22]
  reg  valid_489; // @[ICache.scala 51:22]
  reg  valid_490; // @[ICache.scala 51:22]
  reg  valid_491; // @[ICache.scala 51:22]
  reg  valid_492; // @[ICache.scala 51:22]
  reg  valid_493; // @[ICache.scala 51:22]
  reg  valid_494; // @[ICache.scala 51:22]
  reg  valid_495; // @[ICache.scala 51:22]
  reg  valid_496; // @[ICache.scala 51:22]
  reg  valid_497; // @[ICache.scala 51:22]
  reg  valid_498; // @[ICache.scala 51:22]
  reg  valid_499; // @[ICache.scala 51:22]
  reg  valid_500; // @[ICache.scala 51:22]
  reg  valid_501; // @[ICache.scala 51:22]
  reg  valid_502; // @[ICache.scala 51:22]
  reg  valid_503; // @[ICache.scala 51:22]
  reg  valid_504; // @[ICache.scala 51:22]
  reg  valid_505; // @[ICache.scala 51:22]
  reg  valid_506; // @[ICache.scala 51:22]
  reg  valid_507; // @[ICache.scala 51:22]
  reg  valid_508; // @[ICache.scala 51:22]
  reg  valid_509; // @[ICache.scala 51:22]
  reg  valid_510; // @[ICache.scala 51:22]
  reg  valid_511; // @[ICache.scala 51:22]
  reg  valid_512; // @[ICache.scala 51:22]
  reg  valid_513; // @[ICache.scala 51:22]
  reg  valid_514; // @[ICache.scala 51:22]
  reg  valid_515; // @[ICache.scala 51:22]
  reg  valid_516; // @[ICache.scala 51:22]
  reg  valid_517; // @[ICache.scala 51:22]
  reg  valid_518; // @[ICache.scala 51:22]
  reg  valid_519; // @[ICache.scala 51:22]
  reg  valid_520; // @[ICache.scala 51:22]
  reg  valid_521; // @[ICache.scala 51:22]
  reg  valid_522; // @[ICache.scala 51:22]
  reg  valid_523; // @[ICache.scala 51:22]
  reg  valid_524; // @[ICache.scala 51:22]
  reg  valid_525; // @[ICache.scala 51:22]
  reg  valid_526; // @[ICache.scala 51:22]
  reg  valid_527; // @[ICache.scala 51:22]
  reg  valid_528; // @[ICache.scala 51:22]
  reg  valid_529; // @[ICache.scala 51:22]
  reg  valid_530; // @[ICache.scala 51:22]
  reg  valid_531; // @[ICache.scala 51:22]
  reg  valid_532; // @[ICache.scala 51:22]
  reg  valid_533; // @[ICache.scala 51:22]
  reg  valid_534; // @[ICache.scala 51:22]
  reg  valid_535; // @[ICache.scala 51:22]
  reg  valid_536; // @[ICache.scala 51:22]
  reg  valid_537; // @[ICache.scala 51:22]
  reg  valid_538; // @[ICache.scala 51:22]
  reg  valid_539; // @[ICache.scala 51:22]
  reg  valid_540; // @[ICache.scala 51:22]
  reg  valid_541; // @[ICache.scala 51:22]
  reg  valid_542; // @[ICache.scala 51:22]
  reg  valid_543; // @[ICache.scala 51:22]
  reg  valid_544; // @[ICache.scala 51:22]
  reg  valid_545; // @[ICache.scala 51:22]
  reg  valid_546; // @[ICache.scala 51:22]
  reg  valid_547; // @[ICache.scala 51:22]
  reg  valid_548; // @[ICache.scala 51:22]
  reg  valid_549; // @[ICache.scala 51:22]
  reg  valid_550; // @[ICache.scala 51:22]
  reg  valid_551; // @[ICache.scala 51:22]
  reg  valid_552; // @[ICache.scala 51:22]
  reg  valid_553; // @[ICache.scala 51:22]
  reg  valid_554; // @[ICache.scala 51:22]
  reg  valid_555; // @[ICache.scala 51:22]
  reg  valid_556; // @[ICache.scala 51:22]
  reg  valid_557; // @[ICache.scala 51:22]
  reg  valid_558; // @[ICache.scala 51:22]
  reg  valid_559; // @[ICache.scala 51:22]
  reg  valid_560; // @[ICache.scala 51:22]
  reg  valid_561; // @[ICache.scala 51:22]
  reg  valid_562; // @[ICache.scala 51:22]
  reg  valid_563; // @[ICache.scala 51:22]
  reg  valid_564; // @[ICache.scala 51:22]
  reg  valid_565; // @[ICache.scala 51:22]
  reg  valid_566; // @[ICache.scala 51:22]
  reg  valid_567; // @[ICache.scala 51:22]
  reg  valid_568; // @[ICache.scala 51:22]
  reg  valid_569; // @[ICache.scala 51:22]
  reg  valid_570; // @[ICache.scala 51:22]
  reg  valid_571; // @[ICache.scala 51:22]
  reg  valid_572; // @[ICache.scala 51:22]
  reg  valid_573; // @[ICache.scala 51:22]
  reg  valid_574; // @[ICache.scala 51:22]
  reg  valid_575; // @[ICache.scala 51:22]
  reg  valid_576; // @[ICache.scala 51:22]
  reg  valid_577; // @[ICache.scala 51:22]
  reg  valid_578; // @[ICache.scala 51:22]
  reg  valid_579; // @[ICache.scala 51:22]
  reg  valid_580; // @[ICache.scala 51:22]
  reg  valid_581; // @[ICache.scala 51:22]
  reg  valid_582; // @[ICache.scala 51:22]
  reg  valid_583; // @[ICache.scala 51:22]
  reg  valid_584; // @[ICache.scala 51:22]
  reg  valid_585; // @[ICache.scala 51:22]
  reg  valid_586; // @[ICache.scala 51:22]
  reg  valid_587; // @[ICache.scala 51:22]
  reg  valid_588; // @[ICache.scala 51:22]
  reg  valid_589; // @[ICache.scala 51:22]
  reg  valid_590; // @[ICache.scala 51:22]
  reg  valid_591; // @[ICache.scala 51:22]
  reg  valid_592; // @[ICache.scala 51:22]
  reg  valid_593; // @[ICache.scala 51:22]
  reg  valid_594; // @[ICache.scala 51:22]
  reg  valid_595; // @[ICache.scala 51:22]
  reg  valid_596; // @[ICache.scala 51:22]
  reg  valid_597; // @[ICache.scala 51:22]
  reg  valid_598; // @[ICache.scala 51:22]
  reg  valid_599; // @[ICache.scala 51:22]
  reg  valid_600; // @[ICache.scala 51:22]
  reg  valid_601; // @[ICache.scala 51:22]
  reg  valid_602; // @[ICache.scala 51:22]
  reg  valid_603; // @[ICache.scala 51:22]
  reg  valid_604; // @[ICache.scala 51:22]
  reg  valid_605; // @[ICache.scala 51:22]
  reg  valid_606; // @[ICache.scala 51:22]
  reg  valid_607; // @[ICache.scala 51:22]
  reg  valid_608; // @[ICache.scala 51:22]
  reg  valid_609; // @[ICache.scala 51:22]
  reg  valid_610; // @[ICache.scala 51:22]
  reg  valid_611; // @[ICache.scala 51:22]
  reg  valid_612; // @[ICache.scala 51:22]
  reg  valid_613; // @[ICache.scala 51:22]
  reg  valid_614; // @[ICache.scala 51:22]
  reg  valid_615; // @[ICache.scala 51:22]
  reg  valid_616; // @[ICache.scala 51:22]
  reg  valid_617; // @[ICache.scala 51:22]
  reg  valid_618; // @[ICache.scala 51:22]
  reg  valid_619; // @[ICache.scala 51:22]
  reg  valid_620; // @[ICache.scala 51:22]
  reg  valid_621; // @[ICache.scala 51:22]
  reg  valid_622; // @[ICache.scala 51:22]
  reg  valid_623; // @[ICache.scala 51:22]
  reg  valid_624; // @[ICache.scala 51:22]
  reg  valid_625; // @[ICache.scala 51:22]
  reg  valid_626; // @[ICache.scala 51:22]
  reg  valid_627; // @[ICache.scala 51:22]
  reg  valid_628; // @[ICache.scala 51:22]
  reg  valid_629; // @[ICache.scala 51:22]
  reg  valid_630; // @[ICache.scala 51:22]
  reg  valid_631; // @[ICache.scala 51:22]
  reg  valid_632; // @[ICache.scala 51:22]
  reg  valid_633; // @[ICache.scala 51:22]
  reg  valid_634; // @[ICache.scala 51:22]
  reg  valid_635; // @[ICache.scala 51:22]
  reg  valid_636; // @[ICache.scala 51:22]
  reg  valid_637; // @[ICache.scala 51:22]
  reg  valid_638; // @[ICache.scala 51:22]
  reg  valid_639; // @[ICache.scala 51:22]
  reg  valid_640; // @[ICache.scala 51:22]
  reg  valid_641; // @[ICache.scala 51:22]
  reg  valid_642; // @[ICache.scala 51:22]
  reg  valid_643; // @[ICache.scala 51:22]
  reg  valid_644; // @[ICache.scala 51:22]
  reg  valid_645; // @[ICache.scala 51:22]
  reg  valid_646; // @[ICache.scala 51:22]
  reg  valid_647; // @[ICache.scala 51:22]
  reg  valid_648; // @[ICache.scala 51:22]
  reg  valid_649; // @[ICache.scala 51:22]
  reg  valid_650; // @[ICache.scala 51:22]
  reg  valid_651; // @[ICache.scala 51:22]
  reg  valid_652; // @[ICache.scala 51:22]
  reg  valid_653; // @[ICache.scala 51:22]
  reg  valid_654; // @[ICache.scala 51:22]
  reg  valid_655; // @[ICache.scala 51:22]
  reg  valid_656; // @[ICache.scala 51:22]
  reg  valid_657; // @[ICache.scala 51:22]
  reg  valid_658; // @[ICache.scala 51:22]
  reg  valid_659; // @[ICache.scala 51:22]
  reg  valid_660; // @[ICache.scala 51:22]
  reg  valid_661; // @[ICache.scala 51:22]
  reg  valid_662; // @[ICache.scala 51:22]
  reg  valid_663; // @[ICache.scala 51:22]
  reg  valid_664; // @[ICache.scala 51:22]
  reg  valid_665; // @[ICache.scala 51:22]
  reg  valid_666; // @[ICache.scala 51:22]
  reg  valid_667; // @[ICache.scala 51:22]
  reg  valid_668; // @[ICache.scala 51:22]
  reg  valid_669; // @[ICache.scala 51:22]
  reg  valid_670; // @[ICache.scala 51:22]
  reg  valid_671; // @[ICache.scala 51:22]
  reg  valid_672; // @[ICache.scala 51:22]
  reg  valid_673; // @[ICache.scala 51:22]
  reg  valid_674; // @[ICache.scala 51:22]
  reg  valid_675; // @[ICache.scala 51:22]
  reg  valid_676; // @[ICache.scala 51:22]
  reg  valid_677; // @[ICache.scala 51:22]
  reg  valid_678; // @[ICache.scala 51:22]
  reg  valid_679; // @[ICache.scala 51:22]
  reg  valid_680; // @[ICache.scala 51:22]
  reg  valid_681; // @[ICache.scala 51:22]
  reg  valid_682; // @[ICache.scala 51:22]
  reg  valid_683; // @[ICache.scala 51:22]
  reg  valid_684; // @[ICache.scala 51:22]
  reg  valid_685; // @[ICache.scala 51:22]
  reg  valid_686; // @[ICache.scala 51:22]
  reg  valid_687; // @[ICache.scala 51:22]
  reg  valid_688; // @[ICache.scala 51:22]
  reg  valid_689; // @[ICache.scala 51:22]
  reg  valid_690; // @[ICache.scala 51:22]
  reg  valid_691; // @[ICache.scala 51:22]
  reg  valid_692; // @[ICache.scala 51:22]
  reg  valid_693; // @[ICache.scala 51:22]
  reg  valid_694; // @[ICache.scala 51:22]
  reg  valid_695; // @[ICache.scala 51:22]
  reg  valid_696; // @[ICache.scala 51:22]
  reg  valid_697; // @[ICache.scala 51:22]
  reg  valid_698; // @[ICache.scala 51:22]
  reg  valid_699; // @[ICache.scala 51:22]
  reg  valid_700; // @[ICache.scala 51:22]
  reg  valid_701; // @[ICache.scala 51:22]
  reg  valid_702; // @[ICache.scala 51:22]
  reg  valid_703; // @[ICache.scala 51:22]
  reg  valid_704; // @[ICache.scala 51:22]
  reg  valid_705; // @[ICache.scala 51:22]
  reg  valid_706; // @[ICache.scala 51:22]
  reg  valid_707; // @[ICache.scala 51:22]
  reg  valid_708; // @[ICache.scala 51:22]
  reg  valid_709; // @[ICache.scala 51:22]
  reg  valid_710; // @[ICache.scala 51:22]
  reg  valid_711; // @[ICache.scala 51:22]
  reg  valid_712; // @[ICache.scala 51:22]
  reg  valid_713; // @[ICache.scala 51:22]
  reg  valid_714; // @[ICache.scala 51:22]
  reg  valid_715; // @[ICache.scala 51:22]
  reg  valid_716; // @[ICache.scala 51:22]
  reg  valid_717; // @[ICache.scala 51:22]
  reg  valid_718; // @[ICache.scala 51:22]
  reg  valid_719; // @[ICache.scala 51:22]
  reg  valid_720; // @[ICache.scala 51:22]
  reg  valid_721; // @[ICache.scala 51:22]
  reg  valid_722; // @[ICache.scala 51:22]
  reg  valid_723; // @[ICache.scala 51:22]
  reg  valid_724; // @[ICache.scala 51:22]
  reg  valid_725; // @[ICache.scala 51:22]
  reg  valid_726; // @[ICache.scala 51:22]
  reg  valid_727; // @[ICache.scala 51:22]
  reg  valid_728; // @[ICache.scala 51:22]
  reg  valid_729; // @[ICache.scala 51:22]
  reg  valid_730; // @[ICache.scala 51:22]
  reg  valid_731; // @[ICache.scala 51:22]
  reg  valid_732; // @[ICache.scala 51:22]
  reg  valid_733; // @[ICache.scala 51:22]
  reg  valid_734; // @[ICache.scala 51:22]
  reg  valid_735; // @[ICache.scala 51:22]
  reg  valid_736; // @[ICache.scala 51:22]
  reg  valid_737; // @[ICache.scala 51:22]
  reg  valid_738; // @[ICache.scala 51:22]
  reg  valid_739; // @[ICache.scala 51:22]
  reg  valid_740; // @[ICache.scala 51:22]
  reg  valid_741; // @[ICache.scala 51:22]
  reg  valid_742; // @[ICache.scala 51:22]
  reg  valid_743; // @[ICache.scala 51:22]
  reg  valid_744; // @[ICache.scala 51:22]
  reg  valid_745; // @[ICache.scala 51:22]
  reg  valid_746; // @[ICache.scala 51:22]
  reg  valid_747; // @[ICache.scala 51:22]
  reg  valid_748; // @[ICache.scala 51:22]
  reg  valid_749; // @[ICache.scala 51:22]
  reg  valid_750; // @[ICache.scala 51:22]
  reg  valid_751; // @[ICache.scala 51:22]
  reg  valid_752; // @[ICache.scala 51:22]
  reg  valid_753; // @[ICache.scala 51:22]
  reg  valid_754; // @[ICache.scala 51:22]
  reg  valid_755; // @[ICache.scala 51:22]
  reg  valid_756; // @[ICache.scala 51:22]
  reg  valid_757; // @[ICache.scala 51:22]
  reg  valid_758; // @[ICache.scala 51:22]
  reg  valid_759; // @[ICache.scala 51:22]
  reg  valid_760; // @[ICache.scala 51:22]
  reg  valid_761; // @[ICache.scala 51:22]
  reg  valid_762; // @[ICache.scala 51:22]
  reg  valid_763; // @[ICache.scala 51:22]
  reg  valid_764; // @[ICache.scala 51:22]
  reg  valid_765; // @[ICache.scala 51:22]
  reg  valid_766; // @[ICache.scala 51:22]
  reg  valid_767; // @[ICache.scala 51:22]
  reg  valid_768; // @[ICache.scala 51:22]
  reg  valid_769; // @[ICache.scala 51:22]
  reg  valid_770; // @[ICache.scala 51:22]
  reg  valid_771; // @[ICache.scala 51:22]
  reg  valid_772; // @[ICache.scala 51:22]
  reg  valid_773; // @[ICache.scala 51:22]
  reg  valid_774; // @[ICache.scala 51:22]
  reg  valid_775; // @[ICache.scala 51:22]
  reg  valid_776; // @[ICache.scala 51:22]
  reg  valid_777; // @[ICache.scala 51:22]
  reg  valid_778; // @[ICache.scala 51:22]
  reg  valid_779; // @[ICache.scala 51:22]
  reg  valid_780; // @[ICache.scala 51:22]
  reg  valid_781; // @[ICache.scala 51:22]
  reg  valid_782; // @[ICache.scala 51:22]
  reg  valid_783; // @[ICache.scala 51:22]
  reg  valid_784; // @[ICache.scala 51:22]
  reg  valid_785; // @[ICache.scala 51:22]
  reg  valid_786; // @[ICache.scala 51:22]
  reg  valid_787; // @[ICache.scala 51:22]
  reg  valid_788; // @[ICache.scala 51:22]
  reg  valid_789; // @[ICache.scala 51:22]
  reg  valid_790; // @[ICache.scala 51:22]
  reg  valid_791; // @[ICache.scala 51:22]
  reg  valid_792; // @[ICache.scala 51:22]
  reg  valid_793; // @[ICache.scala 51:22]
  reg  valid_794; // @[ICache.scala 51:22]
  reg  valid_795; // @[ICache.scala 51:22]
  reg  valid_796; // @[ICache.scala 51:22]
  reg  valid_797; // @[ICache.scala 51:22]
  reg  valid_798; // @[ICache.scala 51:22]
  reg  valid_799; // @[ICache.scala 51:22]
  reg  valid_800; // @[ICache.scala 51:22]
  reg  valid_801; // @[ICache.scala 51:22]
  reg  valid_802; // @[ICache.scala 51:22]
  reg  valid_803; // @[ICache.scala 51:22]
  reg  valid_804; // @[ICache.scala 51:22]
  reg  valid_805; // @[ICache.scala 51:22]
  reg  valid_806; // @[ICache.scala 51:22]
  reg  valid_807; // @[ICache.scala 51:22]
  reg  valid_808; // @[ICache.scala 51:22]
  reg  valid_809; // @[ICache.scala 51:22]
  reg  valid_810; // @[ICache.scala 51:22]
  reg  valid_811; // @[ICache.scala 51:22]
  reg  valid_812; // @[ICache.scala 51:22]
  reg  valid_813; // @[ICache.scala 51:22]
  reg  valid_814; // @[ICache.scala 51:22]
  reg  valid_815; // @[ICache.scala 51:22]
  reg  valid_816; // @[ICache.scala 51:22]
  reg  valid_817; // @[ICache.scala 51:22]
  reg  valid_818; // @[ICache.scala 51:22]
  reg  valid_819; // @[ICache.scala 51:22]
  reg  valid_820; // @[ICache.scala 51:22]
  reg  valid_821; // @[ICache.scala 51:22]
  reg  valid_822; // @[ICache.scala 51:22]
  reg  valid_823; // @[ICache.scala 51:22]
  reg  valid_824; // @[ICache.scala 51:22]
  reg  valid_825; // @[ICache.scala 51:22]
  reg  valid_826; // @[ICache.scala 51:22]
  reg  valid_827; // @[ICache.scala 51:22]
  reg  valid_828; // @[ICache.scala 51:22]
  reg  valid_829; // @[ICache.scala 51:22]
  reg  valid_830; // @[ICache.scala 51:22]
  reg  valid_831; // @[ICache.scala 51:22]
  reg  valid_832; // @[ICache.scala 51:22]
  reg  valid_833; // @[ICache.scala 51:22]
  reg  valid_834; // @[ICache.scala 51:22]
  reg  valid_835; // @[ICache.scala 51:22]
  reg  valid_836; // @[ICache.scala 51:22]
  reg  valid_837; // @[ICache.scala 51:22]
  reg  valid_838; // @[ICache.scala 51:22]
  reg  valid_839; // @[ICache.scala 51:22]
  reg  valid_840; // @[ICache.scala 51:22]
  reg  valid_841; // @[ICache.scala 51:22]
  reg  valid_842; // @[ICache.scala 51:22]
  reg  valid_843; // @[ICache.scala 51:22]
  reg  valid_844; // @[ICache.scala 51:22]
  reg  valid_845; // @[ICache.scala 51:22]
  reg  valid_846; // @[ICache.scala 51:22]
  reg  valid_847; // @[ICache.scala 51:22]
  reg  valid_848; // @[ICache.scala 51:22]
  reg  valid_849; // @[ICache.scala 51:22]
  reg  valid_850; // @[ICache.scala 51:22]
  reg  valid_851; // @[ICache.scala 51:22]
  reg  valid_852; // @[ICache.scala 51:22]
  reg  valid_853; // @[ICache.scala 51:22]
  reg  valid_854; // @[ICache.scala 51:22]
  reg  valid_855; // @[ICache.scala 51:22]
  reg  valid_856; // @[ICache.scala 51:22]
  reg  valid_857; // @[ICache.scala 51:22]
  reg  valid_858; // @[ICache.scala 51:22]
  reg  valid_859; // @[ICache.scala 51:22]
  reg  valid_860; // @[ICache.scala 51:22]
  reg  valid_861; // @[ICache.scala 51:22]
  reg  valid_862; // @[ICache.scala 51:22]
  reg  valid_863; // @[ICache.scala 51:22]
  reg  valid_864; // @[ICache.scala 51:22]
  reg  valid_865; // @[ICache.scala 51:22]
  reg  valid_866; // @[ICache.scala 51:22]
  reg  valid_867; // @[ICache.scala 51:22]
  reg  valid_868; // @[ICache.scala 51:22]
  reg  valid_869; // @[ICache.scala 51:22]
  reg  valid_870; // @[ICache.scala 51:22]
  reg  valid_871; // @[ICache.scala 51:22]
  reg  valid_872; // @[ICache.scala 51:22]
  reg  valid_873; // @[ICache.scala 51:22]
  reg  valid_874; // @[ICache.scala 51:22]
  reg  valid_875; // @[ICache.scala 51:22]
  reg  valid_876; // @[ICache.scala 51:22]
  reg  valid_877; // @[ICache.scala 51:22]
  reg  valid_878; // @[ICache.scala 51:22]
  reg  valid_879; // @[ICache.scala 51:22]
  reg  valid_880; // @[ICache.scala 51:22]
  reg  valid_881; // @[ICache.scala 51:22]
  reg  valid_882; // @[ICache.scala 51:22]
  reg  valid_883; // @[ICache.scala 51:22]
  reg  valid_884; // @[ICache.scala 51:22]
  reg  valid_885; // @[ICache.scala 51:22]
  reg  valid_886; // @[ICache.scala 51:22]
  reg  valid_887; // @[ICache.scala 51:22]
  reg  valid_888; // @[ICache.scala 51:22]
  reg  valid_889; // @[ICache.scala 51:22]
  reg  valid_890; // @[ICache.scala 51:22]
  reg  valid_891; // @[ICache.scala 51:22]
  reg  valid_892; // @[ICache.scala 51:22]
  reg  valid_893; // @[ICache.scala 51:22]
  reg  valid_894; // @[ICache.scala 51:22]
  reg  valid_895; // @[ICache.scala 51:22]
  reg  valid_896; // @[ICache.scala 51:22]
  reg  valid_897; // @[ICache.scala 51:22]
  reg  valid_898; // @[ICache.scala 51:22]
  reg  valid_899; // @[ICache.scala 51:22]
  reg  valid_900; // @[ICache.scala 51:22]
  reg  valid_901; // @[ICache.scala 51:22]
  reg  valid_902; // @[ICache.scala 51:22]
  reg  valid_903; // @[ICache.scala 51:22]
  reg  valid_904; // @[ICache.scala 51:22]
  reg  valid_905; // @[ICache.scala 51:22]
  reg  valid_906; // @[ICache.scala 51:22]
  reg  valid_907; // @[ICache.scala 51:22]
  reg  valid_908; // @[ICache.scala 51:22]
  reg  valid_909; // @[ICache.scala 51:22]
  reg  valid_910; // @[ICache.scala 51:22]
  reg  valid_911; // @[ICache.scala 51:22]
  reg  valid_912; // @[ICache.scala 51:22]
  reg  valid_913; // @[ICache.scala 51:22]
  reg  valid_914; // @[ICache.scala 51:22]
  reg  valid_915; // @[ICache.scala 51:22]
  reg  valid_916; // @[ICache.scala 51:22]
  reg  valid_917; // @[ICache.scala 51:22]
  reg  valid_918; // @[ICache.scala 51:22]
  reg  valid_919; // @[ICache.scala 51:22]
  reg  valid_920; // @[ICache.scala 51:22]
  reg  valid_921; // @[ICache.scala 51:22]
  reg  valid_922; // @[ICache.scala 51:22]
  reg  valid_923; // @[ICache.scala 51:22]
  reg  valid_924; // @[ICache.scala 51:22]
  reg  valid_925; // @[ICache.scala 51:22]
  reg  valid_926; // @[ICache.scala 51:22]
  reg  valid_927; // @[ICache.scala 51:22]
  reg  valid_928; // @[ICache.scala 51:22]
  reg  valid_929; // @[ICache.scala 51:22]
  reg  valid_930; // @[ICache.scala 51:22]
  reg  valid_931; // @[ICache.scala 51:22]
  reg  valid_932; // @[ICache.scala 51:22]
  reg  valid_933; // @[ICache.scala 51:22]
  reg  valid_934; // @[ICache.scala 51:22]
  reg  valid_935; // @[ICache.scala 51:22]
  reg  valid_936; // @[ICache.scala 51:22]
  reg  valid_937; // @[ICache.scala 51:22]
  reg  valid_938; // @[ICache.scala 51:22]
  reg  valid_939; // @[ICache.scala 51:22]
  reg  valid_940; // @[ICache.scala 51:22]
  reg  valid_941; // @[ICache.scala 51:22]
  reg  valid_942; // @[ICache.scala 51:22]
  reg  valid_943; // @[ICache.scala 51:22]
  reg  valid_944; // @[ICache.scala 51:22]
  reg  valid_945; // @[ICache.scala 51:22]
  reg  valid_946; // @[ICache.scala 51:22]
  reg  valid_947; // @[ICache.scala 51:22]
  reg  valid_948; // @[ICache.scala 51:22]
  reg  valid_949; // @[ICache.scala 51:22]
  reg  valid_950; // @[ICache.scala 51:22]
  reg  valid_951; // @[ICache.scala 51:22]
  reg  valid_952; // @[ICache.scala 51:22]
  reg  valid_953; // @[ICache.scala 51:22]
  reg  valid_954; // @[ICache.scala 51:22]
  reg  valid_955; // @[ICache.scala 51:22]
  reg  valid_956; // @[ICache.scala 51:22]
  reg  valid_957; // @[ICache.scala 51:22]
  reg  valid_958; // @[ICache.scala 51:22]
  reg  valid_959; // @[ICache.scala 51:22]
  reg  valid_960; // @[ICache.scala 51:22]
  reg  valid_961; // @[ICache.scala 51:22]
  reg  valid_962; // @[ICache.scala 51:22]
  reg  valid_963; // @[ICache.scala 51:22]
  reg  valid_964; // @[ICache.scala 51:22]
  reg  valid_965; // @[ICache.scala 51:22]
  reg  valid_966; // @[ICache.scala 51:22]
  reg  valid_967; // @[ICache.scala 51:22]
  reg  valid_968; // @[ICache.scala 51:22]
  reg  valid_969; // @[ICache.scala 51:22]
  reg  valid_970; // @[ICache.scala 51:22]
  reg  valid_971; // @[ICache.scala 51:22]
  reg  valid_972; // @[ICache.scala 51:22]
  reg  valid_973; // @[ICache.scala 51:22]
  reg  valid_974; // @[ICache.scala 51:22]
  reg  valid_975; // @[ICache.scala 51:22]
  reg  valid_976; // @[ICache.scala 51:22]
  reg  valid_977; // @[ICache.scala 51:22]
  reg  valid_978; // @[ICache.scala 51:22]
  reg  valid_979; // @[ICache.scala 51:22]
  reg  valid_980; // @[ICache.scala 51:22]
  reg  valid_981; // @[ICache.scala 51:22]
  reg  valid_982; // @[ICache.scala 51:22]
  reg  valid_983; // @[ICache.scala 51:22]
  reg  valid_984; // @[ICache.scala 51:22]
  reg  valid_985; // @[ICache.scala 51:22]
  reg  valid_986; // @[ICache.scala 51:22]
  reg  valid_987; // @[ICache.scala 51:22]
  reg  valid_988; // @[ICache.scala 51:22]
  reg  valid_989; // @[ICache.scala 51:22]
  reg  valid_990; // @[ICache.scala 51:22]
  reg  valid_991; // @[ICache.scala 51:22]
  reg  valid_992; // @[ICache.scala 51:22]
  reg  valid_993; // @[ICache.scala 51:22]
  reg  valid_994; // @[ICache.scala 51:22]
  reg  valid_995; // @[ICache.scala 51:22]
  reg  valid_996; // @[ICache.scala 51:22]
  reg  valid_997; // @[ICache.scala 51:22]
  reg  valid_998; // @[ICache.scala 51:22]
  reg  valid_999; // @[ICache.scala 51:22]
  reg  valid_1000; // @[ICache.scala 51:22]
  reg  valid_1001; // @[ICache.scala 51:22]
  reg  valid_1002; // @[ICache.scala 51:22]
  reg  valid_1003; // @[ICache.scala 51:22]
  reg  valid_1004; // @[ICache.scala 51:22]
  reg  valid_1005; // @[ICache.scala 51:22]
  reg  valid_1006; // @[ICache.scala 51:22]
  reg  valid_1007; // @[ICache.scala 51:22]
  reg  valid_1008; // @[ICache.scala 51:22]
  reg  valid_1009; // @[ICache.scala 51:22]
  reg  valid_1010; // @[ICache.scala 51:22]
  reg  valid_1011; // @[ICache.scala 51:22]
  reg  valid_1012; // @[ICache.scala 51:22]
  reg  valid_1013; // @[ICache.scala 51:22]
  reg  valid_1014; // @[ICache.scala 51:22]
  reg  valid_1015; // @[ICache.scala 51:22]
  reg  valid_1016; // @[ICache.scala 51:22]
  reg  valid_1017; // @[ICache.scala 51:22]
  reg  valid_1018; // @[ICache.scala 51:22]
  reg  valid_1019; // @[ICache.scala 51:22]
  reg  valid_1020; // @[ICache.scala 51:22]
  reg  valid_1021; // @[ICache.scala 51:22]
  reg  valid_1022; // @[ICache.scala 51:22]
  reg  valid_1023; // @[ICache.scala 51:22]
  reg [2:0] state; // @[ICache.scala 78:68]
  wire  _GEN_2 = 10'h1 == req_r_addr[14:5] ? valid_1 : valid_0; // @[ICache.scala 68:{44,44}]
  wire  _GEN_3 = 10'h2 == req_r_addr[14:5] ? valid_2 : _GEN_2; // @[ICache.scala 68:{44,44}]
  wire  _GEN_4 = 10'h3 == req_r_addr[14:5] ? valid_3 : _GEN_3; // @[ICache.scala 68:{44,44}]
  wire  _GEN_5 = 10'h4 == req_r_addr[14:5] ? valid_4 : _GEN_4; // @[ICache.scala 68:{44,44}]
  wire  _GEN_6 = 10'h5 == req_r_addr[14:5] ? valid_5 : _GEN_5; // @[ICache.scala 68:{44,44}]
  wire  _GEN_7 = 10'h6 == req_r_addr[14:5] ? valid_6 : _GEN_6; // @[ICache.scala 68:{44,44}]
  wire  _GEN_8 = 10'h7 == req_r_addr[14:5] ? valid_7 : _GEN_7; // @[ICache.scala 68:{44,44}]
  wire  _GEN_9 = 10'h8 == req_r_addr[14:5] ? valid_8 : _GEN_8; // @[ICache.scala 68:{44,44}]
  wire  _GEN_10 = 10'h9 == req_r_addr[14:5] ? valid_9 : _GEN_9; // @[ICache.scala 68:{44,44}]
  wire  _GEN_11 = 10'ha == req_r_addr[14:5] ? valid_10 : _GEN_10; // @[ICache.scala 68:{44,44}]
  wire  _GEN_12 = 10'hb == req_r_addr[14:5] ? valid_11 : _GEN_11; // @[ICache.scala 68:{44,44}]
  wire  _GEN_13 = 10'hc == req_r_addr[14:5] ? valid_12 : _GEN_12; // @[ICache.scala 68:{44,44}]
  wire  _GEN_14 = 10'hd == req_r_addr[14:5] ? valid_13 : _GEN_13; // @[ICache.scala 68:{44,44}]
  wire  _GEN_15 = 10'he == req_r_addr[14:5] ? valid_14 : _GEN_14; // @[ICache.scala 68:{44,44}]
  wire  _GEN_16 = 10'hf == req_r_addr[14:5] ? valid_15 : _GEN_15; // @[ICache.scala 68:{44,44}]
  wire  _GEN_17 = 10'h10 == req_r_addr[14:5] ? valid_16 : _GEN_16; // @[ICache.scala 68:{44,44}]
  wire  _GEN_18 = 10'h11 == req_r_addr[14:5] ? valid_17 : _GEN_17; // @[ICache.scala 68:{44,44}]
  wire  _GEN_19 = 10'h12 == req_r_addr[14:5] ? valid_18 : _GEN_18; // @[ICache.scala 68:{44,44}]
  wire  _GEN_20 = 10'h13 == req_r_addr[14:5] ? valid_19 : _GEN_19; // @[ICache.scala 68:{44,44}]
  wire  _GEN_21 = 10'h14 == req_r_addr[14:5] ? valid_20 : _GEN_20; // @[ICache.scala 68:{44,44}]
  wire  _GEN_22 = 10'h15 == req_r_addr[14:5] ? valid_21 : _GEN_21; // @[ICache.scala 68:{44,44}]
  wire  _GEN_23 = 10'h16 == req_r_addr[14:5] ? valid_22 : _GEN_22; // @[ICache.scala 68:{44,44}]
  wire  _GEN_24 = 10'h17 == req_r_addr[14:5] ? valid_23 : _GEN_23; // @[ICache.scala 68:{44,44}]
  wire  _GEN_25 = 10'h18 == req_r_addr[14:5] ? valid_24 : _GEN_24; // @[ICache.scala 68:{44,44}]
  wire  _GEN_26 = 10'h19 == req_r_addr[14:5] ? valid_25 : _GEN_25; // @[ICache.scala 68:{44,44}]
  wire  _GEN_27 = 10'h1a == req_r_addr[14:5] ? valid_26 : _GEN_26; // @[ICache.scala 68:{44,44}]
  wire  _GEN_28 = 10'h1b == req_r_addr[14:5] ? valid_27 : _GEN_27; // @[ICache.scala 68:{44,44}]
  wire  _GEN_29 = 10'h1c == req_r_addr[14:5] ? valid_28 : _GEN_28; // @[ICache.scala 68:{44,44}]
  wire  _GEN_30 = 10'h1d == req_r_addr[14:5] ? valid_29 : _GEN_29; // @[ICache.scala 68:{44,44}]
  wire  _GEN_31 = 10'h1e == req_r_addr[14:5] ? valid_30 : _GEN_30; // @[ICache.scala 68:{44,44}]
  wire  _GEN_32 = 10'h1f == req_r_addr[14:5] ? valid_31 : _GEN_31; // @[ICache.scala 68:{44,44}]
  wire  _GEN_33 = 10'h20 == req_r_addr[14:5] ? valid_32 : _GEN_32; // @[ICache.scala 68:{44,44}]
  wire  _GEN_34 = 10'h21 == req_r_addr[14:5] ? valid_33 : _GEN_33; // @[ICache.scala 68:{44,44}]
  wire  _GEN_35 = 10'h22 == req_r_addr[14:5] ? valid_34 : _GEN_34; // @[ICache.scala 68:{44,44}]
  wire  _GEN_36 = 10'h23 == req_r_addr[14:5] ? valid_35 : _GEN_35; // @[ICache.scala 68:{44,44}]
  wire  _GEN_37 = 10'h24 == req_r_addr[14:5] ? valid_36 : _GEN_36; // @[ICache.scala 68:{44,44}]
  wire  _GEN_38 = 10'h25 == req_r_addr[14:5] ? valid_37 : _GEN_37; // @[ICache.scala 68:{44,44}]
  wire  _GEN_39 = 10'h26 == req_r_addr[14:5] ? valid_38 : _GEN_38; // @[ICache.scala 68:{44,44}]
  wire  _GEN_40 = 10'h27 == req_r_addr[14:5] ? valid_39 : _GEN_39; // @[ICache.scala 68:{44,44}]
  wire  _GEN_41 = 10'h28 == req_r_addr[14:5] ? valid_40 : _GEN_40; // @[ICache.scala 68:{44,44}]
  wire  _GEN_42 = 10'h29 == req_r_addr[14:5] ? valid_41 : _GEN_41; // @[ICache.scala 68:{44,44}]
  wire  _GEN_43 = 10'h2a == req_r_addr[14:5] ? valid_42 : _GEN_42; // @[ICache.scala 68:{44,44}]
  wire  _GEN_44 = 10'h2b == req_r_addr[14:5] ? valid_43 : _GEN_43; // @[ICache.scala 68:{44,44}]
  wire  _GEN_45 = 10'h2c == req_r_addr[14:5] ? valid_44 : _GEN_44; // @[ICache.scala 68:{44,44}]
  wire  _GEN_46 = 10'h2d == req_r_addr[14:5] ? valid_45 : _GEN_45; // @[ICache.scala 68:{44,44}]
  wire  _GEN_47 = 10'h2e == req_r_addr[14:5] ? valid_46 : _GEN_46; // @[ICache.scala 68:{44,44}]
  wire  _GEN_48 = 10'h2f == req_r_addr[14:5] ? valid_47 : _GEN_47; // @[ICache.scala 68:{44,44}]
  wire  _GEN_49 = 10'h30 == req_r_addr[14:5] ? valid_48 : _GEN_48; // @[ICache.scala 68:{44,44}]
  wire  _GEN_50 = 10'h31 == req_r_addr[14:5] ? valid_49 : _GEN_49; // @[ICache.scala 68:{44,44}]
  wire  _GEN_51 = 10'h32 == req_r_addr[14:5] ? valid_50 : _GEN_50; // @[ICache.scala 68:{44,44}]
  wire  _GEN_52 = 10'h33 == req_r_addr[14:5] ? valid_51 : _GEN_51; // @[ICache.scala 68:{44,44}]
  wire  _GEN_53 = 10'h34 == req_r_addr[14:5] ? valid_52 : _GEN_52; // @[ICache.scala 68:{44,44}]
  wire  _GEN_54 = 10'h35 == req_r_addr[14:5] ? valid_53 : _GEN_53; // @[ICache.scala 68:{44,44}]
  wire  _GEN_55 = 10'h36 == req_r_addr[14:5] ? valid_54 : _GEN_54; // @[ICache.scala 68:{44,44}]
  wire  _GEN_56 = 10'h37 == req_r_addr[14:5] ? valid_55 : _GEN_55; // @[ICache.scala 68:{44,44}]
  wire  _GEN_57 = 10'h38 == req_r_addr[14:5] ? valid_56 : _GEN_56; // @[ICache.scala 68:{44,44}]
  wire  _GEN_58 = 10'h39 == req_r_addr[14:5] ? valid_57 : _GEN_57; // @[ICache.scala 68:{44,44}]
  wire  _GEN_59 = 10'h3a == req_r_addr[14:5] ? valid_58 : _GEN_58; // @[ICache.scala 68:{44,44}]
  wire  _GEN_60 = 10'h3b == req_r_addr[14:5] ? valid_59 : _GEN_59; // @[ICache.scala 68:{44,44}]
  wire  _GEN_61 = 10'h3c == req_r_addr[14:5] ? valid_60 : _GEN_60; // @[ICache.scala 68:{44,44}]
  wire  _GEN_62 = 10'h3d == req_r_addr[14:5] ? valid_61 : _GEN_61; // @[ICache.scala 68:{44,44}]
  wire  _GEN_63 = 10'h3e == req_r_addr[14:5] ? valid_62 : _GEN_62; // @[ICache.scala 68:{44,44}]
  wire  _GEN_64 = 10'h3f == req_r_addr[14:5] ? valid_63 : _GEN_63; // @[ICache.scala 68:{44,44}]
  wire  _GEN_65 = 10'h40 == req_r_addr[14:5] ? valid_64 : _GEN_64; // @[ICache.scala 68:{44,44}]
  wire  _GEN_66 = 10'h41 == req_r_addr[14:5] ? valid_65 : _GEN_65; // @[ICache.scala 68:{44,44}]
  wire  _GEN_67 = 10'h42 == req_r_addr[14:5] ? valid_66 : _GEN_66; // @[ICache.scala 68:{44,44}]
  wire  _GEN_68 = 10'h43 == req_r_addr[14:5] ? valid_67 : _GEN_67; // @[ICache.scala 68:{44,44}]
  wire  _GEN_69 = 10'h44 == req_r_addr[14:5] ? valid_68 : _GEN_68; // @[ICache.scala 68:{44,44}]
  wire  _GEN_70 = 10'h45 == req_r_addr[14:5] ? valid_69 : _GEN_69; // @[ICache.scala 68:{44,44}]
  wire  _GEN_71 = 10'h46 == req_r_addr[14:5] ? valid_70 : _GEN_70; // @[ICache.scala 68:{44,44}]
  wire  _GEN_72 = 10'h47 == req_r_addr[14:5] ? valid_71 : _GEN_71; // @[ICache.scala 68:{44,44}]
  wire  _GEN_73 = 10'h48 == req_r_addr[14:5] ? valid_72 : _GEN_72; // @[ICache.scala 68:{44,44}]
  wire  _GEN_74 = 10'h49 == req_r_addr[14:5] ? valid_73 : _GEN_73; // @[ICache.scala 68:{44,44}]
  wire  _GEN_75 = 10'h4a == req_r_addr[14:5] ? valid_74 : _GEN_74; // @[ICache.scala 68:{44,44}]
  wire  _GEN_76 = 10'h4b == req_r_addr[14:5] ? valid_75 : _GEN_75; // @[ICache.scala 68:{44,44}]
  wire  _GEN_77 = 10'h4c == req_r_addr[14:5] ? valid_76 : _GEN_76; // @[ICache.scala 68:{44,44}]
  wire  _GEN_78 = 10'h4d == req_r_addr[14:5] ? valid_77 : _GEN_77; // @[ICache.scala 68:{44,44}]
  wire  _GEN_79 = 10'h4e == req_r_addr[14:5] ? valid_78 : _GEN_78; // @[ICache.scala 68:{44,44}]
  wire  _GEN_80 = 10'h4f == req_r_addr[14:5] ? valid_79 : _GEN_79; // @[ICache.scala 68:{44,44}]
  wire  _GEN_81 = 10'h50 == req_r_addr[14:5] ? valid_80 : _GEN_80; // @[ICache.scala 68:{44,44}]
  wire  _GEN_82 = 10'h51 == req_r_addr[14:5] ? valid_81 : _GEN_81; // @[ICache.scala 68:{44,44}]
  wire  _GEN_83 = 10'h52 == req_r_addr[14:5] ? valid_82 : _GEN_82; // @[ICache.scala 68:{44,44}]
  wire  _GEN_84 = 10'h53 == req_r_addr[14:5] ? valid_83 : _GEN_83; // @[ICache.scala 68:{44,44}]
  wire  _GEN_85 = 10'h54 == req_r_addr[14:5] ? valid_84 : _GEN_84; // @[ICache.scala 68:{44,44}]
  wire  _GEN_86 = 10'h55 == req_r_addr[14:5] ? valid_85 : _GEN_85; // @[ICache.scala 68:{44,44}]
  wire  _GEN_87 = 10'h56 == req_r_addr[14:5] ? valid_86 : _GEN_86; // @[ICache.scala 68:{44,44}]
  wire  _GEN_88 = 10'h57 == req_r_addr[14:5] ? valid_87 : _GEN_87; // @[ICache.scala 68:{44,44}]
  wire  _GEN_89 = 10'h58 == req_r_addr[14:5] ? valid_88 : _GEN_88; // @[ICache.scala 68:{44,44}]
  wire  _GEN_90 = 10'h59 == req_r_addr[14:5] ? valid_89 : _GEN_89; // @[ICache.scala 68:{44,44}]
  wire  _GEN_91 = 10'h5a == req_r_addr[14:5] ? valid_90 : _GEN_90; // @[ICache.scala 68:{44,44}]
  wire  _GEN_92 = 10'h5b == req_r_addr[14:5] ? valid_91 : _GEN_91; // @[ICache.scala 68:{44,44}]
  wire  _GEN_93 = 10'h5c == req_r_addr[14:5] ? valid_92 : _GEN_92; // @[ICache.scala 68:{44,44}]
  wire  _GEN_94 = 10'h5d == req_r_addr[14:5] ? valid_93 : _GEN_93; // @[ICache.scala 68:{44,44}]
  wire  _GEN_95 = 10'h5e == req_r_addr[14:5] ? valid_94 : _GEN_94; // @[ICache.scala 68:{44,44}]
  wire  _GEN_96 = 10'h5f == req_r_addr[14:5] ? valid_95 : _GEN_95; // @[ICache.scala 68:{44,44}]
  wire  _GEN_97 = 10'h60 == req_r_addr[14:5] ? valid_96 : _GEN_96; // @[ICache.scala 68:{44,44}]
  wire  _GEN_98 = 10'h61 == req_r_addr[14:5] ? valid_97 : _GEN_97; // @[ICache.scala 68:{44,44}]
  wire  _GEN_99 = 10'h62 == req_r_addr[14:5] ? valid_98 : _GEN_98; // @[ICache.scala 68:{44,44}]
  wire  _GEN_100 = 10'h63 == req_r_addr[14:5] ? valid_99 : _GEN_99; // @[ICache.scala 68:{44,44}]
  wire  _GEN_101 = 10'h64 == req_r_addr[14:5] ? valid_100 : _GEN_100; // @[ICache.scala 68:{44,44}]
  wire  _GEN_102 = 10'h65 == req_r_addr[14:5] ? valid_101 : _GEN_101; // @[ICache.scala 68:{44,44}]
  wire  _GEN_103 = 10'h66 == req_r_addr[14:5] ? valid_102 : _GEN_102; // @[ICache.scala 68:{44,44}]
  wire  _GEN_104 = 10'h67 == req_r_addr[14:5] ? valid_103 : _GEN_103; // @[ICache.scala 68:{44,44}]
  wire  _GEN_105 = 10'h68 == req_r_addr[14:5] ? valid_104 : _GEN_104; // @[ICache.scala 68:{44,44}]
  wire  _GEN_106 = 10'h69 == req_r_addr[14:5] ? valid_105 : _GEN_105; // @[ICache.scala 68:{44,44}]
  wire  _GEN_107 = 10'h6a == req_r_addr[14:5] ? valid_106 : _GEN_106; // @[ICache.scala 68:{44,44}]
  wire  _GEN_108 = 10'h6b == req_r_addr[14:5] ? valid_107 : _GEN_107; // @[ICache.scala 68:{44,44}]
  wire  _GEN_109 = 10'h6c == req_r_addr[14:5] ? valid_108 : _GEN_108; // @[ICache.scala 68:{44,44}]
  wire  _GEN_110 = 10'h6d == req_r_addr[14:5] ? valid_109 : _GEN_109; // @[ICache.scala 68:{44,44}]
  wire  _GEN_111 = 10'h6e == req_r_addr[14:5] ? valid_110 : _GEN_110; // @[ICache.scala 68:{44,44}]
  wire  _GEN_112 = 10'h6f == req_r_addr[14:5] ? valid_111 : _GEN_111; // @[ICache.scala 68:{44,44}]
  wire  _GEN_113 = 10'h70 == req_r_addr[14:5] ? valid_112 : _GEN_112; // @[ICache.scala 68:{44,44}]
  wire  _GEN_114 = 10'h71 == req_r_addr[14:5] ? valid_113 : _GEN_113; // @[ICache.scala 68:{44,44}]
  wire  _GEN_115 = 10'h72 == req_r_addr[14:5] ? valid_114 : _GEN_114; // @[ICache.scala 68:{44,44}]
  wire  _GEN_116 = 10'h73 == req_r_addr[14:5] ? valid_115 : _GEN_115; // @[ICache.scala 68:{44,44}]
  wire  _GEN_117 = 10'h74 == req_r_addr[14:5] ? valid_116 : _GEN_116; // @[ICache.scala 68:{44,44}]
  wire  _GEN_118 = 10'h75 == req_r_addr[14:5] ? valid_117 : _GEN_117; // @[ICache.scala 68:{44,44}]
  wire  _GEN_119 = 10'h76 == req_r_addr[14:5] ? valid_118 : _GEN_118; // @[ICache.scala 68:{44,44}]
  wire  _GEN_120 = 10'h77 == req_r_addr[14:5] ? valid_119 : _GEN_119; // @[ICache.scala 68:{44,44}]
  wire  _GEN_121 = 10'h78 == req_r_addr[14:5] ? valid_120 : _GEN_120; // @[ICache.scala 68:{44,44}]
  wire  _GEN_122 = 10'h79 == req_r_addr[14:5] ? valid_121 : _GEN_121; // @[ICache.scala 68:{44,44}]
  wire  _GEN_123 = 10'h7a == req_r_addr[14:5] ? valid_122 : _GEN_122; // @[ICache.scala 68:{44,44}]
  wire  _GEN_124 = 10'h7b == req_r_addr[14:5] ? valid_123 : _GEN_123; // @[ICache.scala 68:{44,44}]
  wire  _GEN_125 = 10'h7c == req_r_addr[14:5] ? valid_124 : _GEN_124; // @[ICache.scala 68:{44,44}]
  wire  _GEN_126 = 10'h7d == req_r_addr[14:5] ? valid_125 : _GEN_125; // @[ICache.scala 68:{44,44}]
  wire  _GEN_127 = 10'h7e == req_r_addr[14:5] ? valid_126 : _GEN_126; // @[ICache.scala 68:{44,44}]
  wire  _GEN_128 = 10'h7f == req_r_addr[14:5] ? valid_127 : _GEN_127; // @[ICache.scala 68:{44,44}]
  wire  _GEN_129 = 10'h80 == req_r_addr[14:5] ? valid_128 : _GEN_128; // @[ICache.scala 68:{44,44}]
  wire  _GEN_130 = 10'h81 == req_r_addr[14:5] ? valid_129 : _GEN_129; // @[ICache.scala 68:{44,44}]
  wire  _GEN_131 = 10'h82 == req_r_addr[14:5] ? valid_130 : _GEN_130; // @[ICache.scala 68:{44,44}]
  wire  _GEN_132 = 10'h83 == req_r_addr[14:5] ? valid_131 : _GEN_131; // @[ICache.scala 68:{44,44}]
  wire  _GEN_133 = 10'h84 == req_r_addr[14:5] ? valid_132 : _GEN_132; // @[ICache.scala 68:{44,44}]
  wire  _GEN_134 = 10'h85 == req_r_addr[14:5] ? valid_133 : _GEN_133; // @[ICache.scala 68:{44,44}]
  wire  _GEN_135 = 10'h86 == req_r_addr[14:5] ? valid_134 : _GEN_134; // @[ICache.scala 68:{44,44}]
  wire  _GEN_136 = 10'h87 == req_r_addr[14:5] ? valid_135 : _GEN_135; // @[ICache.scala 68:{44,44}]
  wire  _GEN_137 = 10'h88 == req_r_addr[14:5] ? valid_136 : _GEN_136; // @[ICache.scala 68:{44,44}]
  wire  _GEN_138 = 10'h89 == req_r_addr[14:5] ? valid_137 : _GEN_137; // @[ICache.scala 68:{44,44}]
  wire  _GEN_139 = 10'h8a == req_r_addr[14:5] ? valid_138 : _GEN_138; // @[ICache.scala 68:{44,44}]
  wire  _GEN_140 = 10'h8b == req_r_addr[14:5] ? valid_139 : _GEN_139; // @[ICache.scala 68:{44,44}]
  wire  _GEN_141 = 10'h8c == req_r_addr[14:5] ? valid_140 : _GEN_140; // @[ICache.scala 68:{44,44}]
  wire  _GEN_142 = 10'h8d == req_r_addr[14:5] ? valid_141 : _GEN_141; // @[ICache.scala 68:{44,44}]
  wire  _GEN_143 = 10'h8e == req_r_addr[14:5] ? valid_142 : _GEN_142; // @[ICache.scala 68:{44,44}]
  wire  _GEN_144 = 10'h8f == req_r_addr[14:5] ? valid_143 : _GEN_143; // @[ICache.scala 68:{44,44}]
  wire  _GEN_145 = 10'h90 == req_r_addr[14:5] ? valid_144 : _GEN_144; // @[ICache.scala 68:{44,44}]
  wire  _GEN_146 = 10'h91 == req_r_addr[14:5] ? valid_145 : _GEN_145; // @[ICache.scala 68:{44,44}]
  wire  _GEN_147 = 10'h92 == req_r_addr[14:5] ? valid_146 : _GEN_146; // @[ICache.scala 68:{44,44}]
  wire  _GEN_148 = 10'h93 == req_r_addr[14:5] ? valid_147 : _GEN_147; // @[ICache.scala 68:{44,44}]
  wire  _GEN_149 = 10'h94 == req_r_addr[14:5] ? valid_148 : _GEN_148; // @[ICache.scala 68:{44,44}]
  wire  _GEN_150 = 10'h95 == req_r_addr[14:5] ? valid_149 : _GEN_149; // @[ICache.scala 68:{44,44}]
  wire  _GEN_151 = 10'h96 == req_r_addr[14:5] ? valid_150 : _GEN_150; // @[ICache.scala 68:{44,44}]
  wire  _GEN_152 = 10'h97 == req_r_addr[14:5] ? valid_151 : _GEN_151; // @[ICache.scala 68:{44,44}]
  wire  _GEN_153 = 10'h98 == req_r_addr[14:5] ? valid_152 : _GEN_152; // @[ICache.scala 68:{44,44}]
  wire  _GEN_154 = 10'h99 == req_r_addr[14:5] ? valid_153 : _GEN_153; // @[ICache.scala 68:{44,44}]
  wire  _GEN_155 = 10'h9a == req_r_addr[14:5] ? valid_154 : _GEN_154; // @[ICache.scala 68:{44,44}]
  wire  _GEN_156 = 10'h9b == req_r_addr[14:5] ? valid_155 : _GEN_155; // @[ICache.scala 68:{44,44}]
  wire  _GEN_157 = 10'h9c == req_r_addr[14:5] ? valid_156 : _GEN_156; // @[ICache.scala 68:{44,44}]
  wire  _GEN_158 = 10'h9d == req_r_addr[14:5] ? valid_157 : _GEN_157; // @[ICache.scala 68:{44,44}]
  wire  _GEN_159 = 10'h9e == req_r_addr[14:5] ? valid_158 : _GEN_158; // @[ICache.scala 68:{44,44}]
  wire  _GEN_160 = 10'h9f == req_r_addr[14:5] ? valid_159 : _GEN_159; // @[ICache.scala 68:{44,44}]
  wire  _GEN_161 = 10'ha0 == req_r_addr[14:5] ? valid_160 : _GEN_160; // @[ICache.scala 68:{44,44}]
  wire  _GEN_162 = 10'ha1 == req_r_addr[14:5] ? valid_161 : _GEN_161; // @[ICache.scala 68:{44,44}]
  wire  _GEN_163 = 10'ha2 == req_r_addr[14:5] ? valid_162 : _GEN_162; // @[ICache.scala 68:{44,44}]
  wire  _GEN_164 = 10'ha3 == req_r_addr[14:5] ? valid_163 : _GEN_163; // @[ICache.scala 68:{44,44}]
  wire  _GEN_165 = 10'ha4 == req_r_addr[14:5] ? valid_164 : _GEN_164; // @[ICache.scala 68:{44,44}]
  wire  _GEN_166 = 10'ha5 == req_r_addr[14:5] ? valid_165 : _GEN_165; // @[ICache.scala 68:{44,44}]
  wire  _GEN_167 = 10'ha6 == req_r_addr[14:5] ? valid_166 : _GEN_166; // @[ICache.scala 68:{44,44}]
  wire  _GEN_168 = 10'ha7 == req_r_addr[14:5] ? valid_167 : _GEN_167; // @[ICache.scala 68:{44,44}]
  wire  _GEN_169 = 10'ha8 == req_r_addr[14:5] ? valid_168 : _GEN_168; // @[ICache.scala 68:{44,44}]
  wire  _GEN_170 = 10'ha9 == req_r_addr[14:5] ? valid_169 : _GEN_169; // @[ICache.scala 68:{44,44}]
  wire  _GEN_171 = 10'haa == req_r_addr[14:5] ? valid_170 : _GEN_170; // @[ICache.scala 68:{44,44}]
  wire  _GEN_172 = 10'hab == req_r_addr[14:5] ? valid_171 : _GEN_171; // @[ICache.scala 68:{44,44}]
  wire  _GEN_173 = 10'hac == req_r_addr[14:5] ? valid_172 : _GEN_172; // @[ICache.scala 68:{44,44}]
  wire  _GEN_174 = 10'had == req_r_addr[14:5] ? valid_173 : _GEN_173; // @[ICache.scala 68:{44,44}]
  wire  _GEN_175 = 10'hae == req_r_addr[14:5] ? valid_174 : _GEN_174; // @[ICache.scala 68:{44,44}]
  wire  _GEN_176 = 10'haf == req_r_addr[14:5] ? valid_175 : _GEN_175; // @[ICache.scala 68:{44,44}]
  wire  _GEN_177 = 10'hb0 == req_r_addr[14:5] ? valid_176 : _GEN_176; // @[ICache.scala 68:{44,44}]
  wire  _GEN_178 = 10'hb1 == req_r_addr[14:5] ? valid_177 : _GEN_177; // @[ICache.scala 68:{44,44}]
  wire  _GEN_179 = 10'hb2 == req_r_addr[14:5] ? valid_178 : _GEN_178; // @[ICache.scala 68:{44,44}]
  wire  _GEN_180 = 10'hb3 == req_r_addr[14:5] ? valid_179 : _GEN_179; // @[ICache.scala 68:{44,44}]
  wire  _GEN_181 = 10'hb4 == req_r_addr[14:5] ? valid_180 : _GEN_180; // @[ICache.scala 68:{44,44}]
  wire  _GEN_182 = 10'hb5 == req_r_addr[14:5] ? valid_181 : _GEN_181; // @[ICache.scala 68:{44,44}]
  wire  _GEN_183 = 10'hb6 == req_r_addr[14:5] ? valid_182 : _GEN_182; // @[ICache.scala 68:{44,44}]
  wire  _GEN_184 = 10'hb7 == req_r_addr[14:5] ? valid_183 : _GEN_183; // @[ICache.scala 68:{44,44}]
  wire  _GEN_185 = 10'hb8 == req_r_addr[14:5] ? valid_184 : _GEN_184; // @[ICache.scala 68:{44,44}]
  wire  _GEN_186 = 10'hb9 == req_r_addr[14:5] ? valid_185 : _GEN_185; // @[ICache.scala 68:{44,44}]
  wire  _GEN_187 = 10'hba == req_r_addr[14:5] ? valid_186 : _GEN_186; // @[ICache.scala 68:{44,44}]
  wire  _GEN_188 = 10'hbb == req_r_addr[14:5] ? valid_187 : _GEN_187; // @[ICache.scala 68:{44,44}]
  wire  _GEN_189 = 10'hbc == req_r_addr[14:5] ? valid_188 : _GEN_188; // @[ICache.scala 68:{44,44}]
  wire  _GEN_190 = 10'hbd == req_r_addr[14:5] ? valid_189 : _GEN_189; // @[ICache.scala 68:{44,44}]
  wire  _GEN_191 = 10'hbe == req_r_addr[14:5] ? valid_190 : _GEN_190; // @[ICache.scala 68:{44,44}]
  wire  _GEN_192 = 10'hbf == req_r_addr[14:5] ? valid_191 : _GEN_191; // @[ICache.scala 68:{44,44}]
  wire  _GEN_193 = 10'hc0 == req_r_addr[14:5] ? valid_192 : _GEN_192; // @[ICache.scala 68:{44,44}]
  wire  _GEN_194 = 10'hc1 == req_r_addr[14:5] ? valid_193 : _GEN_193; // @[ICache.scala 68:{44,44}]
  wire  _GEN_195 = 10'hc2 == req_r_addr[14:5] ? valid_194 : _GEN_194; // @[ICache.scala 68:{44,44}]
  wire  _GEN_196 = 10'hc3 == req_r_addr[14:5] ? valid_195 : _GEN_195; // @[ICache.scala 68:{44,44}]
  wire  _GEN_197 = 10'hc4 == req_r_addr[14:5] ? valid_196 : _GEN_196; // @[ICache.scala 68:{44,44}]
  wire  _GEN_198 = 10'hc5 == req_r_addr[14:5] ? valid_197 : _GEN_197; // @[ICache.scala 68:{44,44}]
  wire  _GEN_199 = 10'hc6 == req_r_addr[14:5] ? valid_198 : _GEN_198; // @[ICache.scala 68:{44,44}]
  wire  _GEN_200 = 10'hc7 == req_r_addr[14:5] ? valid_199 : _GEN_199; // @[ICache.scala 68:{44,44}]
  wire  _GEN_201 = 10'hc8 == req_r_addr[14:5] ? valid_200 : _GEN_200; // @[ICache.scala 68:{44,44}]
  wire  _GEN_202 = 10'hc9 == req_r_addr[14:5] ? valid_201 : _GEN_201; // @[ICache.scala 68:{44,44}]
  wire  _GEN_203 = 10'hca == req_r_addr[14:5] ? valid_202 : _GEN_202; // @[ICache.scala 68:{44,44}]
  wire  _GEN_204 = 10'hcb == req_r_addr[14:5] ? valid_203 : _GEN_203; // @[ICache.scala 68:{44,44}]
  wire  _GEN_205 = 10'hcc == req_r_addr[14:5] ? valid_204 : _GEN_204; // @[ICache.scala 68:{44,44}]
  wire  _GEN_206 = 10'hcd == req_r_addr[14:5] ? valid_205 : _GEN_205; // @[ICache.scala 68:{44,44}]
  wire  _GEN_207 = 10'hce == req_r_addr[14:5] ? valid_206 : _GEN_206; // @[ICache.scala 68:{44,44}]
  wire  _GEN_208 = 10'hcf == req_r_addr[14:5] ? valid_207 : _GEN_207; // @[ICache.scala 68:{44,44}]
  wire  _GEN_209 = 10'hd0 == req_r_addr[14:5] ? valid_208 : _GEN_208; // @[ICache.scala 68:{44,44}]
  wire  _GEN_210 = 10'hd1 == req_r_addr[14:5] ? valid_209 : _GEN_209; // @[ICache.scala 68:{44,44}]
  wire  _GEN_211 = 10'hd2 == req_r_addr[14:5] ? valid_210 : _GEN_210; // @[ICache.scala 68:{44,44}]
  wire  _GEN_212 = 10'hd3 == req_r_addr[14:5] ? valid_211 : _GEN_211; // @[ICache.scala 68:{44,44}]
  wire  _GEN_213 = 10'hd4 == req_r_addr[14:5] ? valid_212 : _GEN_212; // @[ICache.scala 68:{44,44}]
  wire  _GEN_214 = 10'hd5 == req_r_addr[14:5] ? valid_213 : _GEN_213; // @[ICache.scala 68:{44,44}]
  wire  _GEN_215 = 10'hd6 == req_r_addr[14:5] ? valid_214 : _GEN_214; // @[ICache.scala 68:{44,44}]
  wire  _GEN_216 = 10'hd7 == req_r_addr[14:5] ? valid_215 : _GEN_215; // @[ICache.scala 68:{44,44}]
  wire  _GEN_217 = 10'hd8 == req_r_addr[14:5] ? valid_216 : _GEN_216; // @[ICache.scala 68:{44,44}]
  wire  _GEN_218 = 10'hd9 == req_r_addr[14:5] ? valid_217 : _GEN_217; // @[ICache.scala 68:{44,44}]
  wire  _GEN_219 = 10'hda == req_r_addr[14:5] ? valid_218 : _GEN_218; // @[ICache.scala 68:{44,44}]
  wire  _GEN_220 = 10'hdb == req_r_addr[14:5] ? valid_219 : _GEN_219; // @[ICache.scala 68:{44,44}]
  wire  _GEN_221 = 10'hdc == req_r_addr[14:5] ? valid_220 : _GEN_220; // @[ICache.scala 68:{44,44}]
  wire  _GEN_222 = 10'hdd == req_r_addr[14:5] ? valid_221 : _GEN_221; // @[ICache.scala 68:{44,44}]
  wire  _GEN_223 = 10'hde == req_r_addr[14:5] ? valid_222 : _GEN_222; // @[ICache.scala 68:{44,44}]
  wire  _GEN_224 = 10'hdf == req_r_addr[14:5] ? valid_223 : _GEN_223; // @[ICache.scala 68:{44,44}]
  wire  _GEN_225 = 10'he0 == req_r_addr[14:5] ? valid_224 : _GEN_224; // @[ICache.scala 68:{44,44}]
  wire  _GEN_226 = 10'he1 == req_r_addr[14:5] ? valid_225 : _GEN_225; // @[ICache.scala 68:{44,44}]
  wire  _GEN_227 = 10'he2 == req_r_addr[14:5] ? valid_226 : _GEN_226; // @[ICache.scala 68:{44,44}]
  wire  _GEN_228 = 10'he3 == req_r_addr[14:5] ? valid_227 : _GEN_227; // @[ICache.scala 68:{44,44}]
  wire  _GEN_229 = 10'he4 == req_r_addr[14:5] ? valid_228 : _GEN_228; // @[ICache.scala 68:{44,44}]
  wire  _GEN_230 = 10'he5 == req_r_addr[14:5] ? valid_229 : _GEN_229; // @[ICache.scala 68:{44,44}]
  wire  _GEN_231 = 10'he6 == req_r_addr[14:5] ? valid_230 : _GEN_230; // @[ICache.scala 68:{44,44}]
  wire  _GEN_232 = 10'he7 == req_r_addr[14:5] ? valid_231 : _GEN_231; // @[ICache.scala 68:{44,44}]
  wire  _GEN_233 = 10'he8 == req_r_addr[14:5] ? valid_232 : _GEN_232; // @[ICache.scala 68:{44,44}]
  wire  _GEN_234 = 10'he9 == req_r_addr[14:5] ? valid_233 : _GEN_233; // @[ICache.scala 68:{44,44}]
  wire  _GEN_235 = 10'hea == req_r_addr[14:5] ? valid_234 : _GEN_234; // @[ICache.scala 68:{44,44}]
  wire  _GEN_236 = 10'heb == req_r_addr[14:5] ? valid_235 : _GEN_235; // @[ICache.scala 68:{44,44}]
  wire  _GEN_237 = 10'hec == req_r_addr[14:5] ? valid_236 : _GEN_236; // @[ICache.scala 68:{44,44}]
  wire  _GEN_238 = 10'hed == req_r_addr[14:5] ? valid_237 : _GEN_237; // @[ICache.scala 68:{44,44}]
  wire  _GEN_239 = 10'hee == req_r_addr[14:5] ? valid_238 : _GEN_238; // @[ICache.scala 68:{44,44}]
  wire  _GEN_240 = 10'hef == req_r_addr[14:5] ? valid_239 : _GEN_239; // @[ICache.scala 68:{44,44}]
  wire  _GEN_241 = 10'hf0 == req_r_addr[14:5] ? valid_240 : _GEN_240; // @[ICache.scala 68:{44,44}]
  wire  _GEN_242 = 10'hf1 == req_r_addr[14:5] ? valid_241 : _GEN_241; // @[ICache.scala 68:{44,44}]
  wire  _GEN_243 = 10'hf2 == req_r_addr[14:5] ? valid_242 : _GEN_242; // @[ICache.scala 68:{44,44}]
  wire  _GEN_244 = 10'hf3 == req_r_addr[14:5] ? valid_243 : _GEN_243; // @[ICache.scala 68:{44,44}]
  wire  _GEN_245 = 10'hf4 == req_r_addr[14:5] ? valid_244 : _GEN_244; // @[ICache.scala 68:{44,44}]
  wire  _GEN_246 = 10'hf5 == req_r_addr[14:5] ? valid_245 : _GEN_245; // @[ICache.scala 68:{44,44}]
  wire  _GEN_247 = 10'hf6 == req_r_addr[14:5] ? valid_246 : _GEN_246; // @[ICache.scala 68:{44,44}]
  wire  _GEN_248 = 10'hf7 == req_r_addr[14:5] ? valid_247 : _GEN_247; // @[ICache.scala 68:{44,44}]
  wire  _GEN_249 = 10'hf8 == req_r_addr[14:5] ? valid_248 : _GEN_248; // @[ICache.scala 68:{44,44}]
  wire  _GEN_250 = 10'hf9 == req_r_addr[14:5] ? valid_249 : _GEN_249; // @[ICache.scala 68:{44,44}]
  wire  _GEN_251 = 10'hfa == req_r_addr[14:5] ? valid_250 : _GEN_250; // @[ICache.scala 68:{44,44}]
  wire  _GEN_252 = 10'hfb == req_r_addr[14:5] ? valid_251 : _GEN_251; // @[ICache.scala 68:{44,44}]
  wire  _GEN_253 = 10'hfc == req_r_addr[14:5] ? valid_252 : _GEN_252; // @[ICache.scala 68:{44,44}]
  wire  _GEN_254 = 10'hfd == req_r_addr[14:5] ? valid_253 : _GEN_253; // @[ICache.scala 68:{44,44}]
  wire  _GEN_255 = 10'hfe == req_r_addr[14:5] ? valid_254 : _GEN_254; // @[ICache.scala 68:{44,44}]
  wire  _GEN_256 = 10'hff == req_r_addr[14:5] ? valid_255 : _GEN_255; // @[ICache.scala 68:{44,44}]
  wire  _GEN_257 = 10'h100 == req_r_addr[14:5] ? valid_256 : _GEN_256; // @[ICache.scala 68:{44,44}]
  wire  _GEN_258 = 10'h101 == req_r_addr[14:5] ? valid_257 : _GEN_257; // @[ICache.scala 68:{44,44}]
  wire  _GEN_259 = 10'h102 == req_r_addr[14:5] ? valid_258 : _GEN_258; // @[ICache.scala 68:{44,44}]
  wire  _GEN_260 = 10'h103 == req_r_addr[14:5] ? valid_259 : _GEN_259; // @[ICache.scala 68:{44,44}]
  wire  _GEN_261 = 10'h104 == req_r_addr[14:5] ? valid_260 : _GEN_260; // @[ICache.scala 68:{44,44}]
  wire  _GEN_262 = 10'h105 == req_r_addr[14:5] ? valid_261 : _GEN_261; // @[ICache.scala 68:{44,44}]
  wire  _GEN_263 = 10'h106 == req_r_addr[14:5] ? valid_262 : _GEN_262; // @[ICache.scala 68:{44,44}]
  wire  _GEN_264 = 10'h107 == req_r_addr[14:5] ? valid_263 : _GEN_263; // @[ICache.scala 68:{44,44}]
  wire  _GEN_265 = 10'h108 == req_r_addr[14:5] ? valid_264 : _GEN_264; // @[ICache.scala 68:{44,44}]
  wire  _GEN_266 = 10'h109 == req_r_addr[14:5] ? valid_265 : _GEN_265; // @[ICache.scala 68:{44,44}]
  wire  _GEN_267 = 10'h10a == req_r_addr[14:5] ? valid_266 : _GEN_266; // @[ICache.scala 68:{44,44}]
  wire  _GEN_268 = 10'h10b == req_r_addr[14:5] ? valid_267 : _GEN_267; // @[ICache.scala 68:{44,44}]
  wire  _GEN_269 = 10'h10c == req_r_addr[14:5] ? valid_268 : _GEN_268; // @[ICache.scala 68:{44,44}]
  wire  _GEN_270 = 10'h10d == req_r_addr[14:5] ? valid_269 : _GEN_269; // @[ICache.scala 68:{44,44}]
  wire  _GEN_271 = 10'h10e == req_r_addr[14:5] ? valid_270 : _GEN_270; // @[ICache.scala 68:{44,44}]
  wire  _GEN_272 = 10'h10f == req_r_addr[14:5] ? valid_271 : _GEN_271; // @[ICache.scala 68:{44,44}]
  wire  _GEN_273 = 10'h110 == req_r_addr[14:5] ? valid_272 : _GEN_272; // @[ICache.scala 68:{44,44}]
  wire  _GEN_274 = 10'h111 == req_r_addr[14:5] ? valid_273 : _GEN_273; // @[ICache.scala 68:{44,44}]
  wire  _GEN_275 = 10'h112 == req_r_addr[14:5] ? valid_274 : _GEN_274; // @[ICache.scala 68:{44,44}]
  wire  _GEN_276 = 10'h113 == req_r_addr[14:5] ? valid_275 : _GEN_275; // @[ICache.scala 68:{44,44}]
  wire  _GEN_277 = 10'h114 == req_r_addr[14:5] ? valid_276 : _GEN_276; // @[ICache.scala 68:{44,44}]
  wire  _GEN_278 = 10'h115 == req_r_addr[14:5] ? valid_277 : _GEN_277; // @[ICache.scala 68:{44,44}]
  wire  _GEN_279 = 10'h116 == req_r_addr[14:5] ? valid_278 : _GEN_278; // @[ICache.scala 68:{44,44}]
  wire  _GEN_280 = 10'h117 == req_r_addr[14:5] ? valid_279 : _GEN_279; // @[ICache.scala 68:{44,44}]
  wire  _GEN_281 = 10'h118 == req_r_addr[14:5] ? valid_280 : _GEN_280; // @[ICache.scala 68:{44,44}]
  wire  _GEN_282 = 10'h119 == req_r_addr[14:5] ? valid_281 : _GEN_281; // @[ICache.scala 68:{44,44}]
  wire  _GEN_283 = 10'h11a == req_r_addr[14:5] ? valid_282 : _GEN_282; // @[ICache.scala 68:{44,44}]
  wire  _GEN_284 = 10'h11b == req_r_addr[14:5] ? valid_283 : _GEN_283; // @[ICache.scala 68:{44,44}]
  wire  _GEN_285 = 10'h11c == req_r_addr[14:5] ? valid_284 : _GEN_284; // @[ICache.scala 68:{44,44}]
  wire  _GEN_286 = 10'h11d == req_r_addr[14:5] ? valid_285 : _GEN_285; // @[ICache.scala 68:{44,44}]
  wire  _GEN_287 = 10'h11e == req_r_addr[14:5] ? valid_286 : _GEN_286; // @[ICache.scala 68:{44,44}]
  wire  _GEN_288 = 10'h11f == req_r_addr[14:5] ? valid_287 : _GEN_287; // @[ICache.scala 68:{44,44}]
  wire  _GEN_289 = 10'h120 == req_r_addr[14:5] ? valid_288 : _GEN_288; // @[ICache.scala 68:{44,44}]
  wire  _GEN_290 = 10'h121 == req_r_addr[14:5] ? valid_289 : _GEN_289; // @[ICache.scala 68:{44,44}]
  wire  _GEN_291 = 10'h122 == req_r_addr[14:5] ? valid_290 : _GEN_290; // @[ICache.scala 68:{44,44}]
  wire  _GEN_292 = 10'h123 == req_r_addr[14:5] ? valid_291 : _GEN_291; // @[ICache.scala 68:{44,44}]
  wire  _GEN_293 = 10'h124 == req_r_addr[14:5] ? valid_292 : _GEN_292; // @[ICache.scala 68:{44,44}]
  wire  _GEN_294 = 10'h125 == req_r_addr[14:5] ? valid_293 : _GEN_293; // @[ICache.scala 68:{44,44}]
  wire  _GEN_295 = 10'h126 == req_r_addr[14:5] ? valid_294 : _GEN_294; // @[ICache.scala 68:{44,44}]
  wire  _GEN_296 = 10'h127 == req_r_addr[14:5] ? valid_295 : _GEN_295; // @[ICache.scala 68:{44,44}]
  wire  _GEN_297 = 10'h128 == req_r_addr[14:5] ? valid_296 : _GEN_296; // @[ICache.scala 68:{44,44}]
  wire  _GEN_298 = 10'h129 == req_r_addr[14:5] ? valid_297 : _GEN_297; // @[ICache.scala 68:{44,44}]
  wire  _GEN_299 = 10'h12a == req_r_addr[14:5] ? valid_298 : _GEN_298; // @[ICache.scala 68:{44,44}]
  wire  _GEN_300 = 10'h12b == req_r_addr[14:5] ? valid_299 : _GEN_299; // @[ICache.scala 68:{44,44}]
  wire  _GEN_301 = 10'h12c == req_r_addr[14:5] ? valid_300 : _GEN_300; // @[ICache.scala 68:{44,44}]
  wire  _GEN_302 = 10'h12d == req_r_addr[14:5] ? valid_301 : _GEN_301; // @[ICache.scala 68:{44,44}]
  wire  _GEN_303 = 10'h12e == req_r_addr[14:5] ? valid_302 : _GEN_302; // @[ICache.scala 68:{44,44}]
  wire  _GEN_304 = 10'h12f == req_r_addr[14:5] ? valid_303 : _GEN_303; // @[ICache.scala 68:{44,44}]
  wire  _GEN_305 = 10'h130 == req_r_addr[14:5] ? valid_304 : _GEN_304; // @[ICache.scala 68:{44,44}]
  wire  _GEN_306 = 10'h131 == req_r_addr[14:5] ? valid_305 : _GEN_305; // @[ICache.scala 68:{44,44}]
  wire  _GEN_307 = 10'h132 == req_r_addr[14:5] ? valid_306 : _GEN_306; // @[ICache.scala 68:{44,44}]
  wire  _GEN_308 = 10'h133 == req_r_addr[14:5] ? valid_307 : _GEN_307; // @[ICache.scala 68:{44,44}]
  wire  _GEN_309 = 10'h134 == req_r_addr[14:5] ? valid_308 : _GEN_308; // @[ICache.scala 68:{44,44}]
  wire  _GEN_310 = 10'h135 == req_r_addr[14:5] ? valid_309 : _GEN_309; // @[ICache.scala 68:{44,44}]
  wire  _GEN_311 = 10'h136 == req_r_addr[14:5] ? valid_310 : _GEN_310; // @[ICache.scala 68:{44,44}]
  wire  _GEN_312 = 10'h137 == req_r_addr[14:5] ? valid_311 : _GEN_311; // @[ICache.scala 68:{44,44}]
  wire  _GEN_313 = 10'h138 == req_r_addr[14:5] ? valid_312 : _GEN_312; // @[ICache.scala 68:{44,44}]
  wire  _GEN_314 = 10'h139 == req_r_addr[14:5] ? valid_313 : _GEN_313; // @[ICache.scala 68:{44,44}]
  wire  _GEN_315 = 10'h13a == req_r_addr[14:5] ? valid_314 : _GEN_314; // @[ICache.scala 68:{44,44}]
  wire  _GEN_316 = 10'h13b == req_r_addr[14:5] ? valid_315 : _GEN_315; // @[ICache.scala 68:{44,44}]
  wire  _GEN_317 = 10'h13c == req_r_addr[14:5] ? valid_316 : _GEN_316; // @[ICache.scala 68:{44,44}]
  wire  _GEN_318 = 10'h13d == req_r_addr[14:5] ? valid_317 : _GEN_317; // @[ICache.scala 68:{44,44}]
  wire  _GEN_319 = 10'h13e == req_r_addr[14:5] ? valid_318 : _GEN_318; // @[ICache.scala 68:{44,44}]
  wire  _GEN_320 = 10'h13f == req_r_addr[14:5] ? valid_319 : _GEN_319; // @[ICache.scala 68:{44,44}]
  wire  _GEN_321 = 10'h140 == req_r_addr[14:5] ? valid_320 : _GEN_320; // @[ICache.scala 68:{44,44}]
  wire  _GEN_322 = 10'h141 == req_r_addr[14:5] ? valid_321 : _GEN_321; // @[ICache.scala 68:{44,44}]
  wire  _GEN_323 = 10'h142 == req_r_addr[14:5] ? valid_322 : _GEN_322; // @[ICache.scala 68:{44,44}]
  wire  _GEN_324 = 10'h143 == req_r_addr[14:5] ? valid_323 : _GEN_323; // @[ICache.scala 68:{44,44}]
  wire  _GEN_325 = 10'h144 == req_r_addr[14:5] ? valid_324 : _GEN_324; // @[ICache.scala 68:{44,44}]
  wire  _GEN_326 = 10'h145 == req_r_addr[14:5] ? valid_325 : _GEN_325; // @[ICache.scala 68:{44,44}]
  wire  _GEN_327 = 10'h146 == req_r_addr[14:5] ? valid_326 : _GEN_326; // @[ICache.scala 68:{44,44}]
  wire  _GEN_328 = 10'h147 == req_r_addr[14:5] ? valid_327 : _GEN_327; // @[ICache.scala 68:{44,44}]
  wire  _GEN_329 = 10'h148 == req_r_addr[14:5] ? valid_328 : _GEN_328; // @[ICache.scala 68:{44,44}]
  wire  _GEN_330 = 10'h149 == req_r_addr[14:5] ? valid_329 : _GEN_329; // @[ICache.scala 68:{44,44}]
  wire  _GEN_331 = 10'h14a == req_r_addr[14:5] ? valid_330 : _GEN_330; // @[ICache.scala 68:{44,44}]
  wire  _GEN_332 = 10'h14b == req_r_addr[14:5] ? valid_331 : _GEN_331; // @[ICache.scala 68:{44,44}]
  wire  _GEN_333 = 10'h14c == req_r_addr[14:5] ? valid_332 : _GEN_332; // @[ICache.scala 68:{44,44}]
  wire  _GEN_334 = 10'h14d == req_r_addr[14:5] ? valid_333 : _GEN_333; // @[ICache.scala 68:{44,44}]
  wire  _GEN_335 = 10'h14e == req_r_addr[14:5] ? valid_334 : _GEN_334; // @[ICache.scala 68:{44,44}]
  wire  _GEN_336 = 10'h14f == req_r_addr[14:5] ? valid_335 : _GEN_335; // @[ICache.scala 68:{44,44}]
  wire  _GEN_337 = 10'h150 == req_r_addr[14:5] ? valid_336 : _GEN_336; // @[ICache.scala 68:{44,44}]
  wire  _GEN_338 = 10'h151 == req_r_addr[14:5] ? valid_337 : _GEN_337; // @[ICache.scala 68:{44,44}]
  wire  _GEN_339 = 10'h152 == req_r_addr[14:5] ? valid_338 : _GEN_338; // @[ICache.scala 68:{44,44}]
  wire  _GEN_340 = 10'h153 == req_r_addr[14:5] ? valid_339 : _GEN_339; // @[ICache.scala 68:{44,44}]
  wire  _GEN_341 = 10'h154 == req_r_addr[14:5] ? valid_340 : _GEN_340; // @[ICache.scala 68:{44,44}]
  wire  _GEN_342 = 10'h155 == req_r_addr[14:5] ? valid_341 : _GEN_341; // @[ICache.scala 68:{44,44}]
  wire  _GEN_343 = 10'h156 == req_r_addr[14:5] ? valid_342 : _GEN_342; // @[ICache.scala 68:{44,44}]
  wire  _GEN_344 = 10'h157 == req_r_addr[14:5] ? valid_343 : _GEN_343; // @[ICache.scala 68:{44,44}]
  wire  _GEN_345 = 10'h158 == req_r_addr[14:5] ? valid_344 : _GEN_344; // @[ICache.scala 68:{44,44}]
  wire  _GEN_346 = 10'h159 == req_r_addr[14:5] ? valid_345 : _GEN_345; // @[ICache.scala 68:{44,44}]
  wire  _GEN_347 = 10'h15a == req_r_addr[14:5] ? valid_346 : _GEN_346; // @[ICache.scala 68:{44,44}]
  wire  _GEN_348 = 10'h15b == req_r_addr[14:5] ? valid_347 : _GEN_347; // @[ICache.scala 68:{44,44}]
  wire  _GEN_349 = 10'h15c == req_r_addr[14:5] ? valid_348 : _GEN_348; // @[ICache.scala 68:{44,44}]
  wire  _GEN_350 = 10'h15d == req_r_addr[14:5] ? valid_349 : _GEN_349; // @[ICache.scala 68:{44,44}]
  wire  _GEN_351 = 10'h15e == req_r_addr[14:5] ? valid_350 : _GEN_350; // @[ICache.scala 68:{44,44}]
  wire  _GEN_352 = 10'h15f == req_r_addr[14:5] ? valid_351 : _GEN_351; // @[ICache.scala 68:{44,44}]
  wire  _GEN_353 = 10'h160 == req_r_addr[14:5] ? valid_352 : _GEN_352; // @[ICache.scala 68:{44,44}]
  wire  _GEN_354 = 10'h161 == req_r_addr[14:5] ? valid_353 : _GEN_353; // @[ICache.scala 68:{44,44}]
  wire  _GEN_355 = 10'h162 == req_r_addr[14:5] ? valid_354 : _GEN_354; // @[ICache.scala 68:{44,44}]
  wire  _GEN_356 = 10'h163 == req_r_addr[14:5] ? valid_355 : _GEN_355; // @[ICache.scala 68:{44,44}]
  wire  _GEN_357 = 10'h164 == req_r_addr[14:5] ? valid_356 : _GEN_356; // @[ICache.scala 68:{44,44}]
  wire  _GEN_358 = 10'h165 == req_r_addr[14:5] ? valid_357 : _GEN_357; // @[ICache.scala 68:{44,44}]
  wire  _GEN_359 = 10'h166 == req_r_addr[14:5] ? valid_358 : _GEN_358; // @[ICache.scala 68:{44,44}]
  wire  _GEN_360 = 10'h167 == req_r_addr[14:5] ? valid_359 : _GEN_359; // @[ICache.scala 68:{44,44}]
  wire  _GEN_361 = 10'h168 == req_r_addr[14:5] ? valid_360 : _GEN_360; // @[ICache.scala 68:{44,44}]
  wire  _GEN_362 = 10'h169 == req_r_addr[14:5] ? valid_361 : _GEN_361; // @[ICache.scala 68:{44,44}]
  wire  _GEN_363 = 10'h16a == req_r_addr[14:5] ? valid_362 : _GEN_362; // @[ICache.scala 68:{44,44}]
  wire  _GEN_364 = 10'h16b == req_r_addr[14:5] ? valid_363 : _GEN_363; // @[ICache.scala 68:{44,44}]
  wire  _GEN_365 = 10'h16c == req_r_addr[14:5] ? valid_364 : _GEN_364; // @[ICache.scala 68:{44,44}]
  wire  _GEN_366 = 10'h16d == req_r_addr[14:5] ? valid_365 : _GEN_365; // @[ICache.scala 68:{44,44}]
  wire  _GEN_367 = 10'h16e == req_r_addr[14:5] ? valid_366 : _GEN_366; // @[ICache.scala 68:{44,44}]
  wire  _GEN_368 = 10'h16f == req_r_addr[14:5] ? valid_367 : _GEN_367; // @[ICache.scala 68:{44,44}]
  wire  _GEN_369 = 10'h170 == req_r_addr[14:5] ? valid_368 : _GEN_368; // @[ICache.scala 68:{44,44}]
  wire  _GEN_370 = 10'h171 == req_r_addr[14:5] ? valid_369 : _GEN_369; // @[ICache.scala 68:{44,44}]
  wire  _GEN_371 = 10'h172 == req_r_addr[14:5] ? valid_370 : _GEN_370; // @[ICache.scala 68:{44,44}]
  wire  _GEN_372 = 10'h173 == req_r_addr[14:5] ? valid_371 : _GEN_371; // @[ICache.scala 68:{44,44}]
  wire  _GEN_373 = 10'h174 == req_r_addr[14:5] ? valid_372 : _GEN_372; // @[ICache.scala 68:{44,44}]
  wire  _GEN_374 = 10'h175 == req_r_addr[14:5] ? valid_373 : _GEN_373; // @[ICache.scala 68:{44,44}]
  wire  _GEN_375 = 10'h176 == req_r_addr[14:5] ? valid_374 : _GEN_374; // @[ICache.scala 68:{44,44}]
  wire  _GEN_376 = 10'h177 == req_r_addr[14:5] ? valid_375 : _GEN_375; // @[ICache.scala 68:{44,44}]
  wire  _GEN_377 = 10'h178 == req_r_addr[14:5] ? valid_376 : _GEN_376; // @[ICache.scala 68:{44,44}]
  wire  _GEN_378 = 10'h179 == req_r_addr[14:5] ? valid_377 : _GEN_377; // @[ICache.scala 68:{44,44}]
  wire  _GEN_379 = 10'h17a == req_r_addr[14:5] ? valid_378 : _GEN_378; // @[ICache.scala 68:{44,44}]
  wire  _GEN_380 = 10'h17b == req_r_addr[14:5] ? valid_379 : _GEN_379; // @[ICache.scala 68:{44,44}]
  wire  _GEN_381 = 10'h17c == req_r_addr[14:5] ? valid_380 : _GEN_380; // @[ICache.scala 68:{44,44}]
  wire  _GEN_382 = 10'h17d == req_r_addr[14:5] ? valid_381 : _GEN_381; // @[ICache.scala 68:{44,44}]
  wire  _GEN_383 = 10'h17e == req_r_addr[14:5] ? valid_382 : _GEN_382; // @[ICache.scala 68:{44,44}]
  wire  _GEN_384 = 10'h17f == req_r_addr[14:5] ? valid_383 : _GEN_383; // @[ICache.scala 68:{44,44}]
  wire  _GEN_385 = 10'h180 == req_r_addr[14:5] ? valid_384 : _GEN_384; // @[ICache.scala 68:{44,44}]
  wire  _GEN_386 = 10'h181 == req_r_addr[14:5] ? valid_385 : _GEN_385; // @[ICache.scala 68:{44,44}]
  wire  _GEN_387 = 10'h182 == req_r_addr[14:5] ? valid_386 : _GEN_386; // @[ICache.scala 68:{44,44}]
  wire  _GEN_388 = 10'h183 == req_r_addr[14:5] ? valid_387 : _GEN_387; // @[ICache.scala 68:{44,44}]
  wire  _GEN_389 = 10'h184 == req_r_addr[14:5] ? valid_388 : _GEN_388; // @[ICache.scala 68:{44,44}]
  wire  _GEN_390 = 10'h185 == req_r_addr[14:5] ? valid_389 : _GEN_389; // @[ICache.scala 68:{44,44}]
  wire  _GEN_391 = 10'h186 == req_r_addr[14:5] ? valid_390 : _GEN_390; // @[ICache.scala 68:{44,44}]
  wire  _GEN_392 = 10'h187 == req_r_addr[14:5] ? valid_391 : _GEN_391; // @[ICache.scala 68:{44,44}]
  wire  _GEN_393 = 10'h188 == req_r_addr[14:5] ? valid_392 : _GEN_392; // @[ICache.scala 68:{44,44}]
  wire  _GEN_394 = 10'h189 == req_r_addr[14:5] ? valid_393 : _GEN_393; // @[ICache.scala 68:{44,44}]
  wire  _GEN_395 = 10'h18a == req_r_addr[14:5] ? valid_394 : _GEN_394; // @[ICache.scala 68:{44,44}]
  wire  _GEN_396 = 10'h18b == req_r_addr[14:5] ? valid_395 : _GEN_395; // @[ICache.scala 68:{44,44}]
  wire  _GEN_397 = 10'h18c == req_r_addr[14:5] ? valid_396 : _GEN_396; // @[ICache.scala 68:{44,44}]
  wire  _GEN_398 = 10'h18d == req_r_addr[14:5] ? valid_397 : _GEN_397; // @[ICache.scala 68:{44,44}]
  wire  _GEN_399 = 10'h18e == req_r_addr[14:5] ? valid_398 : _GEN_398; // @[ICache.scala 68:{44,44}]
  wire  _GEN_400 = 10'h18f == req_r_addr[14:5] ? valid_399 : _GEN_399; // @[ICache.scala 68:{44,44}]
  wire  _GEN_401 = 10'h190 == req_r_addr[14:5] ? valid_400 : _GEN_400; // @[ICache.scala 68:{44,44}]
  wire  _GEN_402 = 10'h191 == req_r_addr[14:5] ? valid_401 : _GEN_401; // @[ICache.scala 68:{44,44}]
  wire  _GEN_403 = 10'h192 == req_r_addr[14:5] ? valid_402 : _GEN_402; // @[ICache.scala 68:{44,44}]
  wire  _GEN_404 = 10'h193 == req_r_addr[14:5] ? valid_403 : _GEN_403; // @[ICache.scala 68:{44,44}]
  wire  _GEN_405 = 10'h194 == req_r_addr[14:5] ? valid_404 : _GEN_404; // @[ICache.scala 68:{44,44}]
  wire  _GEN_406 = 10'h195 == req_r_addr[14:5] ? valid_405 : _GEN_405; // @[ICache.scala 68:{44,44}]
  wire  _GEN_407 = 10'h196 == req_r_addr[14:5] ? valid_406 : _GEN_406; // @[ICache.scala 68:{44,44}]
  wire  _GEN_408 = 10'h197 == req_r_addr[14:5] ? valid_407 : _GEN_407; // @[ICache.scala 68:{44,44}]
  wire  _GEN_409 = 10'h198 == req_r_addr[14:5] ? valid_408 : _GEN_408; // @[ICache.scala 68:{44,44}]
  wire  _GEN_410 = 10'h199 == req_r_addr[14:5] ? valid_409 : _GEN_409; // @[ICache.scala 68:{44,44}]
  wire  _GEN_411 = 10'h19a == req_r_addr[14:5] ? valid_410 : _GEN_410; // @[ICache.scala 68:{44,44}]
  wire  _GEN_412 = 10'h19b == req_r_addr[14:5] ? valid_411 : _GEN_411; // @[ICache.scala 68:{44,44}]
  wire  _GEN_413 = 10'h19c == req_r_addr[14:5] ? valid_412 : _GEN_412; // @[ICache.scala 68:{44,44}]
  wire  _GEN_414 = 10'h19d == req_r_addr[14:5] ? valid_413 : _GEN_413; // @[ICache.scala 68:{44,44}]
  wire  _GEN_415 = 10'h19e == req_r_addr[14:5] ? valid_414 : _GEN_414; // @[ICache.scala 68:{44,44}]
  wire  _GEN_416 = 10'h19f == req_r_addr[14:5] ? valid_415 : _GEN_415; // @[ICache.scala 68:{44,44}]
  wire  _GEN_417 = 10'h1a0 == req_r_addr[14:5] ? valid_416 : _GEN_416; // @[ICache.scala 68:{44,44}]
  wire  _GEN_418 = 10'h1a1 == req_r_addr[14:5] ? valid_417 : _GEN_417; // @[ICache.scala 68:{44,44}]
  wire  _GEN_419 = 10'h1a2 == req_r_addr[14:5] ? valid_418 : _GEN_418; // @[ICache.scala 68:{44,44}]
  wire  _GEN_420 = 10'h1a3 == req_r_addr[14:5] ? valid_419 : _GEN_419; // @[ICache.scala 68:{44,44}]
  wire  _GEN_421 = 10'h1a4 == req_r_addr[14:5] ? valid_420 : _GEN_420; // @[ICache.scala 68:{44,44}]
  wire  _GEN_422 = 10'h1a5 == req_r_addr[14:5] ? valid_421 : _GEN_421; // @[ICache.scala 68:{44,44}]
  wire  _GEN_423 = 10'h1a6 == req_r_addr[14:5] ? valid_422 : _GEN_422; // @[ICache.scala 68:{44,44}]
  wire  _GEN_424 = 10'h1a7 == req_r_addr[14:5] ? valid_423 : _GEN_423; // @[ICache.scala 68:{44,44}]
  wire  _GEN_425 = 10'h1a8 == req_r_addr[14:5] ? valid_424 : _GEN_424; // @[ICache.scala 68:{44,44}]
  wire  _GEN_426 = 10'h1a9 == req_r_addr[14:5] ? valid_425 : _GEN_425; // @[ICache.scala 68:{44,44}]
  wire  _GEN_427 = 10'h1aa == req_r_addr[14:5] ? valid_426 : _GEN_426; // @[ICache.scala 68:{44,44}]
  wire  _GEN_428 = 10'h1ab == req_r_addr[14:5] ? valid_427 : _GEN_427; // @[ICache.scala 68:{44,44}]
  wire  _GEN_429 = 10'h1ac == req_r_addr[14:5] ? valid_428 : _GEN_428; // @[ICache.scala 68:{44,44}]
  wire  _GEN_430 = 10'h1ad == req_r_addr[14:5] ? valid_429 : _GEN_429; // @[ICache.scala 68:{44,44}]
  wire  _GEN_431 = 10'h1ae == req_r_addr[14:5] ? valid_430 : _GEN_430; // @[ICache.scala 68:{44,44}]
  wire  _GEN_432 = 10'h1af == req_r_addr[14:5] ? valid_431 : _GEN_431; // @[ICache.scala 68:{44,44}]
  wire  _GEN_433 = 10'h1b0 == req_r_addr[14:5] ? valid_432 : _GEN_432; // @[ICache.scala 68:{44,44}]
  wire  _GEN_434 = 10'h1b1 == req_r_addr[14:5] ? valid_433 : _GEN_433; // @[ICache.scala 68:{44,44}]
  wire  _GEN_435 = 10'h1b2 == req_r_addr[14:5] ? valid_434 : _GEN_434; // @[ICache.scala 68:{44,44}]
  wire  _GEN_436 = 10'h1b3 == req_r_addr[14:5] ? valid_435 : _GEN_435; // @[ICache.scala 68:{44,44}]
  wire  _GEN_437 = 10'h1b4 == req_r_addr[14:5] ? valid_436 : _GEN_436; // @[ICache.scala 68:{44,44}]
  wire  _GEN_438 = 10'h1b5 == req_r_addr[14:5] ? valid_437 : _GEN_437; // @[ICache.scala 68:{44,44}]
  wire  _GEN_439 = 10'h1b6 == req_r_addr[14:5] ? valid_438 : _GEN_438; // @[ICache.scala 68:{44,44}]
  wire  _GEN_440 = 10'h1b7 == req_r_addr[14:5] ? valid_439 : _GEN_439; // @[ICache.scala 68:{44,44}]
  wire  _GEN_441 = 10'h1b8 == req_r_addr[14:5] ? valid_440 : _GEN_440; // @[ICache.scala 68:{44,44}]
  wire  _GEN_442 = 10'h1b9 == req_r_addr[14:5] ? valid_441 : _GEN_441; // @[ICache.scala 68:{44,44}]
  wire  _GEN_443 = 10'h1ba == req_r_addr[14:5] ? valid_442 : _GEN_442; // @[ICache.scala 68:{44,44}]
  wire  _GEN_444 = 10'h1bb == req_r_addr[14:5] ? valid_443 : _GEN_443; // @[ICache.scala 68:{44,44}]
  wire  _GEN_445 = 10'h1bc == req_r_addr[14:5] ? valid_444 : _GEN_444; // @[ICache.scala 68:{44,44}]
  wire  _GEN_446 = 10'h1bd == req_r_addr[14:5] ? valid_445 : _GEN_445; // @[ICache.scala 68:{44,44}]
  wire  _GEN_447 = 10'h1be == req_r_addr[14:5] ? valid_446 : _GEN_446; // @[ICache.scala 68:{44,44}]
  wire  _GEN_448 = 10'h1bf == req_r_addr[14:5] ? valid_447 : _GEN_447; // @[ICache.scala 68:{44,44}]
  wire  _GEN_449 = 10'h1c0 == req_r_addr[14:5] ? valid_448 : _GEN_448; // @[ICache.scala 68:{44,44}]
  wire  _GEN_450 = 10'h1c1 == req_r_addr[14:5] ? valid_449 : _GEN_449; // @[ICache.scala 68:{44,44}]
  wire  _GEN_451 = 10'h1c2 == req_r_addr[14:5] ? valid_450 : _GEN_450; // @[ICache.scala 68:{44,44}]
  wire  _GEN_452 = 10'h1c3 == req_r_addr[14:5] ? valid_451 : _GEN_451; // @[ICache.scala 68:{44,44}]
  wire  _GEN_453 = 10'h1c4 == req_r_addr[14:5] ? valid_452 : _GEN_452; // @[ICache.scala 68:{44,44}]
  wire  _GEN_454 = 10'h1c5 == req_r_addr[14:5] ? valid_453 : _GEN_453; // @[ICache.scala 68:{44,44}]
  wire  _GEN_455 = 10'h1c6 == req_r_addr[14:5] ? valid_454 : _GEN_454; // @[ICache.scala 68:{44,44}]
  wire  _GEN_456 = 10'h1c7 == req_r_addr[14:5] ? valid_455 : _GEN_455; // @[ICache.scala 68:{44,44}]
  wire  _GEN_457 = 10'h1c8 == req_r_addr[14:5] ? valid_456 : _GEN_456; // @[ICache.scala 68:{44,44}]
  wire  _GEN_458 = 10'h1c9 == req_r_addr[14:5] ? valid_457 : _GEN_457; // @[ICache.scala 68:{44,44}]
  wire  _GEN_459 = 10'h1ca == req_r_addr[14:5] ? valid_458 : _GEN_458; // @[ICache.scala 68:{44,44}]
  wire  _GEN_460 = 10'h1cb == req_r_addr[14:5] ? valid_459 : _GEN_459; // @[ICache.scala 68:{44,44}]
  wire  _GEN_461 = 10'h1cc == req_r_addr[14:5] ? valid_460 : _GEN_460; // @[ICache.scala 68:{44,44}]
  wire  _GEN_462 = 10'h1cd == req_r_addr[14:5] ? valid_461 : _GEN_461; // @[ICache.scala 68:{44,44}]
  wire  _GEN_463 = 10'h1ce == req_r_addr[14:5] ? valid_462 : _GEN_462; // @[ICache.scala 68:{44,44}]
  wire  _GEN_464 = 10'h1cf == req_r_addr[14:5] ? valid_463 : _GEN_463; // @[ICache.scala 68:{44,44}]
  wire  _GEN_465 = 10'h1d0 == req_r_addr[14:5] ? valid_464 : _GEN_464; // @[ICache.scala 68:{44,44}]
  wire  _GEN_466 = 10'h1d1 == req_r_addr[14:5] ? valid_465 : _GEN_465; // @[ICache.scala 68:{44,44}]
  wire  _GEN_467 = 10'h1d2 == req_r_addr[14:5] ? valid_466 : _GEN_466; // @[ICache.scala 68:{44,44}]
  wire  _GEN_468 = 10'h1d3 == req_r_addr[14:5] ? valid_467 : _GEN_467; // @[ICache.scala 68:{44,44}]
  wire  _GEN_469 = 10'h1d4 == req_r_addr[14:5] ? valid_468 : _GEN_468; // @[ICache.scala 68:{44,44}]
  wire  _GEN_470 = 10'h1d5 == req_r_addr[14:5] ? valid_469 : _GEN_469; // @[ICache.scala 68:{44,44}]
  wire  _GEN_471 = 10'h1d6 == req_r_addr[14:5] ? valid_470 : _GEN_470; // @[ICache.scala 68:{44,44}]
  wire  _GEN_472 = 10'h1d7 == req_r_addr[14:5] ? valid_471 : _GEN_471; // @[ICache.scala 68:{44,44}]
  wire  _GEN_473 = 10'h1d8 == req_r_addr[14:5] ? valid_472 : _GEN_472; // @[ICache.scala 68:{44,44}]
  wire  _GEN_474 = 10'h1d9 == req_r_addr[14:5] ? valid_473 : _GEN_473; // @[ICache.scala 68:{44,44}]
  wire  _GEN_475 = 10'h1da == req_r_addr[14:5] ? valid_474 : _GEN_474; // @[ICache.scala 68:{44,44}]
  wire  _GEN_476 = 10'h1db == req_r_addr[14:5] ? valid_475 : _GEN_475; // @[ICache.scala 68:{44,44}]
  wire  _GEN_477 = 10'h1dc == req_r_addr[14:5] ? valid_476 : _GEN_476; // @[ICache.scala 68:{44,44}]
  wire  _GEN_478 = 10'h1dd == req_r_addr[14:5] ? valid_477 : _GEN_477; // @[ICache.scala 68:{44,44}]
  wire  _GEN_479 = 10'h1de == req_r_addr[14:5] ? valid_478 : _GEN_478; // @[ICache.scala 68:{44,44}]
  wire  _GEN_480 = 10'h1df == req_r_addr[14:5] ? valid_479 : _GEN_479; // @[ICache.scala 68:{44,44}]
  wire  _GEN_481 = 10'h1e0 == req_r_addr[14:5] ? valid_480 : _GEN_480; // @[ICache.scala 68:{44,44}]
  wire  _GEN_482 = 10'h1e1 == req_r_addr[14:5] ? valid_481 : _GEN_481; // @[ICache.scala 68:{44,44}]
  wire  _GEN_483 = 10'h1e2 == req_r_addr[14:5] ? valid_482 : _GEN_482; // @[ICache.scala 68:{44,44}]
  wire  _GEN_484 = 10'h1e3 == req_r_addr[14:5] ? valid_483 : _GEN_483; // @[ICache.scala 68:{44,44}]
  wire  _GEN_485 = 10'h1e4 == req_r_addr[14:5] ? valid_484 : _GEN_484; // @[ICache.scala 68:{44,44}]
  wire  _GEN_486 = 10'h1e5 == req_r_addr[14:5] ? valid_485 : _GEN_485; // @[ICache.scala 68:{44,44}]
  wire  _GEN_487 = 10'h1e6 == req_r_addr[14:5] ? valid_486 : _GEN_486; // @[ICache.scala 68:{44,44}]
  wire  _GEN_488 = 10'h1e7 == req_r_addr[14:5] ? valid_487 : _GEN_487; // @[ICache.scala 68:{44,44}]
  wire  _GEN_489 = 10'h1e8 == req_r_addr[14:5] ? valid_488 : _GEN_488; // @[ICache.scala 68:{44,44}]
  wire  _GEN_490 = 10'h1e9 == req_r_addr[14:5] ? valid_489 : _GEN_489; // @[ICache.scala 68:{44,44}]
  wire  _GEN_491 = 10'h1ea == req_r_addr[14:5] ? valid_490 : _GEN_490; // @[ICache.scala 68:{44,44}]
  wire  _GEN_492 = 10'h1eb == req_r_addr[14:5] ? valid_491 : _GEN_491; // @[ICache.scala 68:{44,44}]
  wire  _GEN_493 = 10'h1ec == req_r_addr[14:5] ? valid_492 : _GEN_492; // @[ICache.scala 68:{44,44}]
  wire  _GEN_494 = 10'h1ed == req_r_addr[14:5] ? valid_493 : _GEN_493; // @[ICache.scala 68:{44,44}]
  wire  _GEN_495 = 10'h1ee == req_r_addr[14:5] ? valid_494 : _GEN_494; // @[ICache.scala 68:{44,44}]
  wire  _GEN_496 = 10'h1ef == req_r_addr[14:5] ? valid_495 : _GEN_495; // @[ICache.scala 68:{44,44}]
  wire  _GEN_497 = 10'h1f0 == req_r_addr[14:5] ? valid_496 : _GEN_496; // @[ICache.scala 68:{44,44}]
  wire  _GEN_498 = 10'h1f1 == req_r_addr[14:5] ? valid_497 : _GEN_497; // @[ICache.scala 68:{44,44}]
  wire  _GEN_499 = 10'h1f2 == req_r_addr[14:5] ? valid_498 : _GEN_498; // @[ICache.scala 68:{44,44}]
  wire  _GEN_500 = 10'h1f3 == req_r_addr[14:5] ? valid_499 : _GEN_499; // @[ICache.scala 68:{44,44}]
  wire  _GEN_501 = 10'h1f4 == req_r_addr[14:5] ? valid_500 : _GEN_500; // @[ICache.scala 68:{44,44}]
  wire  _GEN_502 = 10'h1f5 == req_r_addr[14:5] ? valid_501 : _GEN_501; // @[ICache.scala 68:{44,44}]
  wire  _GEN_503 = 10'h1f6 == req_r_addr[14:5] ? valid_502 : _GEN_502; // @[ICache.scala 68:{44,44}]
  wire  _GEN_504 = 10'h1f7 == req_r_addr[14:5] ? valid_503 : _GEN_503; // @[ICache.scala 68:{44,44}]
  wire  _GEN_505 = 10'h1f8 == req_r_addr[14:5] ? valid_504 : _GEN_504; // @[ICache.scala 68:{44,44}]
  wire  _GEN_506 = 10'h1f9 == req_r_addr[14:5] ? valid_505 : _GEN_505; // @[ICache.scala 68:{44,44}]
  wire  _GEN_507 = 10'h1fa == req_r_addr[14:5] ? valid_506 : _GEN_506; // @[ICache.scala 68:{44,44}]
  wire  _GEN_508 = 10'h1fb == req_r_addr[14:5] ? valid_507 : _GEN_507; // @[ICache.scala 68:{44,44}]
  wire  _GEN_509 = 10'h1fc == req_r_addr[14:5] ? valid_508 : _GEN_508; // @[ICache.scala 68:{44,44}]
  wire  _GEN_510 = 10'h1fd == req_r_addr[14:5] ? valid_509 : _GEN_509; // @[ICache.scala 68:{44,44}]
  wire  _GEN_511 = 10'h1fe == req_r_addr[14:5] ? valid_510 : _GEN_510; // @[ICache.scala 68:{44,44}]
  wire  _GEN_512 = 10'h1ff == req_r_addr[14:5] ? valid_511 : _GEN_511; // @[ICache.scala 68:{44,44}]
  wire  _GEN_513 = 10'h200 == req_r_addr[14:5] ? valid_512 : _GEN_512; // @[ICache.scala 68:{44,44}]
  wire  _GEN_514 = 10'h201 == req_r_addr[14:5] ? valid_513 : _GEN_513; // @[ICache.scala 68:{44,44}]
  wire  _GEN_515 = 10'h202 == req_r_addr[14:5] ? valid_514 : _GEN_514; // @[ICache.scala 68:{44,44}]
  wire  _GEN_516 = 10'h203 == req_r_addr[14:5] ? valid_515 : _GEN_515; // @[ICache.scala 68:{44,44}]
  wire  _GEN_517 = 10'h204 == req_r_addr[14:5] ? valid_516 : _GEN_516; // @[ICache.scala 68:{44,44}]
  wire  _GEN_518 = 10'h205 == req_r_addr[14:5] ? valid_517 : _GEN_517; // @[ICache.scala 68:{44,44}]
  wire  _GEN_519 = 10'h206 == req_r_addr[14:5] ? valid_518 : _GEN_518; // @[ICache.scala 68:{44,44}]
  wire  _GEN_520 = 10'h207 == req_r_addr[14:5] ? valid_519 : _GEN_519; // @[ICache.scala 68:{44,44}]
  wire  _GEN_521 = 10'h208 == req_r_addr[14:5] ? valid_520 : _GEN_520; // @[ICache.scala 68:{44,44}]
  wire  _GEN_522 = 10'h209 == req_r_addr[14:5] ? valid_521 : _GEN_521; // @[ICache.scala 68:{44,44}]
  wire  _GEN_523 = 10'h20a == req_r_addr[14:5] ? valid_522 : _GEN_522; // @[ICache.scala 68:{44,44}]
  wire  _GEN_524 = 10'h20b == req_r_addr[14:5] ? valid_523 : _GEN_523; // @[ICache.scala 68:{44,44}]
  wire  _GEN_525 = 10'h20c == req_r_addr[14:5] ? valid_524 : _GEN_524; // @[ICache.scala 68:{44,44}]
  wire  _GEN_526 = 10'h20d == req_r_addr[14:5] ? valid_525 : _GEN_525; // @[ICache.scala 68:{44,44}]
  wire  _GEN_527 = 10'h20e == req_r_addr[14:5] ? valid_526 : _GEN_526; // @[ICache.scala 68:{44,44}]
  wire  _GEN_528 = 10'h20f == req_r_addr[14:5] ? valid_527 : _GEN_527; // @[ICache.scala 68:{44,44}]
  wire  _GEN_529 = 10'h210 == req_r_addr[14:5] ? valid_528 : _GEN_528; // @[ICache.scala 68:{44,44}]
  wire  _GEN_530 = 10'h211 == req_r_addr[14:5] ? valid_529 : _GEN_529; // @[ICache.scala 68:{44,44}]
  wire  _GEN_531 = 10'h212 == req_r_addr[14:5] ? valid_530 : _GEN_530; // @[ICache.scala 68:{44,44}]
  wire  _GEN_532 = 10'h213 == req_r_addr[14:5] ? valid_531 : _GEN_531; // @[ICache.scala 68:{44,44}]
  wire  _GEN_533 = 10'h214 == req_r_addr[14:5] ? valid_532 : _GEN_532; // @[ICache.scala 68:{44,44}]
  wire  _GEN_534 = 10'h215 == req_r_addr[14:5] ? valid_533 : _GEN_533; // @[ICache.scala 68:{44,44}]
  wire  _GEN_535 = 10'h216 == req_r_addr[14:5] ? valid_534 : _GEN_534; // @[ICache.scala 68:{44,44}]
  wire  _GEN_536 = 10'h217 == req_r_addr[14:5] ? valid_535 : _GEN_535; // @[ICache.scala 68:{44,44}]
  wire  _GEN_537 = 10'h218 == req_r_addr[14:5] ? valid_536 : _GEN_536; // @[ICache.scala 68:{44,44}]
  wire  _GEN_538 = 10'h219 == req_r_addr[14:5] ? valid_537 : _GEN_537; // @[ICache.scala 68:{44,44}]
  wire  _GEN_539 = 10'h21a == req_r_addr[14:5] ? valid_538 : _GEN_538; // @[ICache.scala 68:{44,44}]
  wire  _GEN_540 = 10'h21b == req_r_addr[14:5] ? valid_539 : _GEN_539; // @[ICache.scala 68:{44,44}]
  wire  _GEN_541 = 10'h21c == req_r_addr[14:5] ? valid_540 : _GEN_540; // @[ICache.scala 68:{44,44}]
  wire  _GEN_542 = 10'h21d == req_r_addr[14:5] ? valid_541 : _GEN_541; // @[ICache.scala 68:{44,44}]
  wire  _GEN_543 = 10'h21e == req_r_addr[14:5] ? valid_542 : _GEN_542; // @[ICache.scala 68:{44,44}]
  wire  _GEN_544 = 10'h21f == req_r_addr[14:5] ? valid_543 : _GEN_543; // @[ICache.scala 68:{44,44}]
  wire  _GEN_545 = 10'h220 == req_r_addr[14:5] ? valid_544 : _GEN_544; // @[ICache.scala 68:{44,44}]
  wire  _GEN_546 = 10'h221 == req_r_addr[14:5] ? valid_545 : _GEN_545; // @[ICache.scala 68:{44,44}]
  wire  _GEN_547 = 10'h222 == req_r_addr[14:5] ? valid_546 : _GEN_546; // @[ICache.scala 68:{44,44}]
  wire  _GEN_548 = 10'h223 == req_r_addr[14:5] ? valid_547 : _GEN_547; // @[ICache.scala 68:{44,44}]
  wire  _GEN_549 = 10'h224 == req_r_addr[14:5] ? valid_548 : _GEN_548; // @[ICache.scala 68:{44,44}]
  wire  _GEN_550 = 10'h225 == req_r_addr[14:5] ? valid_549 : _GEN_549; // @[ICache.scala 68:{44,44}]
  wire  _GEN_551 = 10'h226 == req_r_addr[14:5] ? valid_550 : _GEN_550; // @[ICache.scala 68:{44,44}]
  wire  _GEN_552 = 10'h227 == req_r_addr[14:5] ? valid_551 : _GEN_551; // @[ICache.scala 68:{44,44}]
  wire  _GEN_553 = 10'h228 == req_r_addr[14:5] ? valid_552 : _GEN_552; // @[ICache.scala 68:{44,44}]
  wire  _GEN_554 = 10'h229 == req_r_addr[14:5] ? valid_553 : _GEN_553; // @[ICache.scala 68:{44,44}]
  wire  _GEN_555 = 10'h22a == req_r_addr[14:5] ? valid_554 : _GEN_554; // @[ICache.scala 68:{44,44}]
  wire  _GEN_556 = 10'h22b == req_r_addr[14:5] ? valid_555 : _GEN_555; // @[ICache.scala 68:{44,44}]
  wire  _GEN_557 = 10'h22c == req_r_addr[14:5] ? valid_556 : _GEN_556; // @[ICache.scala 68:{44,44}]
  wire  _GEN_558 = 10'h22d == req_r_addr[14:5] ? valid_557 : _GEN_557; // @[ICache.scala 68:{44,44}]
  wire  _GEN_559 = 10'h22e == req_r_addr[14:5] ? valid_558 : _GEN_558; // @[ICache.scala 68:{44,44}]
  wire  _GEN_560 = 10'h22f == req_r_addr[14:5] ? valid_559 : _GEN_559; // @[ICache.scala 68:{44,44}]
  wire  _GEN_561 = 10'h230 == req_r_addr[14:5] ? valid_560 : _GEN_560; // @[ICache.scala 68:{44,44}]
  wire  _GEN_562 = 10'h231 == req_r_addr[14:5] ? valid_561 : _GEN_561; // @[ICache.scala 68:{44,44}]
  wire  _GEN_563 = 10'h232 == req_r_addr[14:5] ? valid_562 : _GEN_562; // @[ICache.scala 68:{44,44}]
  wire  _GEN_564 = 10'h233 == req_r_addr[14:5] ? valid_563 : _GEN_563; // @[ICache.scala 68:{44,44}]
  wire  _GEN_565 = 10'h234 == req_r_addr[14:5] ? valid_564 : _GEN_564; // @[ICache.scala 68:{44,44}]
  wire  _GEN_566 = 10'h235 == req_r_addr[14:5] ? valid_565 : _GEN_565; // @[ICache.scala 68:{44,44}]
  wire  _GEN_567 = 10'h236 == req_r_addr[14:5] ? valid_566 : _GEN_566; // @[ICache.scala 68:{44,44}]
  wire  _GEN_568 = 10'h237 == req_r_addr[14:5] ? valid_567 : _GEN_567; // @[ICache.scala 68:{44,44}]
  wire  _GEN_569 = 10'h238 == req_r_addr[14:5] ? valid_568 : _GEN_568; // @[ICache.scala 68:{44,44}]
  wire  _GEN_570 = 10'h239 == req_r_addr[14:5] ? valid_569 : _GEN_569; // @[ICache.scala 68:{44,44}]
  wire  _GEN_571 = 10'h23a == req_r_addr[14:5] ? valid_570 : _GEN_570; // @[ICache.scala 68:{44,44}]
  wire  _GEN_572 = 10'h23b == req_r_addr[14:5] ? valid_571 : _GEN_571; // @[ICache.scala 68:{44,44}]
  wire  _GEN_573 = 10'h23c == req_r_addr[14:5] ? valid_572 : _GEN_572; // @[ICache.scala 68:{44,44}]
  wire  _GEN_574 = 10'h23d == req_r_addr[14:5] ? valid_573 : _GEN_573; // @[ICache.scala 68:{44,44}]
  wire  _GEN_575 = 10'h23e == req_r_addr[14:5] ? valid_574 : _GEN_574; // @[ICache.scala 68:{44,44}]
  wire  _GEN_576 = 10'h23f == req_r_addr[14:5] ? valid_575 : _GEN_575; // @[ICache.scala 68:{44,44}]
  wire  _GEN_577 = 10'h240 == req_r_addr[14:5] ? valid_576 : _GEN_576; // @[ICache.scala 68:{44,44}]
  wire  _GEN_578 = 10'h241 == req_r_addr[14:5] ? valid_577 : _GEN_577; // @[ICache.scala 68:{44,44}]
  wire  _GEN_579 = 10'h242 == req_r_addr[14:5] ? valid_578 : _GEN_578; // @[ICache.scala 68:{44,44}]
  wire  _GEN_580 = 10'h243 == req_r_addr[14:5] ? valid_579 : _GEN_579; // @[ICache.scala 68:{44,44}]
  wire  _GEN_581 = 10'h244 == req_r_addr[14:5] ? valid_580 : _GEN_580; // @[ICache.scala 68:{44,44}]
  wire  _GEN_582 = 10'h245 == req_r_addr[14:5] ? valid_581 : _GEN_581; // @[ICache.scala 68:{44,44}]
  wire  _GEN_583 = 10'h246 == req_r_addr[14:5] ? valid_582 : _GEN_582; // @[ICache.scala 68:{44,44}]
  wire  _GEN_584 = 10'h247 == req_r_addr[14:5] ? valid_583 : _GEN_583; // @[ICache.scala 68:{44,44}]
  wire  _GEN_585 = 10'h248 == req_r_addr[14:5] ? valid_584 : _GEN_584; // @[ICache.scala 68:{44,44}]
  wire  _GEN_586 = 10'h249 == req_r_addr[14:5] ? valid_585 : _GEN_585; // @[ICache.scala 68:{44,44}]
  wire  _GEN_587 = 10'h24a == req_r_addr[14:5] ? valid_586 : _GEN_586; // @[ICache.scala 68:{44,44}]
  wire  _GEN_588 = 10'h24b == req_r_addr[14:5] ? valid_587 : _GEN_587; // @[ICache.scala 68:{44,44}]
  wire  _GEN_589 = 10'h24c == req_r_addr[14:5] ? valid_588 : _GEN_588; // @[ICache.scala 68:{44,44}]
  wire  _GEN_590 = 10'h24d == req_r_addr[14:5] ? valid_589 : _GEN_589; // @[ICache.scala 68:{44,44}]
  wire  _GEN_591 = 10'h24e == req_r_addr[14:5] ? valid_590 : _GEN_590; // @[ICache.scala 68:{44,44}]
  wire  _GEN_592 = 10'h24f == req_r_addr[14:5] ? valid_591 : _GEN_591; // @[ICache.scala 68:{44,44}]
  wire  _GEN_593 = 10'h250 == req_r_addr[14:5] ? valid_592 : _GEN_592; // @[ICache.scala 68:{44,44}]
  wire  _GEN_594 = 10'h251 == req_r_addr[14:5] ? valid_593 : _GEN_593; // @[ICache.scala 68:{44,44}]
  wire  _GEN_595 = 10'h252 == req_r_addr[14:5] ? valid_594 : _GEN_594; // @[ICache.scala 68:{44,44}]
  wire  _GEN_596 = 10'h253 == req_r_addr[14:5] ? valid_595 : _GEN_595; // @[ICache.scala 68:{44,44}]
  wire  _GEN_597 = 10'h254 == req_r_addr[14:5] ? valid_596 : _GEN_596; // @[ICache.scala 68:{44,44}]
  wire  _GEN_598 = 10'h255 == req_r_addr[14:5] ? valid_597 : _GEN_597; // @[ICache.scala 68:{44,44}]
  wire  _GEN_599 = 10'h256 == req_r_addr[14:5] ? valid_598 : _GEN_598; // @[ICache.scala 68:{44,44}]
  wire  _GEN_600 = 10'h257 == req_r_addr[14:5] ? valid_599 : _GEN_599; // @[ICache.scala 68:{44,44}]
  wire  _GEN_601 = 10'h258 == req_r_addr[14:5] ? valid_600 : _GEN_600; // @[ICache.scala 68:{44,44}]
  wire  _GEN_602 = 10'h259 == req_r_addr[14:5] ? valid_601 : _GEN_601; // @[ICache.scala 68:{44,44}]
  wire  _GEN_603 = 10'h25a == req_r_addr[14:5] ? valid_602 : _GEN_602; // @[ICache.scala 68:{44,44}]
  wire  _GEN_604 = 10'h25b == req_r_addr[14:5] ? valid_603 : _GEN_603; // @[ICache.scala 68:{44,44}]
  wire  _GEN_605 = 10'h25c == req_r_addr[14:5] ? valid_604 : _GEN_604; // @[ICache.scala 68:{44,44}]
  wire  _GEN_606 = 10'h25d == req_r_addr[14:5] ? valid_605 : _GEN_605; // @[ICache.scala 68:{44,44}]
  wire  _GEN_607 = 10'h25e == req_r_addr[14:5] ? valid_606 : _GEN_606; // @[ICache.scala 68:{44,44}]
  wire  _GEN_608 = 10'h25f == req_r_addr[14:5] ? valid_607 : _GEN_607; // @[ICache.scala 68:{44,44}]
  wire  _GEN_609 = 10'h260 == req_r_addr[14:5] ? valid_608 : _GEN_608; // @[ICache.scala 68:{44,44}]
  wire  _GEN_610 = 10'h261 == req_r_addr[14:5] ? valid_609 : _GEN_609; // @[ICache.scala 68:{44,44}]
  wire  _GEN_611 = 10'h262 == req_r_addr[14:5] ? valid_610 : _GEN_610; // @[ICache.scala 68:{44,44}]
  wire  _GEN_612 = 10'h263 == req_r_addr[14:5] ? valid_611 : _GEN_611; // @[ICache.scala 68:{44,44}]
  wire  _GEN_613 = 10'h264 == req_r_addr[14:5] ? valid_612 : _GEN_612; // @[ICache.scala 68:{44,44}]
  wire  _GEN_614 = 10'h265 == req_r_addr[14:5] ? valid_613 : _GEN_613; // @[ICache.scala 68:{44,44}]
  wire  _GEN_615 = 10'h266 == req_r_addr[14:5] ? valid_614 : _GEN_614; // @[ICache.scala 68:{44,44}]
  wire  _GEN_616 = 10'h267 == req_r_addr[14:5] ? valid_615 : _GEN_615; // @[ICache.scala 68:{44,44}]
  wire  _GEN_617 = 10'h268 == req_r_addr[14:5] ? valid_616 : _GEN_616; // @[ICache.scala 68:{44,44}]
  wire  _GEN_618 = 10'h269 == req_r_addr[14:5] ? valid_617 : _GEN_617; // @[ICache.scala 68:{44,44}]
  wire  _GEN_619 = 10'h26a == req_r_addr[14:5] ? valid_618 : _GEN_618; // @[ICache.scala 68:{44,44}]
  wire  _GEN_620 = 10'h26b == req_r_addr[14:5] ? valid_619 : _GEN_619; // @[ICache.scala 68:{44,44}]
  wire  _GEN_621 = 10'h26c == req_r_addr[14:5] ? valid_620 : _GEN_620; // @[ICache.scala 68:{44,44}]
  wire  _GEN_622 = 10'h26d == req_r_addr[14:5] ? valid_621 : _GEN_621; // @[ICache.scala 68:{44,44}]
  wire  _GEN_623 = 10'h26e == req_r_addr[14:5] ? valid_622 : _GEN_622; // @[ICache.scala 68:{44,44}]
  wire  _GEN_624 = 10'h26f == req_r_addr[14:5] ? valid_623 : _GEN_623; // @[ICache.scala 68:{44,44}]
  wire  _GEN_625 = 10'h270 == req_r_addr[14:5] ? valid_624 : _GEN_624; // @[ICache.scala 68:{44,44}]
  wire  _GEN_626 = 10'h271 == req_r_addr[14:5] ? valid_625 : _GEN_625; // @[ICache.scala 68:{44,44}]
  wire  _GEN_627 = 10'h272 == req_r_addr[14:5] ? valid_626 : _GEN_626; // @[ICache.scala 68:{44,44}]
  wire  _GEN_628 = 10'h273 == req_r_addr[14:5] ? valid_627 : _GEN_627; // @[ICache.scala 68:{44,44}]
  wire  _GEN_629 = 10'h274 == req_r_addr[14:5] ? valid_628 : _GEN_628; // @[ICache.scala 68:{44,44}]
  wire  _GEN_630 = 10'h275 == req_r_addr[14:5] ? valid_629 : _GEN_629; // @[ICache.scala 68:{44,44}]
  wire  _GEN_631 = 10'h276 == req_r_addr[14:5] ? valid_630 : _GEN_630; // @[ICache.scala 68:{44,44}]
  wire  _GEN_632 = 10'h277 == req_r_addr[14:5] ? valid_631 : _GEN_631; // @[ICache.scala 68:{44,44}]
  wire  _GEN_633 = 10'h278 == req_r_addr[14:5] ? valid_632 : _GEN_632; // @[ICache.scala 68:{44,44}]
  wire  _GEN_634 = 10'h279 == req_r_addr[14:5] ? valid_633 : _GEN_633; // @[ICache.scala 68:{44,44}]
  wire  _GEN_635 = 10'h27a == req_r_addr[14:5] ? valid_634 : _GEN_634; // @[ICache.scala 68:{44,44}]
  wire  _GEN_636 = 10'h27b == req_r_addr[14:5] ? valid_635 : _GEN_635; // @[ICache.scala 68:{44,44}]
  wire  _GEN_637 = 10'h27c == req_r_addr[14:5] ? valid_636 : _GEN_636; // @[ICache.scala 68:{44,44}]
  wire  _GEN_638 = 10'h27d == req_r_addr[14:5] ? valid_637 : _GEN_637; // @[ICache.scala 68:{44,44}]
  wire  _GEN_639 = 10'h27e == req_r_addr[14:5] ? valid_638 : _GEN_638; // @[ICache.scala 68:{44,44}]
  wire  _GEN_640 = 10'h27f == req_r_addr[14:5] ? valid_639 : _GEN_639; // @[ICache.scala 68:{44,44}]
  wire  _GEN_641 = 10'h280 == req_r_addr[14:5] ? valid_640 : _GEN_640; // @[ICache.scala 68:{44,44}]
  wire  _GEN_642 = 10'h281 == req_r_addr[14:5] ? valid_641 : _GEN_641; // @[ICache.scala 68:{44,44}]
  wire  _GEN_643 = 10'h282 == req_r_addr[14:5] ? valid_642 : _GEN_642; // @[ICache.scala 68:{44,44}]
  wire  _GEN_644 = 10'h283 == req_r_addr[14:5] ? valid_643 : _GEN_643; // @[ICache.scala 68:{44,44}]
  wire  _GEN_645 = 10'h284 == req_r_addr[14:5] ? valid_644 : _GEN_644; // @[ICache.scala 68:{44,44}]
  wire  _GEN_646 = 10'h285 == req_r_addr[14:5] ? valid_645 : _GEN_645; // @[ICache.scala 68:{44,44}]
  wire  _GEN_647 = 10'h286 == req_r_addr[14:5] ? valid_646 : _GEN_646; // @[ICache.scala 68:{44,44}]
  wire  _GEN_648 = 10'h287 == req_r_addr[14:5] ? valid_647 : _GEN_647; // @[ICache.scala 68:{44,44}]
  wire  _GEN_649 = 10'h288 == req_r_addr[14:5] ? valid_648 : _GEN_648; // @[ICache.scala 68:{44,44}]
  wire  _GEN_650 = 10'h289 == req_r_addr[14:5] ? valid_649 : _GEN_649; // @[ICache.scala 68:{44,44}]
  wire  _GEN_651 = 10'h28a == req_r_addr[14:5] ? valid_650 : _GEN_650; // @[ICache.scala 68:{44,44}]
  wire  _GEN_652 = 10'h28b == req_r_addr[14:5] ? valid_651 : _GEN_651; // @[ICache.scala 68:{44,44}]
  wire  _GEN_653 = 10'h28c == req_r_addr[14:5] ? valid_652 : _GEN_652; // @[ICache.scala 68:{44,44}]
  wire  _GEN_654 = 10'h28d == req_r_addr[14:5] ? valid_653 : _GEN_653; // @[ICache.scala 68:{44,44}]
  wire  _GEN_655 = 10'h28e == req_r_addr[14:5] ? valid_654 : _GEN_654; // @[ICache.scala 68:{44,44}]
  wire  _GEN_656 = 10'h28f == req_r_addr[14:5] ? valid_655 : _GEN_655; // @[ICache.scala 68:{44,44}]
  wire  _GEN_657 = 10'h290 == req_r_addr[14:5] ? valid_656 : _GEN_656; // @[ICache.scala 68:{44,44}]
  wire  _GEN_658 = 10'h291 == req_r_addr[14:5] ? valid_657 : _GEN_657; // @[ICache.scala 68:{44,44}]
  wire  _GEN_659 = 10'h292 == req_r_addr[14:5] ? valid_658 : _GEN_658; // @[ICache.scala 68:{44,44}]
  wire  _GEN_660 = 10'h293 == req_r_addr[14:5] ? valid_659 : _GEN_659; // @[ICache.scala 68:{44,44}]
  wire  _GEN_661 = 10'h294 == req_r_addr[14:5] ? valid_660 : _GEN_660; // @[ICache.scala 68:{44,44}]
  wire  _GEN_662 = 10'h295 == req_r_addr[14:5] ? valid_661 : _GEN_661; // @[ICache.scala 68:{44,44}]
  wire  _GEN_663 = 10'h296 == req_r_addr[14:5] ? valid_662 : _GEN_662; // @[ICache.scala 68:{44,44}]
  wire  _GEN_664 = 10'h297 == req_r_addr[14:5] ? valid_663 : _GEN_663; // @[ICache.scala 68:{44,44}]
  wire  _GEN_665 = 10'h298 == req_r_addr[14:5] ? valid_664 : _GEN_664; // @[ICache.scala 68:{44,44}]
  wire  _GEN_666 = 10'h299 == req_r_addr[14:5] ? valid_665 : _GEN_665; // @[ICache.scala 68:{44,44}]
  wire  _GEN_667 = 10'h29a == req_r_addr[14:5] ? valid_666 : _GEN_666; // @[ICache.scala 68:{44,44}]
  wire  _GEN_668 = 10'h29b == req_r_addr[14:5] ? valid_667 : _GEN_667; // @[ICache.scala 68:{44,44}]
  wire  _GEN_669 = 10'h29c == req_r_addr[14:5] ? valid_668 : _GEN_668; // @[ICache.scala 68:{44,44}]
  wire  _GEN_670 = 10'h29d == req_r_addr[14:5] ? valid_669 : _GEN_669; // @[ICache.scala 68:{44,44}]
  wire  _GEN_671 = 10'h29e == req_r_addr[14:5] ? valid_670 : _GEN_670; // @[ICache.scala 68:{44,44}]
  wire  _GEN_672 = 10'h29f == req_r_addr[14:5] ? valid_671 : _GEN_671; // @[ICache.scala 68:{44,44}]
  wire  _GEN_673 = 10'h2a0 == req_r_addr[14:5] ? valid_672 : _GEN_672; // @[ICache.scala 68:{44,44}]
  wire  _GEN_674 = 10'h2a1 == req_r_addr[14:5] ? valid_673 : _GEN_673; // @[ICache.scala 68:{44,44}]
  wire  _GEN_675 = 10'h2a2 == req_r_addr[14:5] ? valid_674 : _GEN_674; // @[ICache.scala 68:{44,44}]
  wire  _GEN_676 = 10'h2a3 == req_r_addr[14:5] ? valid_675 : _GEN_675; // @[ICache.scala 68:{44,44}]
  wire  _GEN_677 = 10'h2a4 == req_r_addr[14:5] ? valid_676 : _GEN_676; // @[ICache.scala 68:{44,44}]
  wire  _GEN_678 = 10'h2a5 == req_r_addr[14:5] ? valid_677 : _GEN_677; // @[ICache.scala 68:{44,44}]
  wire  _GEN_679 = 10'h2a6 == req_r_addr[14:5] ? valid_678 : _GEN_678; // @[ICache.scala 68:{44,44}]
  wire  _GEN_680 = 10'h2a7 == req_r_addr[14:5] ? valid_679 : _GEN_679; // @[ICache.scala 68:{44,44}]
  wire  _GEN_681 = 10'h2a8 == req_r_addr[14:5] ? valid_680 : _GEN_680; // @[ICache.scala 68:{44,44}]
  wire  _GEN_682 = 10'h2a9 == req_r_addr[14:5] ? valid_681 : _GEN_681; // @[ICache.scala 68:{44,44}]
  wire  _GEN_683 = 10'h2aa == req_r_addr[14:5] ? valid_682 : _GEN_682; // @[ICache.scala 68:{44,44}]
  wire  _GEN_684 = 10'h2ab == req_r_addr[14:5] ? valid_683 : _GEN_683; // @[ICache.scala 68:{44,44}]
  wire  _GEN_685 = 10'h2ac == req_r_addr[14:5] ? valid_684 : _GEN_684; // @[ICache.scala 68:{44,44}]
  wire  _GEN_686 = 10'h2ad == req_r_addr[14:5] ? valid_685 : _GEN_685; // @[ICache.scala 68:{44,44}]
  wire  _GEN_687 = 10'h2ae == req_r_addr[14:5] ? valid_686 : _GEN_686; // @[ICache.scala 68:{44,44}]
  wire  _GEN_688 = 10'h2af == req_r_addr[14:5] ? valid_687 : _GEN_687; // @[ICache.scala 68:{44,44}]
  wire  _GEN_689 = 10'h2b0 == req_r_addr[14:5] ? valid_688 : _GEN_688; // @[ICache.scala 68:{44,44}]
  wire  _GEN_690 = 10'h2b1 == req_r_addr[14:5] ? valid_689 : _GEN_689; // @[ICache.scala 68:{44,44}]
  wire  _GEN_691 = 10'h2b2 == req_r_addr[14:5] ? valid_690 : _GEN_690; // @[ICache.scala 68:{44,44}]
  wire  _GEN_692 = 10'h2b3 == req_r_addr[14:5] ? valid_691 : _GEN_691; // @[ICache.scala 68:{44,44}]
  wire  _GEN_693 = 10'h2b4 == req_r_addr[14:5] ? valid_692 : _GEN_692; // @[ICache.scala 68:{44,44}]
  wire  _GEN_694 = 10'h2b5 == req_r_addr[14:5] ? valid_693 : _GEN_693; // @[ICache.scala 68:{44,44}]
  wire  _GEN_695 = 10'h2b6 == req_r_addr[14:5] ? valid_694 : _GEN_694; // @[ICache.scala 68:{44,44}]
  wire  _GEN_696 = 10'h2b7 == req_r_addr[14:5] ? valid_695 : _GEN_695; // @[ICache.scala 68:{44,44}]
  wire  _GEN_697 = 10'h2b8 == req_r_addr[14:5] ? valid_696 : _GEN_696; // @[ICache.scala 68:{44,44}]
  wire  _GEN_698 = 10'h2b9 == req_r_addr[14:5] ? valid_697 : _GEN_697; // @[ICache.scala 68:{44,44}]
  wire  _GEN_699 = 10'h2ba == req_r_addr[14:5] ? valid_698 : _GEN_698; // @[ICache.scala 68:{44,44}]
  wire  _GEN_700 = 10'h2bb == req_r_addr[14:5] ? valid_699 : _GEN_699; // @[ICache.scala 68:{44,44}]
  wire  _GEN_701 = 10'h2bc == req_r_addr[14:5] ? valid_700 : _GEN_700; // @[ICache.scala 68:{44,44}]
  wire  _GEN_702 = 10'h2bd == req_r_addr[14:5] ? valid_701 : _GEN_701; // @[ICache.scala 68:{44,44}]
  wire  _GEN_703 = 10'h2be == req_r_addr[14:5] ? valid_702 : _GEN_702; // @[ICache.scala 68:{44,44}]
  wire  _GEN_704 = 10'h2bf == req_r_addr[14:5] ? valid_703 : _GEN_703; // @[ICache.scala 68:{44,44}]
  wire  _GEN_705 = 10'h2c0 == req_r_addr[14:5] ? valid_704 : _GEN_704; // @[ICache.scala 68:{44,44}]
  wire  _GEN_706 = 10'h2c1 == req_r_addr[14:5] ? valid_705 : _GEN_705; // @[ICache.scala 68:{44,44}]
  wire  _GEN_707 = 10'h2c2 == req_r_addr[14:5] ? valid_706 : _GEN_706; // @[ICache.scala 68:{44,44}]
  wire  _GEN_708 = 10'h2c3 == req_r_addr[14:5] ? valid_707 : _GEN_707; // @[ICache.scala 68:{44,44}]
  wire  _GEN_709 = 10'h2c4 == req_r_addr[14:5] ? valid_708 : _GEN_708; // @[ICache.scala 68:{44,44}]
  wire  _GEN_710 = 10'h2c5 == req_r_addr[14:5] ? valid_709 : _GEN_709; // @[ICache.scala 68:{44,44}]
  wire  _GEN_711 = 10'h2c6 == req_r_addr[14:5] ? valid_710 : _GEN_710; // @[ICache.scala 68:{44,44}]
  wire  _GEN_712 = 10'h2c7 == req_r_addr[14:5] ? valid_711 : _GEN_711; // @[ICache.scala 68:{44,44}]
  wire  _GEN_713 = 10'h2c8 == req_r_addr[14:5] ? valid_712 : _GEN_712; // @[ICache.scala 68:{44,44}]
  wire  _GEN_714 = 10'h2c9 == req_r_addr[14:5] ? valid_713 : _GEN_713; // @[ICache.scala 68:{44,44}]
  wire  _GEN_715 = 10'h2ca == req_r_addr[14:5] ? valid_714 : _GEN_714; // @[ICache.scala 68:{44,44}]
  wire  _GEN_716 = 10'h2cb == req_r_addr[14:5] ? valid_715 : _GEN_715; // @[ICache.scala 68:{44,44}]
  wire  _GEN_717 = 10'h2cc == req_r_addr[14:5] ? valid_716 : _GEN_716; // @[ICache.scala 68:{44,44}]
  wire  _GEN_718 = 10'h2cd == req_r_addr[14:5] ? valid_717 : _GEN_717; // @[ICache.scala 68:{44,44}]
  wire  _GEN_719 = 10'h2ce == req_r_addr[14:5] ? valid_718 : _GEN_718; // @[ICache.scala 68:{44,44}]
  wire  _GEN_720 = 10'h2cf == req_r_addr[14:5] ? valid_719 : _GEN_719; // @[ICache.scala 68:{44,44}]
  wire  _GEN_721 = 10'h2d0 == req_r_addr[14:5] ? valid_720 : _GEN_720; // @[ICache.scala 68:{44,44}]
  wire  _GEN_722 = 10'h2d1 == req_r_addr[14:5] ? valid_721 : _GEN_721; // @[ICache.scala 68:{44,44}]
  wire  _GEN_723 = 10'h2d2 == req_r_addr[14:5] ? valid_722 : _GEN_722; // @[ICache.scala 68:{44,44}]
  wire  _GEN_724 = 10'h2d3 == req_r_addr[14:5] ? valid_723 : _GEN_723; // @[ICache.scala 68:{44,44}]
  wire  _GEN_725 = 10'h2d4 == req_r_addr[14:5] ? valid_724 : _GEN_724; // @[ICache.scala 68:{44,44}]
  wire  _GEN_726 = 10'h2d5 == req_r_addr[14:5] ? valid_725 : _GEN_725; // @[ICache.scala 68:{44,44}]
  wire  _GEN_727 = 10'h2d6 == req_r_addr[14:5] ? valid_726 : _GEN_726; // @[ICache.scala 68:{44,44}]
  wire  _GEN_728 = 10'h2d7 == req_r_addr[14:5] ? valid_727 : _GEN_727; // @[ICache.scala 68:{44,44}]
  wire  _GEN_729 = 10'h2d8 == req_r_addr[14:5] ? valid_728 : _GEN_728; // @[ICache.scala 68:{44,44}]
  wire  _GEN_730 = 10'h2d9 == req_r_addr[14:5] ? valid_729 : _GEN_729; // @[ICache.scala 68:{44,44}]
  wire  _GEN_731 = 10'h2da == req_r_addr[14:5] ? valid_730 : _GEN_730; // @[ICache.scala 68:{44,44}]
  wire  _GEN_732 = 10'h2db == req_r_addr[14:5] ? valid_731 : _GEN_731; // @[ICache.scala 68:{44,44}]
  wire  _GEN_733 = 10'h2dc == req_r_addr[14:5] ? valid_732 : _GEN_732; // @[ICache.scala 68:{44,44}]
  wire  _GEN_734 = 10'h2dd == req_r_addr[14:5] ? valid_733 : _GEN_733; // @[ICache.scala 68:{44,44}]
  wire  _GEN_735 = 10'h2de == req_r_addr[14:5] ? valid_734 : _GEN_734; // @[ICache.scala 68:{44,44}]
  wire  _GEN_736 = 10'h2df == req_r_addr[14:5] ? valid_735 : _GEN_735; // @[ICache.scala 68:{44,44}]
  wire  _GEN_737 = 10'h2e0 == req_r_addr[14:5] ? valid_736 : _GEN_736; // @[ICache.scala 68:{44,44}]
  wire  _GEN_738 = 10'h2e1 == req_r_addr[14:5] ? valid_737 : _GEN_737; // @[ICache.scala 68:{44,44}]
  wire  _GEN_739 = 10'h2e2 == req_r_addr[14:5] ? valid_738 : _GEN_738; // @[ICache.scala 68:{44,44}]
  wire  _GEN_740 = 10'h2e3 == req_r_addr[14:5] ? valid_739 : _GEN_739; // @[ICache.scala 68:{44,44}]
  wire  _GEN_741 = 10'h2e4 == req_r_addr[14:5] ? valid_740 : _GEN_740; // @[ICache.scala 68:{44,44}]
  wire  _GEN_742 = 10'h2e5 == req_r_addr[14:5] ? valid_741 : _GEN_741; // @[ICache.scala 68:{44,44}]
  wire  _GEN_743 = 10'h2e6 == req_r_addr[14:5] ? valid_742 : _GEN_742; // @[ICache.scala 68:{44,44}]
  wire  _GEN_744 = 10'h2e7 == req_r_addr[14:5] ? valid_743 : _GEN_743; // @[ICache.scala 68:{44,44}]
  wire  _GEN_745 = 10'h2e8 == req_r_addr[14:5] ? valid_744 : _GEN_744; // @[ICache.scala 68:{44,44}]
  wire  _GEN_746 = 10'h2e9 == req_r_addr[14:5] ? valid_745 : _GEN_745; // @[ICache.scala 68:{44,44}]
  wire  _GEN_747 = 10'h2ea == req_r_addr[14:5] ? valid_746 : _GEN_746; // @[ICache.scala 68:{44,44}]
  wire  _GEN_748 = 10'h2eb == req_r_addr[14:5] ? valid_747 : _GEN_747; // @[ICache.scala 68:{44,44}]
  wire  _GEN_749 = 10'h2ec == req_r_addr[14:5] ? valid_748 : _GEN_748; // @[ICache.scala 68:{44,44}]
  wire  _GEN_750 = 10'h2ed == req_r_addr[14:5] ? valid_749 : _GEN_749; // @[ICache.scala 68:{44,44}]
  wire  _GEN_751 = 10'h2ee == req_r_addr[14:5] ? valid_750 : _GEN_750; // @[ICache.scala 68:{44,44}]
  wire  _GEN_752 = 10'h2ef == req_r_addr[14:5] ? valid_751 : _GEN_751; // @[ICache.scala 68:{44,44}]
  wire  _GEN_753 = 10'h2f0 == req_r_addr[14:5] ? valid_752 : _GEN_752; // @[ICache.scala 68:{44,44}]
  wire  _GEN_754 = 10'h2f1 == req_r_addr[14:5] ? valid_753 : _GEN_753; // @[ICache.scala 68:{44,44}]
  wire  _GEN_755 = 10'h2f2 == req_r_addr[14:5] ? valid_754 : _GEN_754; // @[ICache.scala 68:{44,44}]
  wire  _GEN_756 = 10'h2f3 == req_r_addr[14:5] ? valid_755 : _GEN_755; // @[ICache.scala 68:{44,44}]
  wire  _GEN_757 = 10'h2f4 == req_r_addr[14:5] ? valid_756 : _GEN_756; // @[ICache.scala 68:{44,44}]
  wire  _GEN_758 = 10'h2f5 == req_r_addr[14:5] ? valid_757 : _GEN_757; // @[ICache.scala 68:{44,44}]
  wire  _GEN_759 = 10'h2f6 == req_r_addr[14:5] ? valid_758 : _GEN_758; // @[ICache.scala 68:{44,44}]
  wire  _GEN_760 = 10'h2f7 == req_r_addr[14:5] ? valid_759 : _GEN_759; // @[ICache.scala 68:{44,44}]
  wire  _GEN_761 = 10'h2f8 == req_r_addr[14:5] ? valid_760 : _GEN_760; // @[ICache.scala 68:{44,44}]
  wire  _GEN_762 = 10'h2f9 == req_r_addr[14:5] ? valid_761 : _GEN_761; // @[ICache.scala 68:{44,44}]
  wire  _GEN_763 = 10'h2fa == req_r_addr[14:5] ? valid_762 : _GEN_762; // @[ICache.scala 68:{44,44}]
  wire  _GEN_764 = 10'h2fb == req_r_addr[14:5] ? valid_763 : _GEN_763; // @[ICache.scala 68:{44,44}]
  wire  _GEN_765 = 10'h2fc == req_r_addr[14:5] ? valid_764 : _GEN_764; // @[ICache.scala 68:{44,44}]
  wire  _GEN_766 = 10'h2fd == req_r_addr[14:5] ? valid_765 : _GEN_765; // @[ICache.scala 68:{44,44}]
  wire  _GEN_767 = 10'h2fe == req_r_addr[14:5] ? valid_766 : _GEN_766; // @[ICache.scala 68:{44,44}]
  wire  _GEN_768 = 10'h2ff == req_r_addr[14:5] ? valid_767 : _GEN_767; // @[ICache.scala 68:{44,44}]
  wire  _GEN_769 = 10'h300 == req_r_addr[14:5] ? valid_768 : _GEN_768; // @[ICache.scala 68:{44,44}]
  wire  _GEN_770 = 10'h301 == req_r_addr[14:5] ? valid_769 : _GEN_769; // @[ICache.scala 68:{44,44}]
  wire  _GEN_771 = 10'h302 == req_r_addr[14:5] ? valid_770 : _GEN_770; // @[ICache.scala 68:{44,44}]
  wire  _GEN_772 = 10'h303 == req_r_addr[14:5] ? valid_771 : _GEN_771; // @[ICache.scala 68:{44,44}]
  wire  _GEN_773 = 10'h304 == req_r_addr[14:5] ? valid_772 : _GEN_772; // @[ICache.scala 68:{44,44}]
  wire  _GEN_774 = 10'h305 == req_r_addr[14:5] ? valid_773 : _GEN_773; // @[ICache.scala 68:{44,44}]
  wire  _GEN_775 = 10'h306 == req_r_addr[14:5] ? valid_774 : _GEN_774; // @[ICache.scala 68:{44,44}]
  wire  _GEN_776 = 10'h307 == req_r_addr[14:5] ? valid_775 : _GEN_775; // @[ICache.scala 68:{44,44}]
  wire  _GEN_777 = 10'h308 == req_r_addr[14:5] ? valid_776 : _GEN_776; // @[ICache.scala 68:{44,44}]
  wire  _GEN_778 = 10'h309 == req_r_addr[14:5] ? valid_777 : _GEN_777; // @[ICache.scala 68:{44,44}]
  wire  _GEN_779 = 10'h30a == req_r_addr[14:5] ? valid_778 : _GEN_778; // @[ICache.scala 68:{44,44}]
  wire  _GEN_780 = 10'h30b == req_r_addr[14:5] ? valid_779 : _GEN_779; // @[ICache.scala 68:{44,44}]
  wire  _GEN_781 = 10'h30c == req_r_addr[14:5] ? valid_780 : _GEN_780; // @[ICache.scala 68:{44,44}]
  wire  _GEN_782 = 10'h30d == req_r_addr[14:5] ? valid_781 : _GEN_781; // @[ICache.scala 68:{44,44}]
  wire  _GEN_783 = 10'h30e == req_r_addr[14:5] ? valid_782 : _GEN_782; // @[ICache.scala 68:{44,44}]
  wire  _GEN_784 = 10'h30f == req_r_addr[14:5] ? valid_783 : _GEN_783; // @[ICache.scala 68:{44,44}]
  wire  _GEN_785 = 10'h310 == req_r_addr[14:5] ? valid_784 : _GEN_784; // @[ICache.scala 68:{44,44}]
  wire  _GEN_786 = 10'h311 == req_r_addr[14:5] ? valid_785 : _GEN_785; // @[ICache.scala 68:{44,44}]
  wire  _GEN_787 = 10'h312 == req_r_addr[14:5] ? valid_786 : _GEN_786; // @[ICache.scala 68:{44,44}]
  wire  _GEN_788 = 10'h313 == req_r_addr[14:5] ? valid_787 : _GEN_787; // @[ICache.scala 68:{44,44}]
  wire  _GEN_789 = 10'h314 == req_r_addr[14:5] ? valid_788 : _GEN_788; // @[ICache.scala 68:{44,44}]
  wire  _GEN_790 = 10'h315 == req_r_addr[14:5] ? valid_789 : _GEN_789; // @[ICache.scala 68:{44,44}]
  wire  _GEN_791 = 10'h316 == req_r_addr[14:5] ? valid_790 : _GEN_790; // @[ICache.scala 68:{44,44}]
  wire  _GEN_792 = 10'h317 == req_r_addr[14:5] ? valid_791 : _GEN_791; // @[ICache.scala 68:{44,44}]
  wire  _GEN_793 = 10'h318 == req_r_addr[14:5] ? valid_792 : _GEN_792; // @[ICache.scala 68:{44,44}]
  wire  _GEN_794 = 10'h319 == req_r_addr[14:5] ? valid_793 : _GEN_793; // @[ICache.scala 68:{44,44}]
  wire  _GEN_795 = 10'h31a == req_r_addr[14:5] ? valid_794 : _GEN_794; // @[ICache.scala 68:{44,44}]
  wire  _GEN_796 = 10'h31b == req_r_addr[14:5] ? valid_795 : _GEN_795; // @[ICache.scala 68:{44,44}]
  wire  _GEN_797 = 10'h31c == req_r_addr[14:5] ? valid_796 : _GEN_796; // @[ICache.scala 68:{44,44}]
  wire  _GEN_798 = 10'h31d == req_r_addr[14:5] ? valid_797 : _GEN_797; // @[ICache.scala 68:{44,44}]
  wire  _GEN_799 = 10'h31e == req_r_addr[14:5] ? valid_798 : _GEN_798; // @[ICache.scala 68:{44,44}]
  wire  _GEN_800 = 10'h31f == req_r_addr[14:5] ? valid_799 : _GEN_799; // @[ICache.scala 68:{44,44}]
  wire  _GEN_801 = 10'h320 == req_r_addr[14:5] ? valid_800 : _GEN_800; // @[ICache.scala 68:{44,44}]
  wire  _GEN_802 = 10'h321 == req_r_addr[14:5] ? valid_801 : _GEN_801; // @[ICache.scala 68:{44,44}]
  wire  _GEN_803 = 10'h322 == req_r_addr[14:5] ? valid_802 : _GEN_802; // @[ICache.scala 68:{44,44}]
  wire  _GEN_804 = 10'h323 == req_r_addr[14:5] ? valid_803 : _GEN_803; // @[ICache.scala 68:{44,44}]
  wire  _GEN_805 = 10'h324 == req_r_addr[14:5] ? valid_804 : _GEN_804; // @[ICache.scala 68:{44,44}]
  wire  _GEN_806 = 10'h325 == req_r_addr[14:5] ? valid_805 : _GEN_805; // @[ICache.scala 68:{44,44}]
  wire  _GEN_807 = 10'h326 == req_r_addr[14:5] ? valid_806 : _GEN_806; // @[ICache.scala 68:{44,44}]
  wire  _GEN_808 = 10'h327 == req_r_addr[14:5] ? valid_807 : _GEN_807; // @[ICache.scala 68:{44,44}]
  wire  _GEN_809 = 10'h328 == req_r_addr[14:5] ? valid_808 : _GEN_808; // @[ICache.scala 68:{44,44}]
  wire  _GEN_810 = 10'h329 == req_r_addr[14:5] ? valid_809 : _GEN_809; // @[ICache.scala 68:{44,44}]
  wire  _GEN_811 = 10'h32a == req_r_addr[14:5] ? valid_810 : _GEN_810; // @[ICache.scala 68:{44,44}]
  wire  _GEN_812 = 10'h32b == req_r_addr[14:5] ? valid_811 : _GEN_811; // @[ICache.scala 68:{44,44}]
  wire  _GEN_813 = 10'h32c == req_r_addr[14:5] ? valid_812 : _GEN_812; // @[ICache.scala 68:{44,44}]
  wire  _GEN_814 = 10'h32d == req_r_addr[14:5] ? valid_813 : _GEN_813; // @[ICache.scala 68:{44,44}]
  wire  _GEN_815 = 10'h32e == req_r_addr[14:5] ? valid_814 : _GEN_814; // @[ICache.scala 68:{44,44}]
  wire  _GEN_816 = 10'h32f == req_r_addr[14:5] ? valid_815 : _GEN_815; // @[ICache.scala 68:{44,44}]
  wire  _GEN_817 = 10'h330 == req_r_addr[14:5] ? valid_816 : _GEN_816; // @[ICache.scala 68:{44,44}]
  wire  _GEN_818 = 10'h331 == req_r_addr[14:5] ? valid_817 : _GEN_817; // @[ICache.scala 68:{44,44}]
  wire  _GEN_819 = 10'h332 == req_r_addr[14:5] ? valid_818 : _GEN_818; // @[ICache.scala 68:{44,44}]
  wire  _GEN_820 = 10'h333 == req_r_addr[14:5] ? valid_819 : _GEN_819; // @[ICache.scala 68:{44,44}]
  wire  _GEN_821 = 10'h334 == req_r_addr[14:5] ? valid_820 : _GEN_820; // @[ICache.scala 68:{44,44}]
  wire  _GEN_822 = 10'h335 == req_r_addr[14:5] ? valid_821 : _GEN_821; // @[ICache.scala 68:{44,44}]
  wire  _GEN_823 = 10'h336 == req_r_addr[14:5] ? valid_822 : _GEN_822; // @[ICache.scala 68:{44,44}]
  wire  _GEN_824 = 10'h337 == req_r_addr[14:5] ? valid_823 : _GEN_823; // @[ICache.scala 68:{44,44}]
  wire  _GEN_825 = 10'h338 == req_r_addr[14:5] ? valid_824 : _GEN_824; // @[ICache.scala 68:{44,44}]
  wire  _GEN_826 = 10'h339 == req_r_addr[14:5] ? valid_825 : _GEN_825; // @[ICache.scala 68:{44,44}]
  wire  _GEN_827 = 10'h33a == req_r_addr[14:5] ? valid_826 : _GEN_826; // @[ICache.scala 68:{44,44}]
  wire  _GEN_828 = 10'h33b == req_r_addr[14:5] ? valid_827 : _GEN_827; // @[ICache.scala 68:{44,44}]
  wire  _GEN_829 = 10'h33c == req_r_addr[14:5] ? valid_828 : _GEN_828; // @[ICache.scala 68:{44,44}]
  wire  _GEN_830 = 10'h33d == req_r_addr[14:5] ? valid_829 : _GEN_829; // @[ICache.scala 68:{44,44}]
  wire  _GEN_831 = 10'h33e == req_r_addr[14:5] ? valid_830 : _GEN_830; // @[ICache.scala 68:{44,44}]
  wire  _GEN_832 = 10'h33f == req_r_addr[14:5] ? valid_831 : _GEN_831; // @[ICache.scala 68:{44,44}]
  wire  _GEN_833 = 10'h340 == req_r_addr[14:5] ? valid_832 : _GEN_832; // @[ICache.scala 68:{44,44}]
  wire  _GEN_834 = 10'h341 == req_r_addr[14:5] ? valid_833 : _GEN_833; // @[ICache.scala 68:{44,44}]
  wire  _GEN_835 = 10'h342 == req_r_addr[14:5] ? valid_834 : _GEN_834; // @[ICache.scala 68:{44,44}]
  wire  _GEN_836 = 10'h343 == req_r_addr[14:5] ? valid_835 : _GEN_835; // @[ICache.scala 68:{44,44}]
  wire  _GEN_837 = 10'h344 == req_r_addr[14:5] ? valid_836 : _GEN_836; // @[ICache.scala 68:{44,44}]
  wire  _GEN_838 = 10'h345 == req_r_addr[14:5] ? valid_837 : _GEN_837; // @[ICache.scala 68:{44,44}]
  wire  _GEN_839 = 10'h346 == req_r_addr[14:5] ? valid_838 : _GEN_838; // @[ICache.scala 68:{44,44}]
  wire  _GEN_840 = 10'h347 == req_r_addr[14:5] ? valid_839 : _GEN_839; // @[ICache.scala 68:{44,44}]
  wire  _GEN_841 = 10'h348 == req_r_addr[14:5] ? valid_840 : _GEN_840; // @[ICache.scala 68:{44,44}]
  wire  _GEN_842 = 10'h349 == req_r_addr[14:5] ? valid_841 : _GEN_841; // @[ICache.scala 68:{44,44}]
  wire  _GEN_843 = 10'h34a == req_r_addr[14:5] ? valid_842 : _GEN_842; // @[ICache.scala 68:{44,44}]
  wire  _GEN_844 = 10'h34b == req_r_addr[14:5] ? valid_843 : _GEN_843; // @[ICache.scala 68:{44,44}]
  wire  _GEN_845 = 10'h34c == req_r_addr[14:5] ? valid_844 : _GEN_844; // @[ICache.scala 68:{44,44}]
  wire  _GEN_846 = 10'h34d == req_r_addr[14:5] ? valid_845 : _GEN_845; // @[ICache.scala 68:{44,44}]
  wire  _GEN_847 = 10'h34e == req_r_addr[14:5] ? valid_846 : _GEN_846; // @[ICache.scala 68:{44,44}]
  wire  _GEN_848 = 10'h34f == req_r_addr[14:5] ? valid_847 : _GEN_847; // @[ICache.scala 68:{44,44}]
  wire  _GEN_849 = 10'h350 == req_r_addr[14:5] ? valid_848 : _GEN_848; // @[ICache.scala 68:{44,44}]
  wire  _GEN_850 = 10'h351 == req_r_addr[14:5] ? valid_849 : _GEN_849; // @[ICache.scala 68:{44,44}]
  wire  _GEN_851 = 10'h352 == req_r_addr[14:5] ? valid_850 : _GEN_850; // @[ICache.scala 68:{44,44}]
  wire  _GEN_852 = 10'h353 == req_r_addr[14:5] ? valid_851 : _GEN_851; // @[ICache.scala 68:{44,44}]
  wire  _GEN_853 = 10'h354 == req_r_addr[14:5] ? valid_852 : _GEN_852; // @[ICache.scala 68:{44,44}]
  wire  _GEN_854 = 10'h355 == req_r_addr[14:5] ? valid_853 : _GEN_853; // @[ICache.scala 68:{44,44}]
  wire  _GEN_855 = 10'h356 == req_r_addr[14:5] ? valid_854 : _GEN_854; // @[ICache.scala 68:{44,44}]
  wire  _GEN_856 = 10'h357 == req_r_addr[14:5] ? valid_855 : _GEN_855; // @[ICache.scala 68:{44,44}]
  wire  _GEN_857 = 10'h358 == req_r_addr[14:5] ? valid_856 : _GEN_856; // @[ICache.scala 68:{44,44}]
  wire  _GEN_858 = 10'h359 == req_r_addr[14:5] ? valid_857 : _GEN_857; // @[ICache.scala 68:{44,44}]
  wire  _GEN_859 = 10'h35a == req_r_addr[14:5] ? valid_858 : _GEN_858; // @[ICache.scala 68:{44,44}]
  wire  _GEN_860 = 10'h35b == req_r_addr[14:5] ? valid_859 : _GEN_859; // @[ICache.scala 68:{44,44}]
  wire  _GEN_861 = 10'h35c == req_r_addr[14:5] ? valid_860 : _GEN_860; // @[ICache.scala 68:{44,44}]
  wire  _GEN_862 = 10'h35d == req_r_addr[14:5] ? valid_861 : _GEN_861; // @[ICache.scala 68:{44,44}]
  wire  _GEN_863 = 10'h35e == req_r_addr[14:5] ? valid_862 : _GEN_862; // @[ICache.scala 68:{44,44}]
  wire  _GEN_864 = 10'h35f == req_r_addr[14:5] ? valid_863 : _GEN_863; // @[ICache.scala 68:{44,44}]
  wire  _GEN_865 = 10'h360 == req_r_addr[14:5] ? valid_864 : _GEN_864; // @[ICache.scala 68:{44,44}]
  wire  _GEN_866 = 10'h361 == req_r_addr[14:5] ? valid_865 : _GEN_865; // @[ICache.scala 68:{44,44}]
  wire  _GEN_867 = 10'h362 == req_r_addr[14:5] ? valid_866 : _GEN_866; // @[ICache.scala 68:{44,44}]
  wire  _GEN_868 = 10'h363 == req_r_addr[14:5] ? valid_867 : _GEN_867; // @[ICache.scala 68:{44,44}]
  wire  _GEN_869 = 10'h364 == req_r_addr[14:5] ? valid_868 : _GEN_868; // @[ICache.scala 68:{44,44}]
  wire  _GEN_870 = 10'h365 == req_r_addr[14:5] ? valid_869 : _GEN_869; // @[ICache.scala 68:{44,44}]
  wire  _GEN_871 = 10'h366 == req_r_addr[14:5] ? valid_870 : _GEN_870; // @[ICache.scala 68:{44,44}]
  wire  _GEN_872 = 10'h367 == req_r_addr[14:5] ? valid_871 : _GEN_871; // @[ICache.scala 68:{44,44}]
  wire  _GEN_873 = 10'h368 == req_r_addr[14:5] ? valid_872 : _GEN_872; // @[ICache.scala 68:{44,44}]
  wire  _GEN_874 = 10'h369 == req_r_addr[14:5] ? valid_873 : _GEN_873; // @[ICache.scala 68:{44,44}]
  wire  _GEN_875 = 10'h36a == req_r_addr[14:5] ? valid_874 : _GEN_874; // @[ICache.scala 68:{44,44}]
  wire  _GEN_876 = 10'h36b == req_r_addr[14:5] ? valid_875 : _GEN_875; // @[ICache.scala 68:{44,44}]
  wire  _GEN_877 = 10'h36c == req_r_addr[14:5] ? valid_876 : _GEN_876; // @[ICache.scala 68:{44,44}]
  wire  _GEN_878 = 10'h36d == req_r_addr[14:5] ? valid_877 : _GEN_877; // @[ICache.scala 68:{44,44}]
  wire  _GEN_879 = 10'h36e == req_r_addr[14:5] ? valid_878 : _GEN_878; // @[ICache.scala 68:{44,44}]
  wire  _GEN_880 = 10'h36f == req_r_addr[14:5] ? valid_879 : _GEN_879; // @[ICache.scala 68:{44,44}]
  wire  _GEN_881 = 10'h370 == req_r_addr[14:5] ? valid_880 : _GEN_880; // @[ICache.scala 68:{44,44}]
  wire  _GEN_882 = 10'h371 == req_r_addr[14:5] ? valid_881 : _GEN_881; // @[ICache.scala 68:{44,44}]
  wire  _GEN_883 = 10'h372 == req_r_addr[14:5] ? valid_882 : _GEN_882; // @[ICache.scala 68:{44,44}]
  wire  _GEN_884 = 10'h373 == req_r_addr[14:5] ? valid_883 : _GEN_883; // @[ICache.scala 68:{44,44}]
  wire  _GEN_885 = 10'h374 == req_r_addr[14:5] ? valid_884 : _GEN_884; // @[ICache.scala 68:{44,44}]
  wire  _GEN_886 = 10'h375 == req_r_addr[14:5] ? valid_885 : _GEN_885; // @[ICache.scala 68:{44,44}]
  wire  _GEN_887 = 10'h376 == req_r_addr[14:5] ? valid_886 : _GEN_886; // @[ICache.scala 68:{44,44}]
  wire  _GEN_888 = 10'h377 == req_r_addr[14:5] ? valid_887 : _GEN_887; // @[ICache.scala 68:{44,44}]
  wire  _GEN_889 = 10'h378 == req_r_addr[14:5] ? valid_888 : _GEN_888; // @[ICache.scala 68:{44,44}]
  wire  _GEN_890 = 10'h379 == req_r_addr[14:5] ? valid_889 : _GEN_889; // @[ICache.scala 68:{44,44}]
  wire  _GEN_891 = 10'h37a == req_r_addr[14:5] ? valid_890 : _GEN_890; // @[ICache.scala 68:{44,44}]
  wire  _GEN_892 = 10'h37b == req_r_addr[14:5] ? valid_891 : _GEN_891; // @[ICache.scala 68:{44,44}]
  wire  _GEN_893 = 10'h37c == req_r_addr[14:5] ? valid_892 : _GEN_892; // @[ICache.scala 68:{44,44}]
  wire  _GEN_894 = 10'h37d == req_r_addr[14:5] ? valid_893 : _GEN_893; // @[ICache.scala 68:{44,44}]
  wire  _GEN_895 = 10'h37e == req_r_addr[14:5] ? valid_894 : _GEN_894; // @[ICache.scala 68:{44,44}]
  wire  _GEN_896 = 10'h37f == req_r_addr[14:5] ? valid_895 : _GEN_895; // @[ICache.scala 68:{44,44}]
  wire  _GEN_897 = 10'h380 == req_r_addr[14:5] ? valid_896 : _GEN_896; // @[ICache.scala 68:{44,44}]
  wire  _GEN_898 = 10'h381 == req_r_addr[14:5] ? valid_897 : _GEN_897; // @[ICache.scala 68:{44,44}]
  wire  _GEN_899 = 10'h382 == req_r_addr[14:5] ? valid_898 : _GEN_898; // @[ICache.scala 68:{44,44}]
  wire  _GEN_900 = 10'h383 == req_r_addr[14:5] ? valid_899 : _GEN_899; // @[ICache.scala 68:{44,44}]
  wire  _GEN_901 = 10'h384 == req_r_addr[14:5] ? valid_900 : _GEN_900; // @[ICache.scala 68:{44,44}]
  wire  _GEN_902 = 10'h385 == req_r_addr[14:5] ? valid_901 : _GEN_901; // @[ICache.scala 68:{44,44}]
  wire  _GEN_903 = 10'h386 == req_r_addr[14:5] ? valid_902 : _GEN_902; // @[ICache.scala 68:{44,44}]
  wire  _GEN_904 = 10'h387 == req_r_addr[14:5] ? valid_903 : _GEN_903; // @[ICache.scala 68:{44,44}]
  wire  _GEN_905 = 10'h388 == req_r_addr[14:5] ? valid_904 : _GEN_904; // @[ICache.scala 68:{44,44}]
  wire  _GEN_906 = 10'h389 == req_r_addr[14:5] ? valid_905 : _GEN_905; // @[ICache.scala 68:{44,44}]
  wire  _GEN_907 = 10'h38a == req_r_addr[14:5] ? valid_906 : _GEN_906; // @[ICache.scala 68:{44,44}]
  wire  _GEN_908 = 10'h38b == req_r_addr[14:5] ? valid_907 : _GEN_907; // @[ICache.scala 68:{44,44}]
  wire  _GEN_909 = 10'h38c == req_r_addr[14:5] ? valid_908 : _GEN_908; // @[ICache.scala 68:{44,44}]
  wire  _GEN_910 = 10'h38d == req_r_addr[14:5] ? valid_909 : _GEN_909; // @[ICache.scala 68:{44,44}]
  wire  _GEN_911 = 10'h38e == req_r_addr[14:5] ? valid_910 : _GEN_910; // @[ICache.scala 68:{44,44}]
  wire  _GEN_912 = 10'h38f == req_r_addr[14:5] ? valid_911 : _GEN_911; // @[ICache.scala 68:{44,44}]
  wire  _GEN_913 = 10'h390 == req_r_addr[14:5] ? valid_912 : _GEN_912; // @[ICache.scala 68:{44,44}]
  wire  _GEN_914 = 10'h391 == req_r_addr[14:5] ? valid_913 : _GEN_913; // @[ICache.scala 68:{44,44}]
  wire  _GEN_915 = 10'h392 == req_r_addr[14:5] ? valid_914 : _GEN_914; // @[ICache.scala 68:{44,44}]
  wire  _GEN_916 = 10'h393 == req_r_addr[14:5] ? valid_915 : _GEN_915; // @[ICache.scala 68:{44,44}]
  wire  _GEN_917 = 10'h394 == req_r_addr[14:5] ? valid_916 : _GEN_916; // @[ICache.scala 68:{44,44}]
  wire  _GEN_918 = 10'h395 == req_r_addr[14:5] ? valid_917 : _GEN_917; // @[ICache.scala 68:{44,44}]
  wire  _GEN_919 = 10'h396 == req_r_addr[14:5] ? valid_918 : _GEN_918; // @[ICache.scala 68:{44,44}]
  wire  _GEN_920 = 10'h397 == req_r_addr[14:5] ? valid_919 : _GEN_919; // @[ICache.scala 68:{44,44}]
  wire  _GEN_921 = 10'h398 == req_r_addr[14:5] ? valid_920 : _GEN_920; // @[ICache.scala 68:{44,44}]
  wire  _GEN_922 = 10'h399 == req_r_addr[14:5] ? valid_921 : _GEN_921; // @[ICache.scala 68:{44,44}]
  wire  _GEN_923 = 10'h39a == req_r_addr[14:5] ? valid_922 : _GEN_922; // @[ICache.scala 68:{44,44}]
  wire  _GEN_924 = 10'h39b == req_r_addr[14:5] ? valid_923 : _GEN_923; // @[ICache.scala 68:{44,44}]
  wire  _GEN_925 = 10'h39c == req_r_addr[14:5] ? valid_924 : _GEN_924; // @[ICache.scala 68:{44,44}]
  wire  _GEN_926 = 10'h39d == req_r_addr[14:5] ? valid_925 : _GEN_925; // @[ICache.scala 68:{44,44}]
  wire  _GEN_927 = 10'h39e == req_r_addr[14:5] ? valid_926 : _GEN_926; // @[ICache.scala 68:{44,44}]
  wire  _GEN_928 = 10'h39f == req_r_addr[14:5] ? valid_927 : _GEN_927; // @[ICache.scala 68:{44,44}]
  wire  _GEN_929 = 10'h3a0 == req_r_addr[14:5] ? valid_928 : _GEN_928; // @[ICache.scala 68:{44,44}]
  wire  _GEN_930 = 10'h3a1 == req_r_addr[14:5] ? valid_929 : _GEN_929; // @[ICache.scala 68:{44,44}]
  wire  _GEN_931 = 10'h3a2 == req_r_addr[14:5] ? valid_930 : _GEN_930; // @[ICache.scala 68:{44,44}]
  wire  _GEN_932 = 10'h3a3 == req_r_addr[14:5] ? valid_931 : _GEN_931; // @[ICache.scala 68:{44,44}]
  wire  _GEN_933 = 10'h3a4 == req_r_addr[14:5] ? valid_932 : _GEN_932; // @[ICache.scala 68:{44,44}]
  wire  _GEN_934 = 10'h3a5 == req_r_addr[14:5] ? valid_933 : _GEN_933; // @[ICache.scala 68:{44,44}]
  wire  _GEN_935 = 10'h3a6 == req_r_addr[14:5] ? valid_934 : _GEN_934; // @[ICache.scala 68:{44,44}]
  wire  _GEN_936 = 10'h3a7 == req_r_addr[14:5] ? valid_935 : _GEN_935; // @[ICache.scala 68:{44,44}]
  wire  _GEN_937 = 10'h3a8 == req_r_addr[14:5] ? valid_936 : _GEN_936; // @[ICache.scala 68:{44,44}]
  wire  _GEN_938 = 10'h3a9 == req_r_addr[14:5] ? valid_937 : _GEN_937; // @[ICache.scala 68:{44,44}]
  wire  _GEN_939 = 10'h3aa == req_r_addr[14:5] ? valid_938 : _GEN_938; // @[ICache.scala 68:{44,44}]
  wire  _GEN_940 = 10'h3ab == req_r_addr[14:5] ? valid_939 : _GEN_939; // @[ICache.scala 68:{44,44}]
  wire  _GEN_941 = 10'h3ac == req_r_addr[14:5] ? valid_940 : _GEN_940; // @[ICache.scala 68:{44,44}]
  wire  _GEN_942 = 10'h3ad == req_r_addr[14:5] ? valid_941 : _GEN_941; // @[ICache.scala 68:{44,44}]
  wire  _GEN_943 = 10'h3ae == req_r_addr[14:5] ? valid_942 : _GEN_942; // @[ICache.scala 68:{44,44}]
  wire  _GEN_944 = 10'h3af == req_r_addr[14:5] ? valid_943 : _GEN_943; // @[ICache.scala 68:{44,44}]
  wire  _GEN_945 = 10'h3b0 == req_r_addr[14:5] ? valid_944 : _GEN_944; // @[ICache.scala 68:{44,44}]
  wire  _GEN_946 = 10'h3b1 == req_r_addr[14:5] ? valid_945 : _GEN_945; // @[ICache.scala 68:{44,44}]
  wire  _GEN_947 = 10'h3b2 == req_r_addr[14:5] ? valid_946 : _GEN_946; // @[ICache.scala 68:{44,44}]
  wire  _GEN_948 = 10'h3b3 == req_r_addr[14:5] ? valid_947 : _GEN_947; // @[ICache.scala 68:{44,44}]
  wire  _GEN_949 = 10'h3b4 == req_r_addr[14:5] ? valid_948 : _GEN_948; // @[ICache.scala 68:{44,44}]
  wire  _GEN_950 = 10'h3b5 == req_r_addr[14:5] ? valid_949 : _GEN_949; // @[ICache.scala 68:{44,44}]
  wire  _GEN_951 = 10'h3b6 == req_r_addr[14:5] ? valid_950 : _GEN_950; // @[ICache.scala 68:{44,44}]
  wire  _GEN_952 = 10'h3b7 == req_r_addr[14:5] ? valid_951 : _GEN_951; // @[ICache.scala 68:{44,44}]
  wire  _GEN_953 = 10'h3b8 == req_r_addr[14:5] ? valid_952 : _GEN_952; // @[ICache.scala 68:{44,44}]
  wire  _GEN_954 = 10'h3b9 == req_r_addr[14:5] ? valid_953 : _GEN_953; // @[ICache.scala 68:{44,44}]
  wire  _GEN_955 = 10'h3ba == req_r_addr[14:5] ? valid_954 : _GEN_954; // @[ICache.scala 68:{44,44}]
  wire  _GEN_956 = 10'h3bb == req_r_addr[14:5] ? valid_955 : _GEN_955; // @[ICache.scala 68:{44,44}]
  wire  _GEN_957 = 10'h3bc == req_r_addr[14:5] ? valid_956 : _GEN_956; // @[ICache.scala 68:{44,44}]
  wire  _GEN_958 = 10'h3bd == req_r_addr[14:5] ? valid_957 : _GEN_957; // @[ICache.scala 68:{44,44}]
  wire  _GEN_959 = 10'h3be == req_r_addr[14:5] ? valid_958 : _GEN_958; // @[ICache.scala 68:{44,44}]
  wire  _GEN_960 = 10'h3bf == req_r_addr[14:5] ? valid_959 : _GEN_959; // @[ICache.scala 68:{44,44}]
  wire  _GEN_961 = 10'h3c0 == req_r_addr[14:5] ? valid_960 : _GEN_960; // @[ICache.scala 68:{44,44}]
  wire  _GEN_962 = 10'h3c1 == req_r_addr[14:5] ? valid_961 : _GEN_961; // @[ICache.scala 68:{44,44}]
  wire  _GEN_963 = 10'h3c2 == req_r_addr[14:5] ? valid_962 : _GEN_962; // @[ICache.scala 68:{44,44}]
  wire  _GEN_964 = 10'h3c3 == req_r_addr[14:5] ? valid_963 : _GEN_963; // @[ICache.scala 68:{44,44}]
  wire  _GEN_965 = 10'h3c4 == req_r_addr[14:5] ? valid_964 : _GEN_964; // @[ICache.scala 68:{44,44}]
  wire  _GEN_966 = 10'h3c5 == req_r_addr[14:5] ? valid_965 : _GEN_965; // @[ICache.scala 68:{44,44}]
  wire  _GEN_967 = 10'h3c6 == req_r_addr[14:5] ? valid_966 : _GEN_966; // @[ICache.scala 68:{44,44}]
  wire  _GEN_968 = 10'h3c7 == req_r_addr[14:5] ? valid_967 : _GEN_967; // @[ICache.scala 68:{44,44}]
  wire  _GEN_969 = 10'h3c8 == req_r_addr[14:5] ? valid_968 : _GEN_968; // @[ICache.scala 68:{44,44}]
  wire  _GEN_970 = 10'h3c9 == req_r_addr[14:5] ? valid_969 : _GEN_969; // @[ICache.scala 68:{44,44}]
  wire  _GEN_971 = 10'h3ca == req_r_addr[14:5] ? valid_970 : _GEN_970; // @[ICache.scala 68:{44,44}]
  wire  _GEN_972 = 10'h3cb == req_r_addr[14:5] ? valid_971 : _GEN_971; // @[ICache.scala 68:{44,44}]
  wire  _GEN_973 = 10'h3cc == req_r_addr[14:5] ? valid_972 : _GEN_972; // @[ICache.scala 68:{44,44}]
  wire  _GEN_974 = 10'h3cd == req_r_addr[14:5] ? valid_973 : _GEN_973; // @[ICache.scala 68:{44,44}]
  wire  _GEN_975 = 10'h3ce == req_r_addr[14:5] ? valid_974 : _GEN_974; // @[ICache.scala 68:{44,44}]
  wire  _GEN_976 = 10'h3cf == req_r_addr[14:5] ? valid_975 : _GEN_975; // @[ICache.scala 68:{44,44}]
  wire  _GEN_977 = 10'h3d0 == req_r_addr[14:5] ? valid_976 : _GEN_976; // @[ICache.scala 68:{44,44}]
  wire  _GEN_978 = 10'h3d1 == req_r_addr[14:5] ? valid_977 : _GEN_977; // @[ICache.scala 68:{44,44}]
  wire  _GEN_979 = 10'h3d2 == req_r_addr[14:5] ? valid_978 : _GEN_978; // @[ICache.scala 68:{44,44}]
  wire  _GEN_980 = 10'h3d3 == req_r_addr[14:5] ? valid_979 : _GEN_979; // @[ICache.scala 68:{44,44}]
  wire  _GEN_981 = 10'h3d4 == req_r_addr[14:5] ? valid_980 : _GEN_980; // @[ICache.scala 68:{44,44}]
  wire  _GEN_982 = 10'h3d5 == req_r_addr[14:5] ? valid_981 : _GEN_981; // @[ICache.scala 68:{44,44}]
  wire  _GEN_983 = 10'h3d6 == req_r_addr[14:5] ? valid_982 : _GEN_982; // @[ICache.scala 68:{44,44}]
  wire  _GEN_984 = 10'h3d7 == req_r_addr[14:5] ? valid_983 : _GEN_983; // @[ICache.scala 68:{44,44}]
  wire  _GEN_985 = 10'h3d8 == req_r_addr[14:5] ? valid_984 : _GEN_984; // @[ICache.scala 68:{44,44}]
  wire  _GEN_986 = 10'h3d9 == req_r_addr[14:5] ? valid_985 : _GEN_985; // @[ICache.scala 68:{44,44}]
  wire  _GEN_987 = 10'h3da == req_r_addr[14:5] ? valid_986 : _GEN_986; // @[ICache.scala 68:{44,44}]
  wire  _GEN_988 = 10'h3db == req_r_addr[14:5] ? valid_987 : _GEN_987; // @[ICache.scala 68:{44,44}]
  wire  _GEN_989 = 10'h3dc == req_r_addr[14:5] ? valid_988 : _GEN_988; // @[ICache.scala 68:{44,44}]
  wire  _GEN_990 = 10'h3dd == req_r_addr[14:5] ? valid_989 : _GEN_989; // @[ICache.scala 68:{44,44}]
  wire  _GEN_991 = 10'h3de == req_r_addr[14:5] ? valid_990 : _GEN_990; // @[ICache.scala 68:{44,44}]
  wire  _GEN_992 = 10'h3df == req_r_addr[14:5] ? valid_991 : _GEN_991; // @[ICache.scala 68:{44,44}]
  wire  _GEN_993 = 10'h3e0 == req_r_addr[14:5] ? valid_992 : _GEN_992; // @[ICache.scala 68:{44,44}]
  wire  _GEN_994 = 10'h3e1 == req_r_addr[14:5] ? valid_993 : _GEN_993; // @[ICache.scala 68:{44,44}]
  wire  _GEN_995 = 10'h3e2 == req_r_addr[14:5] ? valid_994 : _GEN_994; // @[ICache.scala 68:{44,44}]
  wire  _GEN_996 = 10'h3e3 == req_r_addr[14:5] ? valid_995 : _GEN_995; // @[ICache.scala 68:{44,44}]
  wire  _GEN_997 = 10'h3e4 == req_r_addr[14:5] ? valid_996 : _GEN_996; // @[ICache.scala 68:{44,44}]
  wire  _GEN_998 = 10'h3e5 == req_r_addr[14:5] ? valid_997 : _GEN_997; // @[ICache.scala 68:{44,44}]
  wire  _GEN_999 = 10'h3e6 == req_r_addr[14:5] ? valid_998 : _GEN_998; // @[ICache.scala 68:{44,44}]
  wire  _GEN_1000 = 10'h3e7 == req_r_addr[14:5] ? valid_999 : _GEN_999; // @[ICache.scala 68:{44,44}]
  wire  _GEN_1001 = 10'h3e8 == req_r_addr[14:5] ? valid_1000 : _GEN_1000; // @[ICache.scala 68:{44,44}]
  wire  _GEN_1002 = 10'h3e9 == req_r_addr[14:5] ? valid_1001 : _GEN_1001; // @[ICache.scala 68:{44,44}]
  wire  _GEN_1003 = 10'h3ea == req_r_addr[14:5] ? valid_1002 : _GEN_1002; // @[ICache.scala 68:{44,44}]
  wire  _GEN_1004 = 10'h3eb == req_r_addr[14:5] ? valid_1003 : _GEN_1003; // @[ICache.scala 68:{44,44}]
  wire  _GEN_1005 = 10'h3ec == req_r_addr[14:5] ? valid_1004 : _GEN_1004; // @[ICache.scala 68:{44,44}]
  wire  _GEN_1006 = 10'h3ed == req_r_addr[14:5] ? valid_1005 : _GEN_1005; // @[ICache.scala 68:{44,44}]
  wire  _GEN_1007 = 10'h3ee == req_r_addr[14:5] ? valid_1006 : _GEN_1006; // @[ICache.scala 68:{44,44}]
  wire  _GEN_1008 = 10'h3ef == req_r_addr[14:5] ? valid_1007 : _GEN_1007; // @[ICache.scala 68:{44,44}]
  wire  _GEN_1009 = 10'h3f0 == req_r_addr[14:5] ? valid_1008 : _GEN_1008; // @[ICache.scala 68:{44,44}]
  wire  _GEN_1010 = 10'h3f1 == req_r_addr[14:5] ? valid_1009 : _GEN_1009; // @[ICache.scala 68:{44,44}]
  wire  _GEN_1011 = 10'h3f2 == req_r_addr[14:5] ? valid_1010 : _GEN_1010; // @[ICache.scala 68:{44,44}]
  wire  _GEN_1012 = 10'h3f3 == req_r_addr[14:5] ? valid_1011 : _GEN_1011; // @[ICache.scala 68:{44,44}]
  wire  _GEN_1013 = 10'h3f4 == req_r_addr[14:5] ? valid_1012 : _GEN_1012; // @[ICache.scala 68:{44,44}]
  wire  _GEN_1014 = 10'h3f5 == req_r_addr[14:5] ? valid_1013 : _GEN_1013; // @[ICache.scala 68:{44,44}]
  wire  _GEN_1015 = 10'h3f6 == req_r_addr[14:5] ? valid_1014 : _GEN_1014; // @[ICache.scala 68:{44,44}]
  wire  _GEN_1016 = 10'h3f7 == req_r_addr[14:5] ? valid_1015 : _GEN_1015; // @[ICache.scala 68:{44,44}]
  wire  _GEN_1017 = 10'h3f8 == req_r_addr[14:5] ? valid_1016 : _GEN_1016; // @[ICache.scala 68:{44,44}]
  wire  _GEN_1018 = 10'h3f9 == req_r_addr[14:5] ? valid_1017 : _GEN_1017; // @[ICache.scala 68:{44,44}]
  wire  _GEN_1019 = 10'h3fa == req_r_addr[14:5] ? valid_1018 : _GEN_1018; // @[ICache.scala 68:{44,44}]
  wire  _GEN_1020 = 10'h3fb == req_r_addr[14:5] ? valid_1019 : _GEN_1019; // @[ICache.scala 68:{44,44}]
  wire  _GEN_1021 = 10'h3fc == req_r_addr[14:5] ? valid_1020 : _GEN_1020; // @[ICache.scala 68:{44,44}]
  wire  _GEN_1022 = 10'h3fd == req_r_addr[14:5] ? valid_1021 : _GEN_1021; // @[ICache.scala 68:{44,44}]
  wire  _GEN_1023 = 10'h3fe == req_r_addr[14:5] ? valid_1022 : _GEN_1022; // @[ICache.scala 68:{44,44}]
  wire  _GEN_1024 = 10'h3ff == req_r_addr[14:5] ? valid_1023 : _GEN_1023; // @[ICache.scala 68:{44,44}]
  reg  array_out_REG; // @[ICache.scala 67:50]
  reg [272:0] array_out_r; // @[Reg.scala 35:20]
  wire [272:0] _array_out_T = array_out_REG ? array_io_rdata : array_out_r; // @[Utils.scala 50:8]
  wire [16:0] array_out_tag = _array_out_T[272:256]; // @[ICache.scala 67:66]
  wire  array_hit = _GEN_1024 & req_r_addr[31:15] == array_out_tag; // @[ICache.scala 68:44]
  wire  _s2_ready_T_1 = state == 3'h0 & array_hit; // @[ICache.scala 143:35]
  wire  _s2_ready_T_2 = state == 3'h3; // @[ICache.scala 143:59]
  wire  s2_ready = (state == 3'h0 & array_hit | state == 3'h3 | state == 3'h4) & io_cache_resp_ready; // @[ICache.scala 143:92]
  wire  fire = io_cache_req_valid & s2_ready; // @[ICache.scala 56:27]
  wire  tl_d_ready = state == 3'h2; // @[ICache.scala 152:24]
  wire  _array_io_en_T = tl_d_ready & auto_out_d_valid; // @[Decoupled.scala 51:35]
  wire [255:0] array_out_data = _array_out_T[255:0]; // @[ICache.scala 67:66]
  wire [9:0] _GEN_1025 = fire ? io_cache_req_bits_addr[14:5] : 10'h0; // @[ICache.scala 71:14 60:18 72:19]
  wire  _state_T = io_cache_resp_ready & io_cache_resp_valid; // @[Decoupled.scala 51:35]
  wire  _state_T_1 = io_cache_req_ready & io_cache_req_valid; // @[Decoupled.scala 51:35]
  wire  _state_T_2 = ~_state_T_1; // @[ICache.scala 82:33]
  wire  tl_a_valid = state == 3'h1; // @[ICache.scala 150:24]
  wire  _T_2 = auto_out_a_ready & tl_a_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_1034 = _array_io_en_T ? 3'h3 : state; // @[ICache.scala 90:23 91:15 78:68]
  wire [2:0] _state_T_8 = _state_T_2 ? 3'h4 : 3'h0; // @[ICache.scala 96:21]
  wire [2:0] _GEN_1035 = _state_T ? _state_T_8 : state; // @[ICache.scala 95:23 96:15 78:68]
  wire [2:0] _GEN_1036 = _state_T_1 ? 3'h0 : state; // @[ICache.scala 100:22 101:15 78:68]
  wire [2:0] _GEN_1037 = 3'h4 == state ? _GEN_1036 : state; // @[ICache.scala 80:17 78:68]
  wire [2:0] _GEN_1038 = 3'h3 == state ? _GEN_1035 : _GEN_1037; // @[ICache.scala 80:17]
  wire [63:0] _array_data_T_6 = 2'h1 == req_r_addr[4:3] ? array_out_data[127:64] : array_out_data[63:0]; // @[Mux.scala 81:58]
  wire [63:0] _array_data_T_8 = 2'h2 == req_r_addr[4:3] ? array_out_data[191:128] : _array_data_T_6; // @[Mux.scala 81:58]
  wire [63:0] _array_data_T_10 = 2'h3 == req_r_addr[4:3] ? array_out_data[255:192] : _array_data_T_8; // @[Mux.scala 81:58]
  reg  array_data_REG; // @[ICache.scala 118:12]
  reg [63:0] array_data_r; // @[Reg.scala 35:20]
  wire [63:0] _GEN_1042 = array_data_REG ? _array_data_T_10 : array_data_r; // @[Reg.scala 36:18 35:20 36:22]
  reg [255:0] wdata; // @[Reg.scala 35:20]
  wire [272:0] _array_io_wdata_T_1 = {req_r_addr[31:15],auto_out_d_bits_data}; // @[Cat.scala 33:92]
  wire  _GEN_1044 = 10'h0 == req_r_addr[14:5] | valid_0; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1045 = 10'h1 == req_r_addr[14:5] | valid_1; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1046 = 10'h2 == req_r_addr[14:5] | valid_2; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1047 = 10'h3 == req_r_addr[14:5] | valid_3; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1048 = 10'h4 == req_r_addr[14:5] | valid_4; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1049 = 10'h5 == req_r_addr[14:5] | valid_5; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1050 = 10'h6 == req_r_addr[14:5] | valid_6; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1051 = 10'h7 == req_r_addr[14:5] | valid_7; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1052 = 10'h8 == req_r_addr[14:5] | valid_8; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1053 = 10'h9 == req_r_addr[14:5] | valid_9; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1054 = 10'ha == req_r_addr[14:5] | valid_10; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1055 = 10'hb == req_r_addr[14:5] | valid_11; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1056 = 10'hc == req_r_addr[14:5] | valid_12; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1057 = 10'hd == req_r_addr[14:5] | valid_13; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1058 = 10'he == req_r_addr[14:5] | valid_14; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1059 = 10'hf == req_r_addr[14:5] | valid_15; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1060 = 10'h10 == req_r_addr[14:5] | valid_16; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1061 = 10'h11 == req_r_addr[14:5] | valid_17; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1062 = 10'h12 == req_r_addr[14:5] | valid_18; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1063 = 10'h13 == req_r_addr[14:5] | valid_19; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1064 = 10'h14 == req_r_addr[14:5] | valid_20; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1065 = 10'h15 == req_r_addr[14:5] | valid_21; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1066 = 10'h16 == req_r_addr[14:5] | valid_22; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1067 = 10'h17 == req_r_addr[14:5] | valid_23; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1068 = 10'h18 == req_r_addr[14:5] | valid_24; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1069 = 10'h19 == req_r_addr[14:5] | valid_25; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1070 = 10'h1a == req_r_addr[14:5] | valid_26; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1071 = 10'h1b == req_r_addr[14:5] | valid_27; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1072 = 10'h1c == req_r_addr[14:5] | valid_28; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1073 = 10'h1d == req_r_addr[14:5] | valid_29; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1074 = 10'h1e == req_r_addr[14:5] | valid_30; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1075 = 10'h1f == req_r_addr[14:5] | valid_31; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1076 = 10'h20 == req_r_addr[14:5] | valid_32; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1077 = 10'h21 == req_r_addr[14:5] | valid_33; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1078 = 10'h22 == req_r_addr[14:5] | valid_34; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1079 = 10'h23 == req_r_addr[14:5] | valid_35; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1080 = 10'h24 == req_r_addr[14:5] | valid_36; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1081 = 10'h25 == req_r_addr[14:5] | valid_37; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1082 = 10'h26 == req_r_addr[14:5] | valid_38; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1083 = 10'h27 == req_r_addr[14:5] | valid_39; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1084 = 10'h28 == req_r_addr[14:5] | valid_40; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1085 = 10'h29 == req_r_addr[14:5] | valid_41; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1086 = 10'h2a == req_r_addr[14:5] | valid_42; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1087 = 10'h2b == req_r_addr[14:5] | valid_43; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1088 = 10'h2c == req_r_addr[14:5] | valid_44; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1089 = 10'h2d == req_r_addr[14:5] | valid_45; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1090 = 10'h2e == req_r_addr[14:5] | valid_46; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1091 = 10'h2f == req_r_addr[14:5] | valid_47; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1092 = 10'h30 == req_r_addr[14:5] | valid_48; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1093 = 10'h31 == req_r_addr[14:5] | valid_49; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1094 = 10'h32 == req_r_addr[14:5] | valid_50; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1095 = 10'h33 == req_r_addr[14:5] | valid_51; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1096 = 10'h34 == req_r_addr[14:5] | valid_52; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1097 = 10'h35 == req_r_addr[14:5] | valid_53; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1098 = 10'h36 == req_r_addr[14:5] | valid_54; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1099 = 10'h37 == req_r_addr[14:5] | valid_55; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1100 = 10'h38 == req_r_addr[14:5] | valid_56; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1101 = 10'h39 == req_r_addr[14:5] | valid_57; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1102 = 10'h3a == req_r_addr[14:5] | valid_58; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1103 = 10'h3b == req_r_addr[14:5] | valid_59; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1104 = 10'h3c == req_r_addr[14:5] | valid_60; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1105 = 10'h3d == req_r_addr[14:5] | valid_61; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1106 = 10'h3e == req_r_addr[14:5] | valid_62; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1107 = 10'h3f == req_r_addr[14:5] | valid_63; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1108 = 10'h40 == req_r_addr[14:5] | valid_64; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1109 = 10'h41 == req_r_addr[14:5] | valid_65; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1110 = 10'h42 == req_r_addr[14:5] | valid_66; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1111 = 10'h43 == req_r_addr[14:5] | valid_67; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1112 = 10'h44 == req_r_addr[14:5] | valid_68; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1113 = 10'h45 == req_r_addr[14:5] | valid_69; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1114 = 10'h46 == req_r_addr[14:5] | valid_70; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1115 = 10'h47 == req_r_addr[14:5] | valid_71; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1116 = 10'h48 == req_r_addr[14:5] | valid_72; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1117 = 10'h49 == req_r_addr[14:5] | valid_73; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1118 = 10'h4a == req_r_addr[14:5] | valid_74; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1119 = 10'h4b == req_r_addr[14:5] | valid_75; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1120 = 10'h4c == req_r_addr[14:5] | valid_76; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1121 = 10'h4d == req_r_addr[14:5] | valid_77; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1122 = 10'h4e == req_r_addr[14:5] | valid_78; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1123 = 10'h4f == req_r_addr[14:5] | valid_79; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1124 = 10'h50 == req_r_addr[14:5] | valid_80; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1125 = 10'h51 == req_r_addr[14:5] | valid_81; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1126 = 10'h52 == req_r_addr[14:5] | valid_82; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1127 = 10'h53 == req_r_addr[14:5] | valid_83; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1128 = 10'h54 == req_r_addr[14:5] | valid_84; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1129 = 10'h55 == req_r_addr[14:5] | valid_85; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1130 = 10'h56 == req_r_addr[14:5] | valid_86; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1131 = 10'h57 == req_r_addr[14:5] | valid_87; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1132 = 10'h58 == req_r_addr[14:5] | valid_88; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1133 = 10'h59 == req_r_addr[14:5] | valid_89; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1134 = 10'h5a == req_r_addr[14:5] | valid_90; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1135 = 10'h5b == req_r_addr[14:5] | valid_91; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1136 = 10'h5c == req_r_addr[14:5] | valid_92; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1137 = 10'h5d == req_r_addr[14:5] | valid_93; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1138 = 10'h5e == req_r_addr[14:5] | valid_94; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1139 = 10'h5f == req_r_addr[14:5] | valid_95; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1140 = 10'h60 == req_r_addr[14:5] | valid_96; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1141 = 10'h61 == req_r_addr[14:5] | valid_97; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1142 = 10'h62 == req_r_addr[14:5] | valid_98; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1143 = 10'h63 == req_r_addr[14:5] | valid_99; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1144 = 10'h64 == req_r_addr[14:5] | valid_100; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1145 = 10'h65 == req_r_addr[14:5] | valid_101; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1146 = 10'h66 == req_r_addr[14:5] | valid_102; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1147 = 10'h67 == req_r_addr[14:5] | valid_103; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1148 = 10'h68 == req_r_addr[14:5] | valid_104; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1149 = 10'h69 == req_r_addr[14:5] | valid_105; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1150 = 10'h6a == req_r_addr[14:5] | valid_106; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1151 = 10'h6b == req_r_addr[14:5] | valid_107; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1152 = 10'h6c == req_r_addr[14:5] | valid_108; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1153 = 10'h6d == req_r_addr[14:5] | valid_109; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1154 = 10'h6e == req_r_addr[14:5] | valid_110; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1155 = 10'h6f == req_r_addr[14:5] | valid_111; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1156 = 10'h70 == req_r_addr[14:5] | valid_112; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1157 = 10'h71 == req_r_addr[14:5] | valid_113; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1158 = 10'h72 == req_r_addr[14:5] | valid_114; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1159 = 10'h73 == req_r_addr[14:5] | valid_115; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1160 = 10'h74 == req_r_addr[14:5] | valid_116; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1161 = 10'h75 == req_r_addr[14:5] | valid_117; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1162 = 10'h76 == req_r_addr[14:5] | valid_118; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1163 = 10'h77 == req_r_addr[14:5] | valid_119; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1164 = 10'h78 == req_r_addr[14:5] | valid_120; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1165 = 10'h79 == req_r_addr[14:5] | valid_121; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1166 = 10'h7a == req_r_addr[14:5] | valid_122; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1167 = 10'h7b == req_r_addr[14:5] | valid_123; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1168 = 10'h7c == req_r_addr[14:5] | valid_124; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1169 = 10'h7d == req_r_addr[14:5] | valid_125; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1170 = 10'h7e == req_r_addr[14:5] | valid_126; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1171 = 10'h7f == req_r_addr[14:5] | valid_127; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1172 = 10'h80 == req_r_addr[14:5] | valid_128; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1173 = 10'h81 == req_r_addr[14:5] | valid_129; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1174 = 10'h82 == req_r_addr[14:5] | valid_130; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1175 = 10'h83 == req_r_addr[14:5] | valid_131; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1176 = 10'h84 == req_r_addr[14:5] | valid_132; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1177 = 10'h85 == req_r_addr[14:5] | valid_133; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1178 = 10'h86 == req_r_addr[14:5] | valid_134; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1179 = 10'h87 == req_r_addr[14:5] | valid_135; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1180 = 10'h88 == req_r_addr[14:5] | valid_136; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1181 = 10'h89 == req_r_addr[14:5] | valid_137; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1182 = 10'h8a == req_r_addr[14:5] | valid_138; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1183 = 10'h8b == req_r_addr[14:5] | valid_139; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1184 = 10'h8c == req_r_addr[14:5] | valid_140; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1185 = 10'h8d == req_r_addr[14:5] | valid_141; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1186 = 10'h8e == req_r_addr[14:5] | valid_142; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1187 = 10'h8f == req_r_addr[14:5] | valid_143; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1188 = 10'h90 == req_r_addr[14:5] | valid_144; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1189 = 10'h91 == req_r_addr[14:5] | valid_145; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1190 = 10'h92 == req_r_addr[14:5] | valid_146; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1191 = 10'h93 == req_r_addr[14:5] | valid_147; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1192 = 10'h94 == req_r_addr[14:5] | valid_148; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1193 = 10'h95 == req_r_addr[14:5] | valid_149; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1194 = 10'h96 == req_r_addr[14:5] | valid_150; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1195 = 10'h97 == req_r_addr[14:5] | valid_151; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1196 = 10'h98 == req_r_addr[14:5] | valid_152; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1197 = 10'h99 == req_r_addr[14:5] | valid_153; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1198 = 10'h9a == req_r_addr[14:5] | valid_154; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1199 = 10'h9b == req_r_addr[14:5] | valid_155; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1200 = 10'h9c == req_r_addr[14:5] | valid_156; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1201 = 10'h9d == req_r_addr[14:5] | valid_157; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1202 = 10'h9e == req_r_addr[14:5] | valid_158; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1203 = 10'h9f == req_r_addr[14:5] | valid_159; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1204 = 10'ha0 == req_r_addr[14:5] | valid_160; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1205 = 10'ha1 == req_r_addr[14:5] | valid_161; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1206 = 10'ha2 == req_r_addr[14:5] | valid_162; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1207 = 10'ha3 == req_r_addr[14:5] | valid_163; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1208 = 10'ha4 == req_r_addr[14:5] | valid_164; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1209 = 10'ha5 == req_r_addr[14:5] | valid_165; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1210 = 10'ha6 == req_r_addr[14:5] | valid_166; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1211 = 10'ha7 == req_r_addr[14:5] | valid_167; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1212 = 10'ha8 == req_r_addr[14:5] | valid_168; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1213 = 10'ha9 == req_r_addr[14:5] | valid_169; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1214 = 10'haa == req_r_addr[14:5] | valid_170; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1215 = 10'hab == req_r_addr[14:5] | valid_171; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1216 = 10'hac == req_r_addr[14:5] | valid_172; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1217 = 10'had == req_r_addr[14:5] | valid_173; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1218 = 10'hae == req_r_addr[14:5] | valid_174; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1219 = 10'haf == req_r_addr[14:5] | valid_175; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1220 = 10'hb0 == req_r_addr[14:5] | valid_176; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1221 = 10'hb1 == req_r_addr[14:5] | valid_177; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1222 = 10'hb2 == req_r_addr[14:5] | valid_178; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1223 = 10'hb3 == req_r_addr[14:5] | valid_179; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1224 = 10'hb4 == req_r_addr[14:5] | valid_180; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1225 = 10'hb5 == req_r_addr[14:5] | valid_181; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1226 = 10'hb6 == req_r_addr[14:5] | valid_182; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1227 = 10'hb7 == req_r_addr[14:5] | valid_183; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1228 = 10'hb8 == req_r_addr[14:5] | valid_184; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1229 = 10'hb9 == req_r_addr[14:5] | valid_185; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1230 = 10'hba == req_r_addr[14:5] | valid_186; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1231 = 10'hbb == req_r_addr[14:5] | valid_187; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1232 = 10'hbc == req_r_addr[14:5] | valid_188; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1233 = 10'hbd == req_r_addr[14:5] | valid_189; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1234 = 10'hbe == req_r_addr[14:5] | valid_190; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1235 = 10'hbf == req_r_addr[14:5] | valid_191; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1236 = 10'hc0 == req_r_addr[14:5] | valid_192; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1237 = 10'hc1 == req_r_addr[14:5] | valid_193; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1238 = 10'hc2 == req_r_addr[14:5] | valid_194; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1239 = 10'hc3 == req_r_addr[14:5] | valid_195; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1240 = 10'hc4 == req_r_addr[14:5] | valid_196; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1241 = 10'hc5 == req_r_addr[14:5] | valid_197; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1242 = 10'hc6 == req_r_addr[14:5] | valid_198; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1243 = 10'hc7 == req_r_addr[14:5] | valid_199; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1244 = 10'hc8 == req_r_addr[14:5] | valid_200; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1245 = 10'hc9 == req_r_addr[14:5] | valid_201; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1246 = 10'hca == req_r_addr[14:5] | valid_202; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1247 = 10'hcb == req_r_addr[14:5] | valid_203; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1248 = 10'hcc == req_r_addr[14:5] | valid_204; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1249 = 10'hcd == req_r_addr[14:5] | valid_205; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1250 = 10'hce == req_r_addr[14:5] | valid_206; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1251 = 10'hcf == req_r_addr[14:5] | valid_207; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1252 = 10'hd0 == req_r_addr[14:5] | valid_208; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1253 = 10'hd1 == req_r_addr[14:5] | valid_209; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1254 = 10'hd2 == req_r_addr[14:5] | valid_210; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1255 = 10'hd3 == req_r_addr[14:5] | valid_211; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1256 = 10'hd4 == req_r_addr[14:5] | valid_212; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1257 = 10'hd5 == req_r_addr[14:5] | valid_213; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1258 = 10'hd6 == req_r_addr[14:5] | valid_214; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1259 = 10'hd7 == req_r_addr[14:5] | valid_215; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1260 = 10'hd8 == req_r_addr[14:5] | valid_216; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1261 = 10'hd9 == req_r_addr[14:5] | valid_217; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1262 = 10'hda == req_r_addr[14:5] | valid_218; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1263 = 10'hdb == req_r_addr[14:5] | valid_219; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1264 = 10'hdc == req_r_addr[14:5] | valid_220; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1265 = 10'hdd == req_r_addr[14:5] | valid_221; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1266 = 10'hde == req_r_addr[14:5] | valid_222; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1267 = 10'hdf == req_r_addr[14:5] | valid_223; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1268 = 10'he0 == req_r_addr[14:5] | valid_224; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1269 = 10'he1 == req_r_addr[14:5] | valid_225; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1270 = 10'he2 == req_r_addr[14:5] | valid_226; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1271 = 10'he3 == req_r_addr[14:5] | valid_227; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1272 = 10'he4 == req_r_addr[14:5] | valid_228; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1273 = 10'he5 == req_r_addr[14:5] | valid_229; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1274 = 10'he6 == req_r_addr[14:5] | valid_230; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1275 = 10'he7 == req_r_addr[14:5] | valid_231; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1276 = 10'he8 == req_r_addr[14:5] | valid_232; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1277 = 10'he9 == req_r_addr[14:5] | valid_233; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1278 = 10'hea == req_r_addr[14:5] | valid_234; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1279 = 10'heb == req_r_addr[14:5] | valid_235; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1280 = 10'hec == req_r_addr[14:5] | valid_236; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1281 = 10'hed == req_r_addr[14:5] | valid_237; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1282 = 10'hee == req_r_addr[14:5] | valid_238; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1283 = 10'hef == req_r_addr[14:5] | valid_239; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1284 = 10'hf0 == req_r_addr[14:5] | valid_240; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1285 = 10'hf1 == req_r_addr[14:5] | valid_241; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1286 = 10'hf2 == req_r_addr[14:5] | valid_242; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1287 = 10'hf3 == req_r_addr[14:5] | valid_243; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1288 = 10'hf4 == req_r_addr[14:5] | valid_244; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1289 = 10'hf5 == req_r_addr[14:5] | valid_245; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1290 = 10'hf6 == req_r_addr[14:5] | valid_246; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1291 = 10'hf7 == req_r_addr[14:5] | valid_247; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1292 = 10'hf8 == req_r_addr[14:5] | valid_248; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1293 = 10'hf9 == req_r_addr[14:5] | valid_249; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1294 = 10'hfa == req_r_addr[14:5] | valid_250; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1295 = 10'hfb == req_r_addr[14:5] | valid_251; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1296 = 10'hfc == req_r_addr[14:5] | valid_252; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1297 = 10'hfd == req_r_addr[14:5] | valid_253; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1298 = 10'hfe == req_r_addr[14:5] | valid_254; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1299 = 10'hff == req_r_addr[14:5] | valid_255; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1300 = 10'h100 == req_r_addr[14:5] | valid_256; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1301 = 10'h101 == req_r_addr[14:5] | valid_257; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1302 = 10'h102 == req_r_addr[14:5] | valid_258; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1303 = 10'h103 == req_r_addr[14:5] | valid_259; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1304 = 10'h104 == req_r_addr[14:5] | valid_260; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1305 = 10'h105 == req_r_addr[14:5] | valid_261; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1306 = 10'h106 == req_r_addr[14:5] | valid_262; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1307 = 10'h107 == req_r_addr[14:5] | valid_263; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1308 = 10'h108 == req_r_addr[14:5] | valid_264; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1309 = 10'h109 == req_r_addr[14:5] | valid_265; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1310 = 10'h10a == req_r_addr[14:5] | valid_266; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1311 = 10'h10b == req_r_addr[14:5] | valid_267; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1312 = 10'h10c == req_r_addr[14:5] | valid_268; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1313 = 10'h10d == req_r_addr[14:5] | valid_269; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1314 = 10'h10e == req_r_addr[14:5] | valid_270; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1315 = 10'h10f == req_r_addr[14:5] | valid_271; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1316 = 10'h110 == req_r_addr[14:5] | valid_272; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1317 = 10'h111 == req_r_addr[14:5] | valid_273; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1318 = 10'h112 == req_r_addr[14:5] | valid_274; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1319 = 10'h113 == req_r_addr[14:5] | valid_275; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1320 = 10'h114 == req_r_addr[14:5] | valid_276; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1321 = 10'h115 == req_r_addr[14:5] | valid_277; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1322 = 10'h116 == req_r_addr[14:5] | valid_278; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1323 = 10'h117 == req_r_addr[14:5] | valid_279; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1324 = 10'h118 == req_r_addr[14:5] | valid_280; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1325 = 10'h119 == req_r_addr[14:5] | valid_281; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1326 = 10'h11a == req_r_addr[14:5] | valid_282; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1327 = 10'h11b == req_r_addr[14:5] | valid_283; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1328 = 10'h11c == req_r_addr[14:5] | valid_284; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1329 = 10'h11d == req_r_addr[14:5] | valid_285; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1330 = 10'h11e == req_r_addr[14:5] | valid_286; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1331 = 10'h11f == req_r_addr[14:5] | valid_287; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1332 = 10'h120 == req_r_addr[14:5] | valid_288; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1333 = 10'h121 == req_r_addr[14:5] | valid_289; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1334 = 10'h122 == req_r_addr[14:5] | valid_290; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1335 = 10'h123 == req_r_addr[14:5] | valid_291; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1336 = 10'h124 == req_r_addr[14:5] | valid_292; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1337 = 10'h125 == req_r_addr[14:5] | valid_293; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1338 = 10'h126 == req_r_addr[14:5] | valid_294; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1339 = 10'h127 == req_r_addr[14:5] | valid_295; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1340 = 10'h128 == req_r_addr[14:5] | valid_296; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1341 = 10'h129 == req_r_addr[14:5] | valid_297; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1342 = 10'h12a == req_r_addr[14:5] | valid_298; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1343 = 10'h12b == req_r_addr[14:5] | valid_299; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1344 = 10'h12c == req_r_addr[14:5] | valid_300; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1345 = 10'h12d == req_r_addr[14:5] | valid_301; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1346 = 10'h12e == req_r_addr[14:5] | valid_302; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1347 = 10'h12f == req_r_addr[14:5] | valid_303; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1348 = 10'h130 == req_r_addr[14:5] | valid_304; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1349 = 10'h131 == req_r_addr[14:5] | valid_305; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1350 = 10'h132 == req_r_addr[14:5] | valid_306; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1351 = 10'h133 == req_r_addr[14:5] | valid_307; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1352 = 10'h134 == req_r_addr[14:5] | valid_308; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1353 = 10'h135 == req_r_addr[14:5] | valid_309; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1354 = 10'h136 == req_r_addr[14:5] | valid_310; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1355 = 10'h137 == req_r_addr[14:5] | valid_311; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1356 = 10'h138 == req_r_addr[14:5] | valid_312; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1357 = 10'h139 == req_r_addr[14:5] | valid_313; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1358 = 10'h13a == req_r_addr[14:5] | valid_314; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1359 = 10'h13b == req_r_addr[14:5] | valid_315; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1360 = 10'h13c == req_r_addr[14:5] | valid_316; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1361 = 10'h13d == req_r_addr[14:5] | valid_317; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1362 = 10'h13e == req_r_addr[14:5] | valid_318; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1363 = 10'h13f == req_r_addr[14:5] | valid_319; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1364 = 10'h140 == req_r_addr[14:5] | valid_320; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1365 = 10'h141 == req_r_addr[14:5] | valid_321; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1366 = 10'h142 == req_r_addr[14:5] | valid_322; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1367 = 10'h143 == req_r_addr[14:5] | valid_323; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1368 = 10'h144 == req_r_addr[14:5] | valid_324; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1369 = 10'h145 == req_r_addr[14:5] | valid_325; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1370 = 10'h146 == req_r_addr[14:5] | valid_326; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1371 = 10'h147 == req_r_addr[14:5] | valid_327; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1372 = 10'h148 == req_r_addr[14:5] | valid_328; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1373 = 10'h149 == req_r_addr[14:5] | valid_329; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1374 = 10'h14a == req_r_addr[14:5] | valid_330; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1375 = 10'h14b == req_r_addr[14:5] | valid_331; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1376 = 10'h14c == req_r_addr[14:5] | valid_332; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1377 = 10'h14d == req_r_addr[14:5] | valid_333; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1378 = 10'h14e == req_r_addr[14:5] | valid_334; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1379 = 10'h14f == req_r_addr[14:5] | valid_335; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1380 = 10'h150 == req_r_addr[14:5] | valid_336; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1381 = 10'h151 == req_r_addr[14:5] | valid_337; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1382 = 10'h152 == req_r_addr[14:5] | valid_338; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1383 = 10'h153 == req_r_addr[14:5] | valid_339; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1384 = 10'h154 == req_r_addr[14:5] | valid_340; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1385 = 10'h155 == req_r_addr[14:5] | valid_341; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1386 = 10'h156 == req_r_addr[14:5] | valid_342; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1387 = 10'h157 == req_r_addr[14:5] | valid_343; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1388 = 10'h158 == req_r_addr[14:5] | valid_344; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1389 = 10'h159 == req_r_addr[14:5] | valid_345; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1390 = 10'h15a == req_r_addr[14:5] | valid_346; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1391 = 10'h15b == req_r_addr[14:5] | valid_347; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1392 = 10'h15c == req_r_addr[14:5] | valid_348; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1393 = 10'h15d == req_r_addr[14:5] | valid_349; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1394 = 10'h15e == req_r_addr[14:5] | valid_350; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1395 = 10'h15f == req_r_addr[14:5] | valid_351; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1396 = 10'h160 == req_r_addr[14:5] | valid_352; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1397 = 10'h161 == req_r_addr[14:5] | valid_353; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1398 = 10'h162 == req_r_addr[14:5] | valid_354; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1399 = 10'h163 == req_r_addr[14:5] | valid_355; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1400 = 10'h164 == req_r_addr[14:5] | valid_356; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1401 = 10'h165 == req_r_addr[14:5] | valid_357; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1402 = 10'h166 == req_r_addr[14:5] | valid_358; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1403 = 10'h167 == req_r_addr[14:5] | valid_359; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1404 = 10'h168 == req_r_addr[14:5] | valid_360; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1405 = 10'h169 == req_r_addr[14:5] | valid_361; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1406 = 10'h16a == req_r_addr[14:5] | valid_362; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1407 = 10'h16b == req_r_addr[14:5] | valid_363; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1408 = 10'h16c == req_r_addr[14:5] | valid_364; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1409 = 10'h16d == req_r_addr[14:5] | valid_365; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1410 = 10'h16e == req_r_addr[14:5] | valid_366; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1411 = 10'h16f == req_r_addr[14:5] | valid_367; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1412 = 10'h170 == req_r_addr[14:5] | valid_368; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1413 = 10'h171 == req_r_addr[14:5] | valid_369; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1414 = 10'h172 == req_r_addr[14:5] | valid_370; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1415 = 10'h173 == req_r_addr[14:5] | valid_371; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1416 = 10'h174 == req_r_addr[14:5] | valid_372; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1417 = 10'h175 == req_r_addr[14:5] | valid_373; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1418 = 10'h176 == req_r_addr[14:5] | valid_374; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1419 = 10'h177 == req_r_addr[14:5] | valid_375; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1420 = 10'h178 == req_r_addr[14:5] | valid_376; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1421 = 10'h179 == req_r_addr[14:5] | valid_377; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1422 = 10'h17a == req_r_addr[14:5] | valid_378; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1423 = 10'h17b == req_r_addr[14:5] | valid_379; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1424 = 10'h17c == req_r_addr[14:5] | valid_380; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1425 = 10'h17d == req_r_addr[14:5] | valid_381; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1426 = 10'h17e == req_r_addr[14:5] | valid_382; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1427 = 10'h17f == req_r_addr[14:5] | valid_383; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1428 = 10'h180 == req_r_addr[14:5] | valid_384; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1429 = 10'h181 == req_r_addr[14:5] | valid_385; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1430 = 10'h182 == req_r_addr[14:5] | valid_386; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1431 = 10'h183 == req_r_addr[14:5] | valid_387; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1432 = 10'h184 == req_r_addr[14:5] | valid_388; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1433 = 10'h185 == req_r_addr[14:5] | valid_389; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1434 = 10'h186 == req_r_addr[14:5] | valid_390; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1435 = 10'h187 == req_r_addr[14:5] | valid_391; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1436 = 10'h188 == req_r_addr[14:5] | valid_392; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1437 = 10'h189 == req_r_addr[14:5] | valid_393; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1438 = 10'h18a == req_r_addr[14:5] | valid_394; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1439 = 10'h18b == req_r_addr[14:5] | valid_395; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1440 = 10'h18c == req_r_addr[14:5] | valid_396; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1441 = 10'h18d == req_r_addr[14:5] | valid_397; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1442 = 10'h18e == req_r_addr[14:5] | valid_398; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1443 = 10'h18f == req_r_addr[14:5] | valid_399; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1444 = 10'h190 == req_r_addr[14:5] | valid_400; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1445 = 10'h191 == req_r_addr[14:5] | valid_401; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1446 = 10'h192 == req_r_addr[14:5] | valid_402; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1447 = 10'h193 == req_r_addr[14:5] | valid_403; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1448 = 10'h194 == req_r_addr[14:5] | valid_404; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1449 = 10'h195 == req_r_addr[14:5] | valid_405; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1450 = 10'h196 == req_r_addr[14:5] | valid_406; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1451 = 10'h197 == req_r_addr[14:5] | valid_407; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1452 = 10'h198 == req_r_addr[14:5] | valid_408; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1453 = 10'h199 == req_r_addr[14:5] | valid_409; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1454 = 10'h19a == req_r_addr[14:5] | valid_410; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1455 = 10'h19b == req_r_addr[14:5] | valid_411; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1456 = 10'h19c == req_r_addr[14:5] | valid_412; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1457 = 10'h19d == req_r_addr[14:5] | valid_413; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1458 = 10'h19e == req_r_addr[14:5] | valid_414; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1459 = 10'h19f == req_r_addr[14:5] | valid_415; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1460 = 10'h1a0 == req_r_addr[14:5] | valid_416; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1461 = 10'h1a1 == req_r_addr[14:5] | valid_417; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1462 = 10'h1a2 == req_r_addr[14:5] | valid_418; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1463 = 10'h1a3 == req_r_addr[14:5] | valid_419; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1464 = 10'h1a4 == req_r_addr[14:5] | valid_420; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1465 = 10'h1a5 == req_r_addr[14:5] | valid_421; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1466 = 10'h1a6 == req_r_addr[14:5] | valid_422; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1467 = 10'h1a7 == req_r_addr[14:5] | valid_423; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1468 = 10'h1a8 == req_r_addr[14:5] | valid_424; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1469 = 10'h1a9 == req_r_addr[14:5] | valid_425; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1470 = 10'h1aa == req_r_addr[14:5] | valid_426; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1471 = 10'h1ab == req_r_addr[14:5] | valid_427; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1472 = 10'h1ac == req_r_addr[14:5] | valid_428; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1473 = 10'h1ad == req_r_addr[14:5] | valid_429; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1474 = 10'h1ae == req_r_addr[14:5] | valid_430; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1475 = 10'h1af == req_r_addr[14:5] | valid_431; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1476 = 10'h1b0 == req_r_addr[14:5] | valid_432; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1477 = 10'h1b1 == req_r_addr[14:5] | valid_433; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1478 = 10'h1b2 == req_r_addr[14:5] | valid_434; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1479 = 10'h1b3 == req_r_addr[14:5] | valid_435; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1480 = 10'h1b4 == req_r_addr[14:5] | valid_436; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1481 = 10'h1b5 == req_r_addr[14:5] | valid_437; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1482 = 10'h1b6 == req_r_addr[14:5] | valid_438; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1483 = 10'h1b7 == req_r_addr[14:5] | valid_439; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1484 = 10'h1b8 == req_r_addr[14:5] | valid_440; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1485 = 10'h1b9 == req_r_addr[14:5] | valid_441; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1486 = 10'h1ba == req_r_addr[14:5] | valid_442; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1487 = 10'h1bb == req_r_addr[14:5] | valid_443; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1488 = 10'h1bc == req_r_addr[14:5] | valid_444; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1489 = 10'h1bd == req_r_addr[14:5] | valid_445; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1490 = 10'h1be == req_r_addr[14:5] | valid_446; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1491 = 10'h1bf == req_r_addr[14:5] | valid_447; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1492 = 10'h1c0 == req_r_addr[14:5] | valid_448; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1493 = 10'h1c1 == req_r_addr[14:5] | valid_449; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1494 = 10'h1c2 == req_r_addr[14:5] | valid_450; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1495 = 10'h1c3 == req_r_addr[14:5] | valid_451; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1496 = 10'h1c4 == req_r_addr[14:5] | valid_452; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1497 = 10'h1c5 == req_r_addr[14:5] | valid_453; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1498 = 10'h1c6 == req_r_addr[14:5] | valid_454; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1499 = 10'h1c7 == req_r_addr[14:5] | valid_455; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1500 = 10'h1c8 == req_r_addr[14:5] | valid_456; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1501 = 10'h1c9 == req_r_addr[14:5] | valid_457; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1502 = 10'h1ca == req_r_addr[14:5] | valid_458; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1503 = 10'h1cb == req_r_addr[14:5] | valid_459; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1504 = 10'h1cc == req_r_addr[14:5] | valid_460; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1505 = 10'h1cd == req_r_addr[14:5] | valid_461; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1506 = 10'h1ce == req_r_addr[14:5] | valid_462; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1507 = 10'h1cf == req_r_addr[14:5] | valid_463; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1508 = 10'h1d0 == req_r_addr[14:5] | valid_464; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1509 = 10'h1d1 == req_r_addr[14:5] | valid_465; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1510 = 10'h1d2 == req_r_addr[14:5] | valid_466; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1511 = 10'h1d3 == req_r_addr[14:5] | valid_467; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1512 = 10'h1d4 == req_r_addr[14:5] | valid_468; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1513 = 10'h1d5 == req_r_addr[14:5] | valid_469; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1514 = 10'h1d6 == req_r_addr[14:5] | valid_470; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1515 = 10'h1d7 == req_r_addr[14:5] | valid_471; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1516 = 10'h1d8 == req_r_addr[14:5] | valid_472; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1517 = 10'h1d9 == req_r_addr[14:5] | valid_473; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1518 = 10'h1da == req_r_addr[14:5] | valid_474; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1519 = 10'h1db == req_r_addr[14:5] | valid_475; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1520 = 10'h1dc == req_r_addr[14:5] | valid_476; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1521 = 10'h1dd == req_r_addr[14:5] | valid_477; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1522 = 10'h1de == req_r_addr[14:5] | valid_478; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1523 = 10'h1df == req_r_addr[14:5] | valid_479; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1524 = 10'h1e0 == req_r_addr[14:5] | valid_480; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1525 = 10'h1e1 == req_r_addr[14:5] | valid_481; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1526 = 10'h1e2 == req_r_addr[14:5] | valid_482; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1527 = 10'h1e3 == req_r_addr[14:5] | valid_483; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1528 = 10'h1e4 == req_r_addr[14:5] | valid_484; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1529 = 10'h1e5 == req_r_addr[14:5] | valid_485; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1530 = 10'h1e6 == req_r_addr[14:5] | valid_486; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1531 = 10'h1e7 == req_r_addr[14:5] | valid_487; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1532 = 10'h1e8 == req_r_addr[14:5] | valid_488; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1533 = 10'h1e9 == req_r_addr[14:5] | valid_489; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1534 = 10'h1ea == req_r_addr[14:5] | valid_490; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1535 = 10'h1eb == req_r_addr[14:5] | valid_491; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1536 = 10'h1ec == req_r_addr[14:5] | valid_492; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1537 = 10'h1ed == req_r_addr[14:5] | valid_493; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1538 = 10'h1ee == req_r_addr[14:5] | valid_494; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1539 = 10'h1ef == req_r_addr[14:5] | valid_495; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1540 = 10'h1f0 == req_r_addr[14:5] | valid_496; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1541 = 10'h1f1 == req_r_addr[14:5] | valid_497; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1542 = 10'h1f2 == req_r_addr[14:5] | valid_498; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1543 = 10'h1f3 == req_r_addr[14:5] | valid_499; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1544 = 10'h1f4 == req_r_addr[14:5] | valid_500; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1545 = 10'h1f5 == req_r_addr[14:5] | valid_501; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1546 = 10'h1f6 == req_r_addr[14:5] | valid_502; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1547 = 10'h1f7 == req_r_addr[14:5] | valid_503; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1548 = 10'h1f8 == req_r_addr[14:5] | valid_504; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1549 = 10'h1f9 == req_r_addr[14:5] | valid_505; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1550 = 10'h1fa == req_r_addr[14:5] | valid_506; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1551 = 10'h1fb == req_r_addr[14:5] | valid_507; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1552 = 10'h1fc == req_r_addr[14:5] | valid_508; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1553 = 10'h1fd == req_r_addr[14:5] | valid_509; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1554 = 10'h1fe == req_r_addr[14:5] | valid_510; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1555 = 10'h1ff == req_r_addr[14:5] | valid_511; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1556 = 10'h200 == req_r_addr[14:5] | valid_512; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1557 = 10'h201 == req_r_addr[14:5] | valid_513; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1558 = 10'h202 == req_r_addr[14:5] | valid_514; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1559 = 10'h203 == req_r_addr[14:5] | valid_515; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1560 = 10'h204 == req_r_addr[14:5] | valid_516; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1561 = 10'h205 == req_r_addr[14:5] | valid_517; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1562 = 10'h206 == req_r_addr[14:5] | valid_518; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1563 = 10'h207 == req_r_addr[14:5] | valid_519; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1564 = 10'h208 == req_r_addr[14:5] | valid_520; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1565 = 10'h209 == req_r_addr[14:5] | valid_521; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1566 = 10'h20a == req_r_addr[14:5] | valid_522; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1567 = 10'h20b == req_r_addr[14:5] | valid_523; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1568 = 10'h20c == req_r_addr[14:5] | valid_524; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1569 = 10'h20d == req_r_addr[14:5] | valid_525; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1570 = 10'h20e == req_r_addr[14:5] | valid_526; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1571 = 10'h20f == req_r_addr[14:5] | valid_527; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1572 = 10'h210 == req_r_addr[14:5] | valid_528; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1573 = 10'h211 == req_r_addr[14:5] | valid_529; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1574 = 10'h212 == req_r_addr[14:5] | valid_530; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1575 = 10'h213 == req_r_addr[14:5] | valid_531; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1576 = 10'h214 == req_r_addr[14:5] | valid_532; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1577 = 10'h215 == req_r_addr[14:5] | valid_533; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1578 = 10'h216 == req_r_addr[14:5] | valid_534; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1579 = 10'h217 == req_r_addr[14:5] | valid_535; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1580 = 10'h218 == req_r_addr[14:5] | valid_536; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1581 = 10'h219 == req_r_addr[14:5] | valid_537; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1582 = 10'h21a == req_r_addr[14:5] | valid_538; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1583 = 10'h21b == req_r_addr[14:5] | valid_539; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1584 = 10'h21c == req_r_addr[14:5] | valid_540; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1585 = 10'h21d == req_r_addr[14:5] | valid_541; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1586 = 10'h21e == req_r_addr[14:5] | valid_542; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1587 = 10'h21f == req_r_addr[14:5] | valid_543; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1588 = 10'h220 == req_r_addr[14:5] | valid_544; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1589 = 10'h221 == req_r_addr[14:5] | valid_545; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1590 = 10'h222 == req_r_addr[14:5] | valid_546; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1591 = 10'h223 == req_r_addr[14:5] | valid_547; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1592 = 10'h224 == req_r_addr[14:5] | valid_548; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1593 = 10'h225 == req_r_addr[14:5] | valid_549; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1594 = 10'h226 == req_r_addr[14:5] | valid_550; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1595 = 10'h227 == req_r_addr[14:5] | valid_551; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1596 = 10'h228 == req_r_addr[14:5] | valid_552; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1597 = 10'h229 == req_r_addr[14:5] | valid_553; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1598 = 10'h22a == req_r_addr[14:5] | valid_554; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1599 = 10'h22b == req_r_addr[14:5] | valid_555; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1600 = 10'h22c == req_r_addr[14:5] | valid_556; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1601 = 10'h22d == req_r_addr[14:5] | valid_557; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1602 = 10'h22e == req_r_addr[14:5] | valid_558; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1603 = 10'h22f == req_r_addr[14:5] | valid_559; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1604 = 10'h230 == req_r_addr[14:5] | valid_560; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1605 = 10'h231 == req_r_addr[14:5] | valid_561; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1606 = 10'h232 == req_r_addr[14:5] | valid_562; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1607 = 10'h233 == req_r_addr[14:5] | valid_563; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1608 = 10'h234 == req_r_addr[14:5] | valid_564; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1609 = 10'h235 == req_r_addr[14:5] | valid_565; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1610 = 10'h236 == req_r_addr[14:5] | valid_566; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1611 = 10'h237 == req_r_addr[14:5] | valid_567; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1612 = 10'h238 == req_r_addr[14:5] | valid_568; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1613 = 10'h239 == req_r_addr[14:5] | valid_569; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1614 = 10'h23a == req_r_addr[14:5] | valid_570; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1615 = 10'h23b == req_r_addr[14:5] | valid_571; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1616 = 10'h23c == req_r_addr[14:5] | valid_572; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1617 = 10'h23d == req_r_addr[14:5] | valid_573; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1618 = 10'h23e == req_r_addr[14:5] | valid_574; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1619 = 10'h23f == req_r_addr[14:5] | valid_575; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1620 = 10'h240 == req_r_addr[14:5] | valid_576; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1621 = 10'h241 == req_r_addr[14:5] | valid_577; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1622 = 10'h242 == req_r_addr[14:5] | valid_578; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1623 = 10'h243 == req_r_addr[14:5] | valid_579; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1624 = 10'h244 == req_r_addr[14:5] | valid_580; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1625 = 10'h245 == req_r_addr[14:5] | valid_581; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1626 = 10'h246 == req_r_addr[14:5] | valid_582; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1627 = 10'h247 == req_r_addr[14:5] | valid_583; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1628 = 10'h248 == req_r_addr[14:5] | valid_584; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1629 = 10'h249 == req_r_addr[14:5] | valid_585; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1630 = 10'h24a == req_r_addr[14:5] | valid_586; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1631 = 10'h24b == req_r_addr[14:5] | valid_587; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1632 = 10'h24c == req_r_addr[14:5] | valid_588; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1633 = 10'h24d == req_r_addr[14:5] | valid_589; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1634 = 10'h24e == req_r_addr[14:5] | valid_590; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1635 = 10'h24f == req_r_addr[14:5] | valid_591; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1636 = 10'h250 == req_r_addr[14:5] | valid_592; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1637 = 10'h251 == req_r_addr[14:5] | valid_593; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1638 = 10'h252 == req_r_addr[14:5] | valid_594; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1639 = 10'h253 == req_r_addr[14:5] | valid_595; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1640 = 10'h254 == req_r_addr[14:5] | valid_596; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1641 = 10'h255 == req_r_addr[14:5] | valid_597; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1642 = 10'h256 == req_r_addr[14:5] | valid_598; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1643 = 10'h257 == req_r_addr[14:5] | valid_599; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1644 = 10'h258 == req_r_addr[14:5] | valid_600; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1645 = 10'h259 == req_r_addr[14:5] | valid_601; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1646 = 10'h25a == req_r_addr[14:5] | valid_602; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1647 = 10'h25b == req_r_addr[14:5] | valid_603; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1648 = 10'h25c == req_r_addr[14:5] | valid_604; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1649 = 10'h25d == req_r_addr[14:5] | valid_605; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1650 = 10'h25e == req_r_addr[14:5] | valid_606; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1651 = 10'h25f == req_r_addr[14:5] | valid_607; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1652 = 10'h260 == req_r_addr[14:5] | valid_608; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1653 = 10'h261 == req_r_addr[14:5] | valid_609; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1654 = 10'h262 == req_r_addr[14:5] | valid_610; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1655 = 10'h263 == req_r_addr[14:5] | valid_611; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1656 = 10'h264 == req_r_addr[14:5] | valid_612; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1657 = 10'h265 == req_r_addr[14:5] | valid_613; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1658 = 10'h266 == req_r_addr[14:5] | valid_614; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1659 = 10'h267 == req_r_addr[14:5] | valid_615; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1660 = 10'h268 == req_r_addr[14:5] | valid_616; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1661 = 10'h269 == req_r_addr[14:5] | valid_617; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1662 = 10'h26a == req_r_addr[14:5] | valid_618; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1663 = 10'h26b == req_r_addr[14:5] | valid_619; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1664 = 10'h26c == req_r_addr[14:5] | valid_620; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1665 = 10'h26d == req_r_addr[14:5] | valid_621; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1666 = 10'h26e == req_r_addr[14:5] | valid_622; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1667 = 10'h26f == req_r_addr[14:5] | valid_623; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1668 = 10'h270 == req_r_addr[14:5] | valid_624; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1669 = 10'h271 == req_r_addr[14:5] | valid_625; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1670 = 10'h272 == req_r_addr[14:5] | valid_626; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1671 = 10'h273 == req_r_addr[14:5] | valid_627; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1672 = 10'h274 == req_r_addr[14:5] | valid_628; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1673 = 10'h275 == req_r_addr[14:5] | valid_629; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1674 = 10'h276 == req_r_addr[14:5] | valid_630; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1675 = 10'h277 == req_r_addr[14:5] | valid_631; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1676 = 10'h278 == req_r_addr[14:5] | valid_632; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1677 = 10'h279 == req_r_addr[14:5] | valid_633; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1678 = 10'h27a == req_r_addr[14:5] | valid_634; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1679 = 10'h27b == req_r_addr[14:5] | valid_635; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1680 = 10'h27c == req_r_addr[14:5] | valid_636; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1681 = 10'h27d == req_r_addr[14:5] | valid_637; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1682 = 10'h27e == req_r_addr[14:5] | valid_638; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1683 = 10'h27f == req_r_addr[14:5] | valid_639; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1684 = 10'h280 == req_r_addr[14:5] | valid_640; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1685 = 10'h281 == req_r_addr[14:5] | valid_641; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1686 = 10'h282 == req_r_addr[14:5] | valid_642; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1687 = 10'h283 == req_r_addr[14:5] | valid_643; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1688 = 10'h284 == req_r_addr[14:5] | valid_644; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1689 = 10'h285 == req_r_addr[14:5] | valid_645; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1690 = 10'h286 == req_r_addr[14:5] | valid_646; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1691 = 10'h287 == req_r_addr[14:5] | valid_647; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1692 = 10'h288 == req_r_addr[14:5] | valid_648; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1693 = 10'h289 == req_r_addr[14:5] | valid_649; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1694 = 10'h28a == req_r_addr[14:5] | valid_650; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1695 = 10'h28b == req_r_addr[14:5] | valid_651; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1696 = 10'h28c == req_r_addr[14:5] | valid_652; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1697 = 10'h28d == req_r_addr[14:5] | valid_653; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1698 = 10'h28e == req_r_addr[14:5] | valid_654; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1699 = 10'h28f == req_r_addr[14:5] | valid_655; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1700 = 10'h290 == req_r_addr[14:5] | valid_656; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1701 = 10'h291 == req_r_addr[14:5] | valid_657; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1702 = 10'h292 == req_r_addr[14:5] | valid_658; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1703 = 10'h293 == req_r_addr[14:5] | valid_659; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1704 = 10'h294 == req_r_addr[14:5] | valid_660; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1705 = 10'h295 == req_r_addr[14:5] | valid_661; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1706 = 10'h296 == req_r_addr[14:5] | valid_662; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1707 = 10'h297 == req_r_addr[14:5] | valid_663; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1708 = 10'h298 == req_r_addr[14:5] | valid_664; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1709 = 10'h299 == req_r_addr[14:5] | valid_665; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1710 = 10'h29a == req_r_addr[14:5] | valid_666; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1711 = 10'h29b == req_r_addr[14:5] | valid_667; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1712 = 10'h29c == req_r_addr[14:5] | valid_668; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1713 = 10'h29d == req_r_addr[14:5] | valid_669; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1714 = 10'h29e == req_r_addr[14:5] | valid_670; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1715 = 10'h29f == req_r_addr[14:5] | valid_671; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1716 = 10'h2a0 == req_r_addr[14:5] | valid_672; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1717 = 10'h2a1 == req_r_addr[14:5] | valid_673; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1718 = 10'h2a2 == req_r_addr[14:5] | valid_674; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1719 = 10'h2a3 == req_r_addr[14:5] | valid_675; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1720 = 10'h2a4 == req_r_addr[14:5] | valid_676; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1721 = 10'h2a5 == req_r_addr[14:5] | valid_677; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1722 = 10'h2a6 == req_r_addr[14:5] | valid_678; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1723 = 10'h2a7 == req_r_addr[14:5] | valid_679; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1724 = 10'h2a8 == req_r_addr[14:5] | valid_680; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1725 = 10'h2a9 == req_r_addr[14:5] | valid_681; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1726 = 10'h2aa == req_r_addr[14:5] | valid_682; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1727 = 10'h2ab == req_r_addr[14:5] | valid_683; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1728 = 10'h2ac == req_r_addr[14:5] | valid_684; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1729 = 10'h2ad == req_r_addr[14:5] | valid_685; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1730 = 10'h2ae == req_r_addr[14:5] | valid_686; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1731 = 10'h2af == req_r_addr[14:5] | valid_687; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1732 = 10'h2b0 == req_r_addr[14:5] | valid_688; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1733 = 10'h2b1 == req_r_addr[14:5] | valid_689; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1734 = 10'h2b2 == req_r_addr[14:5] | valid_690; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1735 = 10'h2b3 == req_r_addr[14:5] | valid_691; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1736 = 10'h2b4 == req_r_addr[14:5] | valid_692; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1737 = 10'h2b5 == req_r_addr[14:5] | valid_693; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1738 = 10'h2b6 == req_r_addr[14:5] | valid_694; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1739 = 10'h2b7 == req_r_addr[14:5] | valid_695; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1740 = 10'h2b8 == req_r_addr[14:5] | valid_696; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1741 = 10'h2b9 == req_r_addr[14:5] | valid_697; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1742 = 10'h2ba == req_r_addr[14:5] | valid_698; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1743 = 10'h2bb == req_r_addr[14:5] | valid_699; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1744 = 10'h2bc == req_r_addr[14:5] | valid_700; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1745 = 10'h2bd == req_r_addr[14:5] | valid_701; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1746 = 10'h2be == req_r_addr[14:5] | valid_702; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1747 = 10'h2bf == req_r_addr[14:5] | valid_703; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1748 = 10'h2c0 == req_r_addr[14:5] | valid_704; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1749 = 10'h2c1 == req_r_addr[14:5] | valid_705; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1750 = 10'h2c2 == req_r_addr[14:5] | valid_706; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1751 = 10'h2c3 == req_r_addr[14:5] | valid_707; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1752 = 10'h2c4 == req_r_addr[14:5] | valid_708; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1753 = 10'h2c5 == req_r_addr[14:5] | valid_709; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1754 = 10'h2c6 == req_r_addr[14:5] | valid_710; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1755 = 10'h2c7 == req_r_addr[14:5] | valid_711; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1756 = 10'h2c8 == req_r_addr[14:5] | valid_712; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1757 = 10'h2c9 == req_r_addr[14:5] | valid_713; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1758 = 10'h2ca == req_r_addr[14:5] | valid_714; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1759 = 10'h2cb == req_r_addr[14:5] | valid_715; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1760 = 10'h2cc == req_r_addr[14:5] | valid_716; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1761 = 10'h2cd == req_r_addr[14:5] | valid_717; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1762 = 10'h2ce == req_r_addr[14:5] | valid_718; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1763 = 10'h2cf == req_r_addr[14:5] | valid_719; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1764 = 10'h2d0 == req_r_addr[14:5] | valid_720; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1765 = 10'h2d1 == req_r_addr[14:5] | valid_721; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1766 = 10'h2d2 == req_r_addr[14:5] | valid_722; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1767 = 10'h2d3 == req_r_addr[14:5] | valid_723; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1768 = 10'h2d4 == req_r_addr[14:5] | valid_724; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1769 = 10'h2d5 == req_r_addr[14:5] | valid_725; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1770 = 10'h2d6 == req_r_addr[14:5] | valid_726; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1771 = 10'h2d7 == req_r_addr[14:5] | valid_727; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1772 = 10'h2d8 == req_r_addr[14:5] | valid_728; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1773 = 10'h2d9 == req_r_addr[14:5] | valid_729; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1774 = 10'h2da == req_r_addr[14:5] | valid_730; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1775 = 10'h2db == req_r_addr[14:5] | valid_731; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1776 = 10'h2dc == req_r_addr[14:5] | valid_732; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1777 = 10'h2dd == req_r_addr[14:5] | valid_733; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1778 = 10'h2de == req_r_addr[14:5] | valid_734; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1779 = 10'h2df == req_r_addr[14:5] | valid_735; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1780 = 10'h2e0 == req_r_addr[14:5] | valid_736; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1781 = 10'h2e1 == req_r_addr[14:5] | valid_737; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1782 = 10'h2e2 == req_r_addr[14:5] | valid_738; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1783 = 10'h2e3 == req_r_addr[14:5] | valid_739; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1784 = 10'h2e4 == req_r_addr[14:5] | valid_740; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1785 = 10'h2e5 == req_r_addr[14:5] | valid_741; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1786 = 10'h2e6 == req_r_addr[14:5] | valid_742; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1787 = 10'h2e7 == req_r_addr[14:5] | valid_743; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1788 = 10'h2e8 == req_r_addr[14:5] | valid_744; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1789 = 10'h2e9 == req_r_addr[14:5] | valid_745; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1790 = 10'h2ea == req_r_addr[14:5] | valid_746; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1791 = 10'h2eb == req_r_addr[14:5] | valid_747; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1792 = 10'h2ec == req_r_addr[14:5] | valid_748; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1793 = 10'h2ed == req_r_addr[14:5] | valid_749; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1794 = 10'h2ee == req_r_addr[14:5] | valid_750; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1795 = 10'h2ef == req_r_addr[14:5] | valid_751; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1796 = 10'h2f0 == req_r_addr[14:5] | valid_752; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1797 = 10'h2f1 == req_r_addr[14:5] | valid_753; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1798 = 10'h2f2 == req_r_addr[14:5] | valid_754; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1799 = 10'h2f3 == req_r_addr[14:5] | valid_755; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1800 = 10'h2f4 == req_r_addr[14:5] | valid_756; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1801 = 10'h2f5 == req_r_addr[14:5] | valid_757; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1802 = 10'h2f6 == req_r_addr[14:5] | valid_758; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1803 = 10'h2f7 == req_r_addr[14:5] | valid_759; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1804 = 10'h2f8 == req_r_addr[14:5] | valid_760; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1805 = 10'h2f9 == req_r_addr[14:5] | valid_761; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1806 = 10'h2fa == req_r_addr[14:5] | valid_762; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1807 = 10'h2fb == req_r_addr[14:5] | valid_763; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1808 = 10'h2fc == req_r_addr[14:5] | valid_764; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1809 = 10'h2fd == req_r_addr[14:5] | valid_765; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1810 = 10'h2fe == req_r_addr[14:5] | valid_766; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1811 = 10'h2ff == req_r_addr[14:5] | valid_767; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1812 = 10'h300 == req_r_addr[14:5] | valid_768; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1813 = 10'h301 == req_r_addr[14:5] | valid_769; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1814 = 10'h302 == req_r_addr[14:5] | valid_770; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1815 = 10'h303 == req_r_addr[14:5] | valid_771; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1816 = 10'h304 == req_r_addr[14:5] | valid_772; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1817 = 10'h305 == req_r_addr[14:5] | valid_773; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1818 = 10'h306 == req_r_addr[14:5] | valid_774; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1819 = 10'h307 == req_r_addr[14:5] | valid_775; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1820 = 10'h308 == req_r_addr[14:5] | valid_776; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1821 = 10'h309 == req_r_addr[14:5] | valid_777; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1822 = 10'h30a == req_r_addr[14:5] | valid_778; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1823 = 10'h30b == req_r_addr[14:5] | valid_779; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1824 = 10'h30c == req_r_addr[14:5] | valid_780; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1825 = 10'h30d == req_r_addr[14:5] | valid_781; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1826 = 10'h30e == req_r_addr[14:5] | valid_782; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1827 = 10'h30f == req_r_addr[14:5] | valid_783; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1828 = 10'h310 == req_r_addr[14:5] | valid_784; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1829 = 10'h311 == req_r_addr[14:5] | valid_785; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1830 = 10'h312 == req_r_addr[14:5] | valid_786; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1831 = 10'h313 == req_r_addr[14:5] | valid_787; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1832 = 10'h314 == req_r_addr[14:5] | valid_788; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1833 = 10'h315 == req_r_addr[14:5] | valid_789; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1834 = 10'h316 == req_r_addr[14:5] | valid_790; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1835 = 10'h317 == req_r_addr[14:5] | valid_791; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1836 = 10'h318 == req_r_addr[14:5] | valid_792; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1837 = 10'h319 == req_r_addr[14:5] | valid_793; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1838 = 10'h31a == req_r_addr[14:5] | valid_794; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1839 = 10'h31b == req_r_addr[14:5] | valid_795; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1840 = 10'h31c == req_r_addr[14:5] | valid_796; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1841 = 10'h31d == req_r_addr[14:5] | valid_797; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1842 = 10'h31e == req_r_addr[14:5] | valid_798; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1843 = 10'h31f == req_r_addr[14:5] | valid_799; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1844 = 10'h320 == req_r_addr[14:5] | valid_800; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1845 = 10'h321 == req_r_addr[14:5] | valid_801; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1846 = 10'h322 == req_r_addr[14:5] | valid_802; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1847 = 10'h323 == req_r_addr[14:5] | valid_803; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1848 = 10'h324 == req_r_addr[14:5] | valid_804; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1849 = 10'h325 == req_r_addr[14:5] | valid_805; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1850 = 10'h326 == req_r_addr[14:5] | valid_806; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1851 = 10'h327 == req_r_addr[14:5] | valid_807; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1852 = 10'h328 == req_r_addr[14:5] | valid_808; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1853 = 10'h329 == req_r_addr[14:5] | valid_809; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1854 = 10'h32a == req_r_addr[14:5] | valid_810; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1855 = 10'h32b == req_r_addr[14:5] | valid_811; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1856 = 10'h32c == req_r_addr[14:5] | valid_812; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1857 = 10'h32d == req_r_addr[14:5] | valid_813; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1858 = 10'h32e == req_r_addr[14:5] | valid_814; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1859 = 10'h32f == req_r_addr[14:5] | valid_815; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1860 = 10'h330 == req_r_addr[14:5] | valid_816; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1861 = 10'h331 == req_r_addr[14:5] | valid_817; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1862 = 10'h332 == req_r_addr[14:5] | valid_818; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1863 = 10'h333 == req_r_addr[14:5] | valid_819; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1864 = 10'h334 == req_r_addr[14:5] | valid_820; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1865 = 10'h335 == req_r_addr[14:5] | valid_821; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1866 = 10'h336 == req_r_addr[14:5] | valid_822; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1867 = 10'h337 == req_r_addr[14:5] | valid_823; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1868 = 10'h338 == req_r_addr[14:5] | valid_824; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1869 = 10'h339 == req_r_addr[14:5] | valid_825; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1870 = 10'h33a == req_r_addr[14:5] | valid_826; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1871 = 10'h33b == req_r_addr[14:5] | valid_827; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1872 = 10'h33c == req_r_addr[14:5] | valid_828; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1873 = 10'h33d == req_r_addr[14:5] | valid_829; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1874 = 10'h33e == req_r_addr[14:5] | valid_830; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1875 = 10'h33f == req_r_addr[14:5] | valid_831; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1876 = 10'h340 == req_r_addr[14:5] | valid_832; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1877 = 10'h341 == req_r_addr[14:5] | valid_833; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1878 = 10'h342 == req_r_addr[14:5] | valid_834; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1879 = 10'h343 == req_r_addr[14:5] | valid_835; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1880 = 10'h344 == req_r_addr[14:5] | valid_836; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1881 = 10'h345 == req_r_addr[14:5] | valid_837; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1882 = 10'h346 == req_r_addr[14:5] | valid_838; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1883 = 10'h347 == req_r_addr[14:5] | valid_839; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1884 = 10'h348 == req_r_addr[14:5] | valid_840; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1885 = 10'h349 == req_r_addr[14:5] | valid_841; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1886 = 10'h34a == req_r_addr[14:5] | valid_842; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1887 = 10'h34b == req_r_addr[14:5] | valid_843; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1888 = 10'h34c == req_r_addr[14:5] | valid_844; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1889 = 10'h34d == req_r_addr[14:5] | valid_845; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1890 = 10'h34e == req_r_addr[14:5] | valid_846; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1891 = 10'h34f == req_r_addr[14:5] | valid_847; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1892 = 10'h350 == req_r_addr[14:5] | valid_848; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1893 = 10'h351 == req_r_addr[14:5] | valid_849; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1894 = 10'h352 == req_r_addr[14:5] | valid_850; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1895 = 10'h353 == req_r_addr[14:5] | valid_851; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1896 = 10'h354 == req_r_addr[14:5] | valid_852; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1897 = 10'h355 == req_r_addr[14:5] | valid_853; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1898 = 10'h356 == req_r_addr[14:5] | valid_854; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1899 = 10'h357 == req_r_addr[14:5] | valid_855; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1900 = 10'h358 == req_r_addr[14:5] | valid_856; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1901 = 10'h359 == req_r_addr[14:5] | valid_857; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1902 = 10'h35a == req_r_addr[14:5] | valid_858; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1903 = 10'h35b == req_r_addr[14:5] | valid_859; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1904 = 10'h35c == req_r_addr[14:5] | valid_860; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1905 = 10'h35d == req_r_addr[14:5] | valid_861; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1906 = 10'h35e == req_r_addr[14:5] | valid_862; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1907 = 10'h35f == req_r_addr[14:5] | valid_863; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1908 = 10'h360 == req_r_addr[14:5] | valid_864; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1909 = 10'h361 == req_r_addr[14:5] | valid_865; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1910 = 10'h362 == req_r_addr[14:5] | valid_866; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1911 = 10'h363 == req_r_addr[14:5] | valid_867; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1912 = 10'h364 == req_r_addr[14:5] | valid_868; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1913 = 10'h365 == req_r_addr[14:5] | valid_869; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1914 = 10'h366 == req_r_addr[14:5] | valid_870; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1915 = 10'h367 == req_r_addr[14:5] | valid_871; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1916 = 10'h368 == req_r_addr[14:5] | valid_872; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1917 = 10'h369 == req_r_addr[14:5] | valid_873; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1918 = 10'h36a == req_r_addr[14:5] | valid_874; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1919 = 10'h36b == req_r_addr[14:5] | valid_875; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1920 = 10'h36c == req_r_addr[14:5] | valid_876; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1921 = 10'h36d == req_r_addr[14:5] | valid_877; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1922 = 10'h36e == req_r_addr[14:5] | valid_878; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1923 = 10'h36f == req_r_addr[14:5] | valid_879; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1924 = 10'h370 == req_r_addr[14:5] | valid_880; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1925 = 10'h371 == req_r_addr[14:5] | valid_881; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1926 = 10'h372 == req_r_addr[14:5] | valid_882; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1927 = 10'h373 == req_r_addr[14:5] | valid_883; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1928 = 10'h374 == req_r_addr[14:5] | valid_884; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1929 = 10'h375 == req_r_addr[14:5] | valid_885; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1930 = 10'h376 == req_r_addr[14:5] | valid_886; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1931 = 10'h377 == req_r_addr[14:5] | valid_887; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1932 = 10'h378 == req_r_addr[14:5] | valid_888; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1933 = 10'h379 == req_r_addr[14:5] | valid_889; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1934 = 10'h37a == req_r_addr[14:5] | valid_890; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1935 = 10'h37b == req_r_addr[14:5] | valid_891; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1936 = 10'h37c == req_r_addr[14:5] | valid_892; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1937 = 10'h37d == req_r_addr[14:5] | valid_893; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1938 = 10'h37e == req_r_addr[14:5] | valid_894; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1939 = 10'h37f == req_r_addr[14:5] | valid_895; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1940 = 10'h380 == req_r_addr[14:5] | valid_896; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1941 = 10'h381 == req_r_addr[14:5] | valid_897; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1942 = 10'h382 == req_r_addr[14:5] | valid_898; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1943 = 10'h383 == req_r_addr[14:5] | valid_899; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1944 = 10'h384 == req_r_addr[14:5] | valid_900; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1945 = 10'h385 == req_r_addr[14:5] | valid_901; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1946 = 10'h386 == req_r_addr[14:5] | valid_902; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1947 = 10'h387 == req_r_addr[14:5] | valid_903; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1948 = 10'h388 == req_r_addr[14:5] | valid_904; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1949 = 10'h389 == req_r_addr[14:5] | valid_905; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1950 = 10'h38a == req_r_addr[14:5] | valid_906; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1951 = 10'h38b == req_r_addr[14:5] | valid_907; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1952 = 10'h38c == req_r_addr[14:5] | valid_908; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1953 = 10'h38d == req_r_addr[14:5] | valid_909; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1954 = 10'h38e == req_r_addr[14:5] | valid_910; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1955 = 10'h38f == req_r_addr[14:5] | valid_911; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1956 = 10'h390 == req_r_addr[14:5] | valid_912; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1957 = 10'h391 == req_r_addr[14:5] | valid_913; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1958 = 10'h392 == req_r_addr[14:5] | valid_914; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1959 = 10'h393 == req_r_addr[14:5] | valid_915; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1960 = 10'h394 == req_r_addr[14:5] | valid_916; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1961 = 10'h395 == req_r_addr[14:5] | valid_917; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1962 = 10'h396 == req_r_addr[14:5] | valid_918; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1963 = 10'h397 == req_r_addr[14:5] | valid_919; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1964 = 10'h398 == req_r_addr[14:5] | valid_920; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1965 = 10'h399 == req_r_addr[14:5] | valid_921; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1966 = 10'h39a == req_r_addr[14:5] | valid_922; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1967 = 10'h39b == req_r_addr[14:5] | valid_923; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1968 = 10'h39c == req_r_addr[14:5] | valid_924; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1969 = 10'h39d == req_r_addr[14:5] | valid_925; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1970 = 10'h39e == req_r_addr[14:5] | valid_926; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1971 = 10'h39f == req_r_addr[14:5] | valid_927; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1972 = 10'h3a0 == req_r_addr[14:5] | valid_928; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1973 = 10'h3a1 == req_r_addr[14:5] | valid_929; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1974 = 10'h3a2 == req_r_addr[14:5] | valid_930; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1975 = 10'h3a3 == req_r_addr[14:5] | valid_931; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1976 = 10'h3a4 == req_r_addr[14:5] | valid_932; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1977 = 10'h3a5 == req_r_addr[14:5] | valid_933; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1978 = 10'h3a6 == req_r_addr[14:5] | valid_934; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1979 = 10'h3a7 == req_r_addr[14:5] | valid_935; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1980 = 10'h3a8 == req_r_addr[14:5] | valid_936; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1981 = 10'h3a9 == req_r_addr[14:5] | valid_937; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1982 = 10'h3aa == req_r_addr[14:5] | valid_938; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1983 = 10'h3ab == req_r_addr[14:5] | valid_939; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1984 = 10'h3ac == req_r_addr[14:5] | valid_940; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1985 = 10'h3ad == req_r_addr[14:5] | valid_941; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1986 = 10'h3ae == req_r_addr[14:5] | valid_942; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1987 = 10'h3af == req_r_addr[14:5] | valid_943; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1988 = 10'h3b0 == req_r_addr[14:5] | valid_944; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1989 = 10'h3b1 == req_r_addr[14:5] | valid_945; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1990 = 10'h3b2 == req_r_addr[14:5] | valid_946; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1991 = 10'h3b3 == req_r_addr[14:5] | valid_947; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1992 = 10'h3b4 == req_r_addr[14:5] | valid_948; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1993 = 10'h3b5 == req_r_addr[14:5] | valid_949; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1994 = 10'h3b6 == req_r_addr[14:5] | valid_950; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1995 = 10'h3b7 == req_r_addr[14:5] | valid_951; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1996 = 10'h3b8 == req_r_addr[14:5] | valid_952; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1997 = 10'h3b9 == req_r_addr[14:5] | valid_953; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1998 = 10'h3ba == req_r_addr[14:5] | valid_954; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_1999 = 10'h3bb == req_r_addr[14:5] | valid_955; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2000 = 10'h3bc == req_r_addr[14:5] | valid_956; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2001 = 10'h3bd == req_r_addr[14:5] | valid_957; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2002 = 10'h3be == req_r_addr[14:5] | valid_958; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2003 = 10'h3bf == req_r_addr[14:5] | valid_959; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2004 = 10'h3c0 == req_r_addr[14:5] | valid_960; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2005 = 10'h3c1 == req_r_addr[14:5] | valid_961; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2006 = 10'h3c2 == req_r_addr[14:5] | valid_962; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2007 = 10'h3c3 == req_r_addr[14:5] | valid_963; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2008 = 10'h3c4 == req_r_addr[14:5] | valid_964; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2009 = 10'h3c5 == req_r_addr[14:5] | valid_965; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2010 = 10'h3c6 == req_r_addr[14:5] | valid_966; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2011 = 10'h3c7 == req_r_addr[14:5] | valid_967; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2012 = 10'h3c8 == req_r_addr[14:5] | valid_968; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2013 = 10'h3c9 == req_r_addr[14:5] | valid_969; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2014 = 10'h3ca == req_r_addr[14:5] | valid_970; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2015 = 10'h3cb == req_r_addr[14:5] | valid_971; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2016 = 10'h3cc == req_r_addr[14:5] | valid_972; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2017 = 10'h3cd == req_r_addr[14:5] | valid_973; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2018 = 10'h3ce == req_r_addr[14:5] | valid_974; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2019 = 10'h3cf == req_r_addr[14:5] | valid_975; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2020 = 10'h3d0 == req_r_addr[14:5] | valid_976; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2021 = 10'h3d1 == req_r_addr[14:5] | valid_977; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2022 = 10'h3d2 == req_r_addr[14:5] | valid_978; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2023 = 10'h3d3 == req_r_addr[14:5] | valid_979; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2024 = 10'h3d4 == req_r_addr[14:5] | valid_980; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2025 = 10'h3d5 == req_r_addr[14:5] | valid_981; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2026 = 10'h3d6 == req_r_addr[14:5] | valid_982; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2027 = 10'h3d7 == req_r_addr[14:5] | valid_983; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2028 = 10'h3d8 == req_r_addr[14:5] | valid_984; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2029 = 10'h3d9 == req_r_addr[14:5] | valid_985; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2030 = 10'h3da == req_r_addr[14:5] | valid_986; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2031 = 10'h3db == req_r_addr[14:5] | valid_987; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2032 = 10'h3dc == req_r_addr[14:5] | valid_988; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2033 = 10'h3dd == req_r_addr[14:5] | valid_989; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2034 = 10'h3de == req_r_addr[14:5] | valid_990; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2035 = 10'h3df == req_r_addr[14:5] | valid_991; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2036 = 10'h3e0 == req_r_addr[14:5] | valid_992; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2037 = 10'h3e1 == req_r_addr[14:5] | valid_993; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2038 = 10'h3e2 == req_r_addr[14:5] | valid_994; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2039 = 10'h3e3 == req_r_addr[14:5] | valid_995; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2040 = 10'h3e4 == req_r_addr[14:5] | valid_996; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2041 = 10'h3e5 == req_r_addr[14:5] | valid_997; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2042 = 10'h3e6 == req_r_addr[14:5] | valid_998; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2043 = 10'h3e7 == req_r_addr[14:5] | valid_999; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2044 = 10'h3e8 == req_r_addr[14:5] | valid_1000; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2045 = 10'h3e9 == req_r_addr[14:5] | valid_1001; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2046 = 10'h3ea == req_r_addr[14:5] | valid_1002; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2047 = 10'h3eb == req_r_addr[14:5] | valid_1003; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2048 = 10'h3ec == req_r_addr[14:5] | valid_1004; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2049 = 10'h3ed == req_r_addr[14:5] | valid_1005; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2050 = 10'h3ee == req_r_addr[14:5] | valid_1006; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2051 = 10'h3ef == req_r_addr[14:5] | valid_1007; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2052 = 10'h3f0 == req_r_addr[14:5] | valid_1008; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2053 = 10'h3f1 == req_r_addr[14:5] | valid_1009; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2054 = 10'h3f2 == req_r_addr[14:5] | valid_1010; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2055 = 10'h3f3 == req_r_addr[14:5] | valid_1011; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2056 = 10'h3f4 == req_r_addr[14:5] | valid_1012; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2057 = 10'h3f5 == req_r_addr[14:5] | valid_1013; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2058 = 10'h3f6 == req_r_addr[14:5] | valid_1014; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2059 = 10'h3f7 == req_r_addr[14:5] | valid_1015; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2060 = 10'h3f8 == req_r_addr[14:5] | valid_1016; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2061 = 10'h3f9 == req_r_addr[14:5] | valid_1017; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2062 = 10'h3fa == req_r_addr[14:5] | valid_1018; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2063 = 10'h3fb == req_r_addr[14:5] | valid_1019; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2064 = 10'h3fc == req_r_addr[14:5] | valid_1020; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2065 = 10'h3fd == req_r_addr[14:5] | valid_1021; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2066 = 10'h3fe == req_r_addr[14:5] | valid_1022; // @[ICache.scala 128:{33,33} 51:22]
  wire  _GEN_2067 = 10'h3ff == req_r_addr[14:5] | valid_1023; // @[ICache.scala 128:{33,33} 51:22]
  wire [63:0] _refill_data_T_6 = 2'h1 == req_r_addr[4:3] ? wdata[127:64] : wdata[63:0]; // @[Mux.scala 81:58]
  wire [63:0] _refill_data_T_8 = 2'h2 == req_r_addr[4:3] ? wdata[191:128] : _refill_data_T_6; // @[Mux.scala 81:58]
  wire [63:0] refill_data = 2'h3 == req_r_addr[4:3] ? wdata[255:192] : _refill_data_T_8; // @[Mux.scala 81:58]
  reg [1:0] source; // @[Counter.scala 61:40]
  wire [1:0] _source_wrap_value_T_1 = source + 2'h1; // @[Counter.scala 77:24]
  SRAM array ( // @[ICache.scala 50:21]
    .clock(array_clock),
    .io_en(array_io_en),
    .io_addr(array_io_addr),
    .io_wdata(array_io_wdata),
    .io_wen(array_io_wen),
    .io_rdata(array_io_rdata)
  );
  assign auto_out_a_valid = state == 3'h1; // @[ICache.scala 150:24]
  assign auto_out_a_bits_source = source; // @[Edges.scala 447:17 451:15]
  assign auto_out_a_bits_address = {req_r_addr[31:5],5'h0}; // @[Cat.scala 33:92]
  assign auto_out_d_ready = state == 3'h2; // @[ICache.scala 152:24]
  assign io_cache_req_ready = (state == 3'h0 & array_hit | state == 3'h3 | state == 3'h4) & io_cache_resp_ready; // @[ICache.scala 143:92]
  assign io_cache_resp_valid = _s2_ready_T_1 | _s2_ready_T_2; // @[ICache.scala 156:55]
  assign io_cache_resp_bits_rdata = _s2_ready_T_2 ? refill_data : _GEN_1042; // @[ICache.scala 158:25]
  assign array_clock = clock;
  assign array_io_en = fire | _array_io_en_T; // @[ICache.scala 59:26]
  assign array_io_addr = _array_io_en_T ? req_r_addr[14:5] : _GEN_1025; // @[ICache.scala 124:19 125:33]
  assign array_io_wdata = _array_io_en_T ? _array_io_wdata_T_1 : 273'h0; // @[ICache.scala 124:19 126:33 61:18]
  assign array_io_wen = tl_d_ready & auto_out_d_valid; // @[Decoupled.scala 51:35]
  always @(posedge clock) begin
    if (reset) begin // @[ICache.scala 48:22]
      req_r_addr <= 39'h0; // @[ICache.scala 48:22]
    end else if (fire) begin // @[ICache.scala 71:14]
      req_r_addr <= io_cache_req_bits_addr; // @[ICache.scala 73:19]
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_0 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_0 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_0 <= _GEN_1044;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_1 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_1 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_1 <= _GEN_1045;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_2 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_2 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_2 <= _GEN_1046;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_3 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_3 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_3 <= _GEN_1047;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_4 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_4 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_4 <= _GEN_1048;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_5 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_5 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_5 <= _GEN_1049;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_6 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_6 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_6 <= _GEN_1050;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_7 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_7 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_7 <= _GEN_1051;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_8 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_8 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_8 <= _GEN_1052;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_9 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_9 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_9 <= _GEN_1053;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_10 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_10 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_10 <= _GEN_1054;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_11 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_11 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_11 <= _GEN_1055;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_12 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_12 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_12 <= _GEN_1056;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_13 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_13 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_13 <= _GEN_1057;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_14 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_14 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_14 <= _GEN_1058;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_15 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_15 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_15 <= _GEN_1059;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_16 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_16 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_16 <= _GEN_1060;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_17 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_17 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_17 <= _GEN_1061;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_18 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_18 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_18 <= _GEN_1062;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_19 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_19 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_19 <= _GEN_1063;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_20 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_20 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_20 <= _GEN_1064;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_21 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_21 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_21 <= _GEN_1065;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_22 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_22 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_22 <= _GEN_1066;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_23 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_23 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_23 <= _GEN_1067;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_24 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_24 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_24 <= _GEN_1068;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_25 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_25 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_25 <= _GEN_1069;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_26 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_26 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_26 <= _GEN_1070;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_27 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_27 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_27 <= _GEN_1071;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_28 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_28 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_28 <= _GEN_1072;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_29 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_29 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_29 <= _GEN_1073;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_30 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_30 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_30 <= _GEN_1074;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_31 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_31 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_31 <= _GEN_1075;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_32 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_32 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_32 <= _GEN_1076;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_33 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_33 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_33 <= _GEN_1077;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_34 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_34 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_34 <= _GEN_1078;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_35 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_35 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_35 <= _GEN_1079;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_36 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_36 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_36 <= _GEN_1080;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_37 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_37 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_37 <= _GEN_1081;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_38 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_38 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_38 <= _GEN_1082;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_39 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_39 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_39 <= _GEN_1083;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_40 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_40 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_40 <= _GEN_1084;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_41 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_41 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_41 <= _GEN_1085;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_42 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_42 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_42 <= _GEN_1086;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_43 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_43 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_43 <= _GEN_1087;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_44 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_44 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_44 <= _GEN_1088;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_45 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_45 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_45 <= _GEN_1089;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_46 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_46 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_46 <= _GEN_1090;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_47 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_47 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_47 <= _GEN_1091;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_48 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_48 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_48 <= _GEN_1092;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_49 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_49 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_49 <= _GEN_1093;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_50 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_50 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_50 <= _GEN_1094;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_51 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_51 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_51 <= _GEN_1095;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_52 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_52 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_52 <= _GEN_1096;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_53 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_53 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_53 <= _GEN_1097;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_54 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_54 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_54 <= _GEN_1098;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_55 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_55 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_55 <= _GEN_1099;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_56 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_56 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_56 <= _GEN_1100;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_57 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_57 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_57 <= _GEN_1101;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_58 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_58 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_58 <= _GEN_1102;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_59 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_59 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_59 <= _GEN_1103;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_60 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_60 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_60 <= _GEN_1104;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_61 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_61 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_61 <= _GEN_1105;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_62 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_62 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_62 <= _GEN_1106;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_63 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_63 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_63 <= _GEN_1107;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_64 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_64 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_64 <= _GEN_1108;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_65 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_65 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_65 <= _GEN_1109;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_66 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_66 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_66 <= _GEN_1110;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_67 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_67 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_67 <= _GEN_1111;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_68 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_68 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_68 <= _GEN_1112;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_69 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_69 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_69 <= _GEN_1113;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_70 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_70 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_70 <= _GEN_1114;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_71 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_71 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_71 <= _GEN_1115;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_72 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_72 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_72 <= _GEN_1116;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_73 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_73 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_73 <= _GEN_1117;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_74 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_74 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_74 <= _GEN_1118;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_75 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_75 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_75 <= _GEN_1119;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_76 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_76 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_76 <= _GEN_1120;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_77 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_77 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_77 <= _GEN_1121;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_78 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_78 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_78 <= _GEN_1122;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_79 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_79 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_79 <= _GEN_1123;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_80 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_80 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_80 <= _GEN_1124;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_81 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_81 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_81 <= _GEN_1125;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_82 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_82 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_82 <= _GEN_1126;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_83 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_83 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_83 <= _GEN_1127;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_84 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_84 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_84 <= _GEN_1128;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_85 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_85 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_85 <= _GEN_1129;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_86 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_86 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_86 <= _GEN_1130;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_87 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_87 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_87 <= _GEN_1131;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_88 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_88 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_88 <= _GEN_1132;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_89 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_89 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_89 <= _GEN_1133;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_90 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_90 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_90 <= _GEN_1134;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_91 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_91 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_91 <= _GEN_1135;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_92 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_92 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_92 <= _GEN_1136;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_93 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_93 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_93 <= _GEN_1137;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_94 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_94 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_94 <= _GEN_1138;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_95 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_95 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_95 <= _GEN_1139;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_96 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_96 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_96 <= _GEN_1140;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_97 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_97 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_97 <= _GEN_1141;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_98 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_98 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_98 <= _GEN_1142;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_99 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_99 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_99 <= _GEN_1143;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_100 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_100 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_100 <= _GEN_1144;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_101 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_101 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_101 <= _GEN_1145;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_102 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_102 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_102 <= _GEN_1146;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_103 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_103 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_103 <= _GEN_1147;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_104 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_104 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_104 <= _GEN_1148;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_105 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_105 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_105 <= _GEN_1149;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_106 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_106 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_106 <= _GEN_1150;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_107 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_107 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_107 <= _GEN_1151;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_108 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_108 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_108 <= _GEN_1152;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_109 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_109 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_109 <= _GEN_1153;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_110 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_110 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_110 <= _GEN_1154;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_111 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_111 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_111 <= _GEN_1155;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_112 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_112 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_112 <= _GEN_1156;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_113 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_113 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_113 <= _GEN_1157;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_114 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_114 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_114 <= _GEN_1158;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_115 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_115 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_115 <= _GEN_1159;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_116 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_116 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_116 <= _GEN_1160;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_117 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_117 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_117 <= _GEN_1161;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_118 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_118 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_118 <= _GEN_1162;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_119 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_119 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_119 <= _GEN_1163;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_120 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_120 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_120 <= _GEN_1164;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_121 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_121 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_121 <= _GEN_1165;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_122 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_122 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_122 <= _GEN_1166;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_123 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_123 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_123 <= _GEN_1167;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_124 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_124 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_124 <= _GEN_1168;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_125 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_125 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_125 <= _GEN_1169;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_126 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_126 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_126 <= _GEN_1170;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_127 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_127 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_127 <= _GEN_1171;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_128 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_128 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_128 <= _GEN_1172;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_129 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_129 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_129 <= _GEN_1173;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_130 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_130 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_130 <= _GEN_1174;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_131 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_131 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_131 <= _GEN_1175;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_132 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_132 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_132 <= _GEN_1176;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_133 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_133 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_133 <= _GEN_1177;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_134 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_134 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_134 <= _GEN_1178;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_135 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_135 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_135 <= _GEN_1179;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_136 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_136 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_136 <= _GEN_1180;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_137 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_137 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_137 <= _GEN_1181;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_138 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_138 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_138 <= _GEN_1182;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_139 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_139 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_139 <= _GEN_1183;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_140 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_140 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_140 <= _GEN_1184;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_141 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_141 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_141 <= _GEN_1185;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_142 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_142 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_142 <= _GEN_1186;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_143 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_143 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_143 <= _GEN_1187;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_144 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_144 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_144 <= _GEN_1188;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_145 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_145 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_145 <= _GEN_1189;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_146 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_146 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_146 <= _GEN_1190;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_147 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_147 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_147 <= _GEN_1191;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_148 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_148 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_148 <= _GEN_1192;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_149 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_149 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_149 <= _GEN_1193;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_150 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_150 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_150 <= _GEN_1194;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_151 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_151 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_151 <= _GEN_1195;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_152 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_152 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_152 <= _GEN_1196;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_153 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_153 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_153 <= _GEN_1197;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_154 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_154 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_154 <= _GEN_1198;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_155 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_155 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_155 <= _GEN_1199;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_156 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_156 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_156 <= _GEN_1200;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_157 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_157 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_157 <= _GEN_1201;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_158 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_158 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_158 <= _GEN_1202;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_159 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_159 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_159 <= _GEN_1203;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_160 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_160 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_160 <= _GEN_1204;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_161 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_161 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_161 <= _GEN_1205;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_162 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_162 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_162 <= _GEN_1206;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_163 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_163 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_163 <= _GEN_1207;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_164 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_164 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_164 <= _GEN_1208;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_165 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_165 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_165 <= _GEN_1209;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_166 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_166 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_166 <= _GEN_1210;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_167 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_167 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_167 <= _GEN_1211;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_168 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_168 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_168 <= _GEN_1212;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_169 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_169 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_169 <= _GEN_1213;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_170 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_170 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_170 <= _GEN_1214;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_171 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_171 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_171 <= _GEN_1215;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_172 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_172 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_172 <= _GEN_1216;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_173 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_173 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_173 <= _GEN_1217;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_174 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_174 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_174 <= _GEN_1218;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_175 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_175 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_175 <= _GEN_1219;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_176 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_176 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_176 <= _GEN_1220;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_177 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_177 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_177 <= _GEN_1221;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_178 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_178 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_178 <= _GEN_1222;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_179 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_179 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_179 <= _GEN_1223;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_180 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_180 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_180 <= _GEN_1224;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_181 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_181 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_181 <= _GEN_1225;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_182 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_182 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_182 <= _GEN_1226;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_183 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_183 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_183 <= _GEN_1227;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_184 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_184 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_184 <= _GEN_1228;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_185 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_185 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_185 <= _GEN_1229;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_186 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_186 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_186 <= _GEN_1230;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_187 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_187 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_187 <= _GEN_1231;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_188 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_188 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_188 <= _GEN_1232;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_189 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_189 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_189 <= _GEN_1233;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_190 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_190 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_190 <= _GEN_1234;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_191 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_191 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_191 <= _GEN_1235;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_192 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_192 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_192 <= _GEN_1236;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_193 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_193 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_193 <= _GEN_1237;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_194 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_194 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_194 <= _GEN_1238;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_195 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_195 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_195 <= _GEN_1239;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_196 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_196 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_196 <= _GEN_1240;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_197 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_197 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_197 <= _GEN_1241;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_198 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_198 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_198 <= _GEN_1242;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_199 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_199 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_199 <= _GEN_1243;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_200 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_200 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_200 <= _GEN_1244;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_201 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_201 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_201 <= _GEN_1245;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_202 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_202 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_202 <= _GEN_1246;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_203 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_203 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_203 <= _GEN_1247;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_204 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_204 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_204 <= _GEN_1248;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_205 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_205 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_205 <= _GEN_1249;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_206 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_206 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_206 <= _GEN_1250;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_207 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_207 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_207 <= _GEN_1251;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_208 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_208 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_208 <= _GEN_1252;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_209 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_209 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_209 <= _GEN_1253;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_210 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_210 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_210 <= _GEN_1254;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_211 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_211 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_211 <= _GEN_1255;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_212 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_212 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_212 <= _GEN_1256;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_213 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_213 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_213 <= _GEN_1257;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_214 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_214 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_214 <= _GEN_1258;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_215 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_215 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_215 <= _GEN_1259;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_216 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_216 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_216 <= _GEN_1260;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_217 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_217 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_217 <= _GEN_1261;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_218 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_218 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_218 <= _GEN_1262;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_219 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_219 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_219 <= _GEN_1263;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_220 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_220 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_220 <= _GEN_1264;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_221 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_221 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_221 <= _GEN_1265;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_222 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_222 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_222 <= _GEN_1266;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_223 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_223 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_223 <= _GEN_1267;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_224 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_224 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_224 <= _GEN_1268;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_225 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_225 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_225 <= _GEN_1269;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_226 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_226 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_226 <= _GEN_1270;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_227 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_227 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_227 <= _GEN_1271;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_228 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_228 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_228 <= _GEN_1272;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_229 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_229 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_229 <= _GEN_1273;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_230 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_230 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_230 <= _GEN_1274;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_231 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_231 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_231 <= _GEN_1275;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_232 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_232 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_232 <= _GEN_1276;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_233 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_233 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_233 <= _GEN_1277;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_234 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_234 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_234 <= _GEN_1278;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_235 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_235 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_235 <= _GEN_1279;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_236 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_236 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_236 <= _GEN_1280;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_237 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_237 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_237 <= _GEN_1281;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_238 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_238 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_238 <= _GEN_1282;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_239 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_239 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_239 <= _GEN_1283;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_240 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_240 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_240 <= _GEN_1284;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_241 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_241 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_241 <= _GEN_1285;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_242 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_242 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_242 <= _GEN_1286;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_243 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_243 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_243 <= _GEN_1287;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_244 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_244 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_244 <= _GEN_1288;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_245 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_245 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_245 <= _GEN_1289;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_246 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_246 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_246 <= _GEN_1290;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_247 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_247 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_247 <= _GEN_1291;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_248 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_248 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_248 <= _GEN_1292;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_249 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_249 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_249 <= _GEN_1293;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_250 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_250 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_250 <= _GEN_1294;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_251 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_251 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_251 <= _GEN_1295;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_252 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_252 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_252 <= _GEN_1296;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_253 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_253 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_253 <= _GEN_1297;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_254 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_254 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_254 <= _GEN_1298;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_255 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_255 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_255 <= _GEN_1299;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_256 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_256 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_256 <= _GEN_1300;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_257 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_257 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_257 <= _GEN_1301;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_258 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_258 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_258 <= _GEN_1302;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_259 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_259 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_259 <= _GEN_1303;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_260 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_260 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_260 <= _GEN_1304;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_261 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_261 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_261 <= _GEN_1305;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_262 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_262 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_262 <= _GEN_1306;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_263 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_263 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_263 <= _GEN_1307;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_264 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_264 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_264 <= _GEN_1308;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_265 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_265 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_265 <= _GEN_1309;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_266 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_266 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_266 <= _GEN_1310;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_267 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_267 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_267 <= _GEN_1311;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_268 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_268 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_268 <= _GEN_1312;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_269 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_269 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_269 <= _GEN_1313;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_270 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_270 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_270 <= _GEN_1314;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_271 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_271 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_271 <= _GEN_1315;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_272 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_272 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_272 <= _GEN_1316;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_273 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_273 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_273 <= _GEN_1317;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_274 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_274 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_274 <= _GEN_1318;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_275 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_275 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_275 <= _GEN_1319;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_276 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_276 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_276 <= _GEN_1320;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_277 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_277 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_277 <= _GEN_1321;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_278 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_278 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_278 <= _GEN_1322;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_279 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_279 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_279 <= _GEN_1323;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_280 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_280 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_280 <= _GEN_1324;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_281 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_281 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_281 <= _GEN_1325;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_282 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_282 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_282 <= _GEN_1326;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_283 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_283 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_283 <= _GEN_1327;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_284 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_284 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_284 <= _GEN_1328;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_285 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_285 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_285 <= _GEN_1329;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_286 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_286 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_286 <= _GEN_1330;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_287 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_287 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_287 <= _GEN_1331;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_288 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_288 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_288 <= _GEN_1332;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_289 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_289 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_289 <= _GEN_1333;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_290 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_290 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_290 <= _GEN_1334;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_291 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_291 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_291 <= _GEN_1335;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_292 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_292 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_292 <= _GEN_1336;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_293 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_293 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_293 <= _GEN_1337;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_294 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_294 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_294 <= _GEN_1338;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_295 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_295 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_295 <= _GEN_1339;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_296 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_296 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_296 <= _GEN_1340;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_297 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_297 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_297 <= _GEN_1341;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_298 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_298 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_298 <= _GEN_1342;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_299 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_299 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_299 <= _GEN_1343;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_300 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_300 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_300 <= _GEN_1344;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_301 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_301 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_301 <= _GEN_1345;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_302 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_302 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_302 <= _GEN_1346;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_303 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_303 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_303 <= _GEN_1347;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_304 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_304 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_304 <= _GEN_1348;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_305 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_305 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_305 <= _GEN_1349;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_306 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_306 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_306 <= _GEN_1350;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_307 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_307 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_307 <= _GEN_1351;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_308 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_308 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_308 <= _GEN_1352;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_309 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_309 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_309 <= _GEN_1353;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_310 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_310 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_310 <= _GEN_1354;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_311 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_311 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_311 <= _GEN_1355;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_312 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_312 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_312 <= _GEN_1356;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_313 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_313 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_313 <= _GEN_1357;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_314 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_314 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_314 <= _GEN_1358;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_315 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_315 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_315 <= _GEN_1359;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_316 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_316 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_316 <= _GEN_1360;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_317 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_317 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_317 <= _GEN_1361;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_318 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_318 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_318 <= _GEN_1362;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_319 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_319 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_319 <= _GEN_1363;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_320 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_320 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_320 <= _GEN_1364;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_321 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_321 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_321 <= _GEN_1365;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_322 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_322 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_322 <= _GEN_1366;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_323 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_323 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_323 <= _GEN_1367;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_324 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_324 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_324 <= _GEN_1368;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_325 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_325 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_325 <= _GEN_1369;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_326 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_326 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_326 <= _GEN_1370;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_327 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_327 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_327 <= _GEN_1371;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_328 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_328 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_328 <= _GEN_1372;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_329 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_329 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_329 <= _GEN_1373;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_330 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_330 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_330 <= _GEN_1374;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_331 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_331 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_331 <= _GEN_1375;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_332 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_332 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_332 <= _GEN_1376;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_333 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_333 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_333 <= _GEN_1377;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_334 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_334 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_334 <= _GEN_1378;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_335 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_335 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_335 <= _GEN_1379;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_336 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_336 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_336 <= _GEN_1380;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_337 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_337 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_337 <= _GEN_1381;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_338 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_338 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_338 <= _GEN_1382;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_339 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_339 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_339 <= _GEN_1383;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_340 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_340 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_340 <= _GEN_1384;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_341 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_341 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_341 <= _GEN_1385;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_342 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_342 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_342 <= _GEN_1386;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_343 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_343 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_343 <= _GEN_1387;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_344 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_344 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_344 <= _GEN_1388;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_345 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_345 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_345 <= _GEN_1389;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_346 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_346 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_346 <= _GEN_1390;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_347 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_347 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_347 <= _GEN_1391;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_348 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_348 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_348 <= _GEN_1392;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_349 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_349 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_349 <= _GEN_1393;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_350 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_350 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_350 <= _GEN_1394;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_351 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_351 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_351 <= _GEN_1395;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_352 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_352 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_352 <= _GEN_1396;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_353 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_353 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_353 <= _GEN_1397;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_354 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_354 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_354 <= _GEN_1398;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_355 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_355 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_355 <= _GEN_1399;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_356 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_356 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_356 <= _GEN_1400;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_357 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_357 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_357 <= _GEN_1401;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_358 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_358 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_358 <= _GEN_1402;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_359 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_359 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_359 <= _GEN_1403;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_360 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_360 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_360 <= _GEN_1404;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_361 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_361 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_361 <= _GEN_1405;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_362 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_362 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_362 <= _GEN_1406;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_363 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_363 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_363 <= _GEN_1407;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_364 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_364 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_364 <= _GEN_1408;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_365 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_365 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_365 <= _GEN_1409;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_366 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_366 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_366 <= _GEN_1410;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_367 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_367 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_367 <= _GEN_1411;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_368 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_368 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_368 <= _GEN_1412;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_369 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_369 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_369 <= _GEN_1413;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_370 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_370 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_370 <= _GEN_1414;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_371 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_371 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_371 <= _GEN_1415;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_372 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_372 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_372 <= _GEN_1416;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_373 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_373 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_373 <= _GEN_1417;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_374 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_374 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_374 <= _GEN_1418;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_375 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_375 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_375 <= _GEN_1419;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_376 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_376 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_376 <= _GEN_1420;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_377 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_377 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_377 <= _GEN_1421;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_378 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_378 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_378 <= _GEN_1422;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_379 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_379 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_379 <= _GEN_1423;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_380 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_380 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_380 <= _GEN_1424;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_381 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_381 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_381 <= _GEN_1425;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_382 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_382 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_382 <= _GEN_1426;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_383 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_383 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_383 <= _GEN_1427;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_384 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_384 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_384 <= _GEN_1428;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_385 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_385 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_385 <= _GEN_1429;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_386 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_386 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_386 <= _GEN_1430;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_387 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_387 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_387 <= _GEN_1431;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_388 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_388 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_388 <= _GEN_1432;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_389 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_389 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_389 <= _GEN_1433;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_390 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_390 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_390 <= _GEN_1434;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_391 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_391 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_391 <= _GEN_1435;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_392 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_392 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_392 <= _GEN_1436;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_393 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_393 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_393 <= _GEN_1437;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_394 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_394 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_394 <= _GEN_1438;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_395 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_395 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_395 <= _GEN_1439;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_396 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_396 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_396 <= _GEN_1440;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_397 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_397 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_397 <= _GEN_1441;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_398 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_398 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_398 <= _GEN_1442;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_399 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_399 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_399 <= _GEN_1443;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_400 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_400 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_400 <= _GEN_1444;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_401 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_401 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_401 <= _GEN_1445;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_402 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_402 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_402 <= _GEN_1446;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_403 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_403 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_403 <= _GEN_1447;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_404 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_404 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_404 <= _GEN_1448;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_405 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_405 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_405 <= _GEN_1449;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_406 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_406 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_406 <= _GEN_1450;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_407 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_407 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_407 <= _GEN_1451;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_408 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_408 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_408 <= _GEN_1452;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_409 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_409 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_409 <= _GEN_1453;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_410 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_410 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_410 <= _GEN_1454;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_411 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_411 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_411 <= _GEN_1455;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_412 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_412 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_412 <= _GEN_1456;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_413 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_413 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_413 <= _GEN_1457;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_414 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_414 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_414 <= _GEN_1458;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_415 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_415 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_415 <= _GEN_1459;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_416 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_416 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_416 <= _GEN_1460;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_417 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_417 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_417 <= _GEN_1461;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_418 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_418 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_418 <= _GEN_1462;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_419 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_419 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_419 <= _GEN_1463;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_420 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_420 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_420 <= _GEN_1464;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_421 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_421 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_421 <= _GEN_1465;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_422 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_422 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_422 <= _GEN_1466;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_423 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_423 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_423 <= _GEN_1467;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_424 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_424 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_424 <= _GEN_1468;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_425 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_425 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_425 <= _GEN_1469;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_426 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_426 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_426 <= _GEN_1470;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_427 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_427 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_427 <= _GEN_1471;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_428 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_428 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_428 <= _GEN_1472;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_429 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_429 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_429 <= _GEN_1473;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_430 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_430 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_430 <= _GEN_1474;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_431 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_431 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_431 <= _GEN_1475;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_432 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_432 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_432 <= _GEN_1476;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_433 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_433 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_433 <= _GEN_1477;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_434 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_434 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_434 <= _GEN_1478;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_435 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_435 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_435 <= _GEN_1479;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_436 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_436 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_436 <= _GEN_1480;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_437 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_437 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_437 <= _GEN_1481;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_438 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_438 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_438 <= _GEN_1482;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_439 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_439 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_439 <= _GEN_1483;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_440 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_440 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_440 <= _GEN_1484;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_441 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_441 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_441 <= _GEN_1485;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_442 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_442 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_442 <= _GEN_1486;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_443 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_443 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_443 <= _GEN_1487;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_444 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_444 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_444 <= _GEN_1488;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_445 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_445 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_445 <= _GEN_1489;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_446 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_446 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_446 <= _GEN_1490;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_447 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_447 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_447 <= _GEN_1491;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_448 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_448 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_448 <= _GEN_1492;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_449 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_449 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_449 <= _GEN_1493;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_450 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_450 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_450 <= _GEN_1494;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_451 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_451 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_451 <= _GEN_1495;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_452 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_452 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_452 <= _GEN_1496;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_453 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_453 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_453 <= _GEN_1497;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_454 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_454 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_454 <= _GEN_1498;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_455 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_455 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_455 <= _GEN_1499;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_456 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_456 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_456 <= _GEN_1500;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_457 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_457 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_457 <= _GEN_1501;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_458 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_458 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_458 <= _GEN_1502;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_459 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_459 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_459 <= _GEN_1503;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_460 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_460 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_460 <= _GEN_1504;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_461 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_461 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_461 <= _GEN_1505;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_462 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_462 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_462 <= _GEN_1506;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_463 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_463 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_463 <= _GEN_1507;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_464 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_464 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_464 <= _GEN_1508;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_465 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_465 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_465 <= _GEN_1509;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_466 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_466 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_466 <= _GEN_1510;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_467 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_467 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_467 <= _GEN_1511;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_468 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_468 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_468 <= _GEN_1512;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_469 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_469 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_469 <= _GEN_1513;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_470 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_470 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_470 <= _GEN_1514;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_471 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_471 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_471 <= _GEN_1515;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_472 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_472 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_472 <= _GEN_1516;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_473 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_473 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_473 <= _GEN_1517;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_474 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_474 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_474 <= _GEN_1518;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_475 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_475 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_475 <= _GEN_1519;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_476 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_476 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_476 <= _GEN_1520;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_477 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_477 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_477 <= _GEN_1521;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_478 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_478 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_478 <= _GEN_1522;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_479 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_479 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_479 <= _GEN_1523;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_480 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_480 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_480 <= _GEN_1524;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_481 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_481 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_481 <= _GEN_1525;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_482 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_482 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_482 <= _GEN_1526;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_483 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_483 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_483 <= _GEN_1527;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_484 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_484 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_484 <= _GEN_1528;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_485 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_485 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_485 <= _GEN_1529;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_486 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_486 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_486 <= _GEN_1530;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_487 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_487 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_487 <= _GEN_1531;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_488 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_488 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_488 <= _GEN_1532;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_489 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_489 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_489 <= _GEN_1533;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_490 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_490 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_490 <= _GEN_1534;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_491 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_491 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_491 <= _GEN_1535;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_492 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_492 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_492 <= _GEN_1536;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_493 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_493 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_493 <= _GEN_1537;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_494 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_494 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_494 <= _GEN_1538;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_495 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_495 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_495 <= _GEN_1539;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_496 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_496 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_496 <= _GEN_1540;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_497 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_497 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_497 <= _GEN_1541;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_498 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_498 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_498 <= _GEN_1542;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_499 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_499 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_499 <= _GEN_1543;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_500 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_500 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_500 <= _GEN_1544;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_501 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_501 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_501 <= _GEN_1545;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_502 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_502 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_502 <= _GEN_1546;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_503 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_503 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_503 <= _GEN_1547;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_504 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_504 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_504 <= _GEN_1548;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_505 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_505 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_505 <= _GEN_1549;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_506 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_506 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_506 <= _GEN_1550;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_507 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_507 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_507 <= _GEN_1551;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_508 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_508 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_508 <= _GEN_1552;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_509 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_509 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_509 <= _GEN_1553;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_510 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_510 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_510 <= _GEN_1554;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_511 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_511 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_511 <= _GEN_1555;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_512 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_512 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_512 <= _GEN_1556;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_513 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_513 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_513 <= _GEN_1557;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_514 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_514 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_514 <= _GEN_1558;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_515 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_515 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_515 <= _GEN_1559;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_516 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_516 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_516 <= _GEN_1560;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_517 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_517 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_517 <= _GEN_1561;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_518 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_518 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_518 <= _GEN_1562;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_519 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_519 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_519 <= _GEN_1563;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_520 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_520 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_520 <= _GEN_1564;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_521 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_521 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_521 <= _GEN_1565;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_522 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_522 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_522 <= _GEN_1566;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_523 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_523 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_523 <= _GEN_1567;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_524 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_524 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_524 <= _GEN_1568;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_525 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_525 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_525 <= _GEN_1569;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_526 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_526 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_526 <= _GEN_1570;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_527 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_527 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_527 <= _GEN_1571;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_528 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_528 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_528 <= _GEN_1572;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_529 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_529 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_529 <= _GEN_1573;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_530 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_530 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_530 <= _GEN_1574;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_531 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_531 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_531 <= _GEN_1575;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_532 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_532 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_532 <= _GEN_1576;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_533 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_533 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_533 <= _GEN_1577;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_534 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_534 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_534 <= _GEN_1578;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_535 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_535 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_535 <= _GEN_1579;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_536 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_536 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_536 <= _GEN_1580;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_537 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_537 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_537 <= _GEN_1581;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_538 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_538 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_538 <= _GEN_1582;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_539 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_539 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_539 <= _GEN_1583;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_540 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_540 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_540 <= _GEN_1584;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_541 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_541 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_541 <= _GEN_1585;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_542 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_542 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_542 <= _GEN_1586;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_543 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_543 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_543 <= _GEN_1587;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_544 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_544 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_544 <= _GEN_1588;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_545 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_545 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_545 <= _GEN_1589;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_546 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_546 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_546 <= _GEN_1590;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_547 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_547 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_547 <= _GEN_1591;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_548 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_548 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_548 <= _GEN_1592;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_549 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_549 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_549 <= _GEN_1593;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_550 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_550 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_550 <= _GEN_1594;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_551 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_551 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_551 <= _GEN_1595;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_552 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_552 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_552 <= _GEN_1596;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_553 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_553 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_553 <= _GEN_1597;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_554 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_554 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_554 <= _GEN_1598;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_555 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_555 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_555 <= _GEN_1599;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_556 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_556 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_556 <= _GEN_1600;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_557 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_557 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_557 <= _GEN_1601;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_558 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_558 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_558 <= _GEN_1602;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_559 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_559 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_559 <= _GEN_1603;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_560 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_560 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_560 <= _GEN_1604;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_561 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_561 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_561 <= _GEN_1605;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_562 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_562 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_562 <= _GEN_1606;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_563 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_563 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_563 <= _GEN_1607;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_564 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_564 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_564 <= _GEN_1608;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_565 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_565 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_565 <= _GEN_1609;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_566 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_566 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_566 <= _GEN_1610;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_567 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_567 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_567 <= _GEN_1611;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_568 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_568 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_568 <= _GEN_1612;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_569 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_569 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_569 <= _GEN_1613;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_570 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_570 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_570 <= _GEN_1614;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_571 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_571 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_571 <= _GEN_1615;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_572 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_572 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_572 <= _GEN_1616;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_573 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_573 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_573 <= _GEN_1617;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_574 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_574 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_574 <= _GEN_1618;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_575 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_575 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_575 <= _GEN_1619;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_576 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_576 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_576 <= _GEN_1620;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_577 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_577 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_577 <= _GEN_1621;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_578 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_578 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_578 <= _GEN_1622;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_579 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_579 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_579 <= _GEN_1623;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_580 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_580 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_580 <= _GEN_1624;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_581 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_581 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_581 <= _GEN_1625;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_582 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_582 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_582 <= _GEN_1626;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_583 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_583 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_583 <= _GEN_1627;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_584 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_584 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_584 <= _GEN_1628;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_585 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_585 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_585 <= _GEN_1629;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_586 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_586 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_586 <= _GEN_1630;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_587 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_587 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_587 <= _GEN_1631;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_588 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_588 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_588 <= _GEN_1632;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_589 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_589 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_589 <= _GEN_1633;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_590 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_590 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_590 <= _GEN_1634;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_591 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_591 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_591 <= _GEN_1635;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_592 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_592 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_592 <= _GEN_1636;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_593 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_593 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_593 <= _GEN_1637;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_594 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_594 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_594 <= _GEN_1638;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_595 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_595 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_595 <= _GEN_1639;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_596 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_596 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_596 <= _GEN_1640;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_597 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_597 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_597 <= _GEN_1641;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_598 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_598 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_598 <= _GEN_1642;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_599 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_599 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_599 <= _GEN_1643;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_600 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_600 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_600 <= _GEN_1644;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_601 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_601 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_601 <= _GEN_1645;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_602 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_602 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_602 <= _GEN_1646;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_603 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_603 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_603 <= _GEN_1647;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_604 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_604 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_604 <= _GEN_1648;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_605 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_605 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_605 <= _GEN_1649;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_606 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_606 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_606 <= _GEN_1650;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_607 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_607 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_607 <= _GEN_1651;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_608 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_608 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_608 <= _GEN_1652;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_609 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_609 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_609 <= _GEN_1653;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_610 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_610 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_610 <= _GEN_1654;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_611 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_611 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_611 <= _GEN_1655;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_612 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_612 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_612 <= _GEN_1656;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_613 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_613 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_613 <= _GEN_1657;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_614 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_614 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_614 <= _GEN_1658;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_615 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_615 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_615 <= _GEN_1659;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_616 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_616 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_616 <= _GEN_1660;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_617 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_617 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_617 <= _GEN_1661;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_618 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_618 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_618 <= _GEN_1662;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_619 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_619 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_619 <= _GEN_1663;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_620 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_620 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_620 <= _GEN_1664;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_621 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_621 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_621 <= _GEN_1665;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_622 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_622 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_622 <= _GEN_1666;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_623 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_623 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_623 <= _GEN_1667;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_624 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_624 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_624 <= _GEN_1668;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_625 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_625 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_625 <= _GEN_1669;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_626 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_626 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_626 <= _GEN_1670;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_627 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_627 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_627 <= _GEN_1671;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_628 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_628 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_628 <= _GEN_1672;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_629 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_629 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_629 <= _GEN_1673;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_630 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_630 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_630 <= _GEN_1674;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_631 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_631 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_631 <= _GEN_1675;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_632 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_632 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_632 <= _GEN_1676;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_633 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_633 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_633 <= _GEN_1677;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_634 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_634 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_634 <= _GEN_1678;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_635 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_635 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_635 <= _GEN_1679;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_636 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_636 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_636 <= _GEN_1680;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_637 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_637 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_637 <= _GEN_1681;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_638 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_638 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_638 <= _GEN_1682;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_639 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_639 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_639 <= _GEN_1683;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_640 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_640 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_640 <= _GEN_1684;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_641 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_641 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_641 <= _GEN_1685;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_642 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_642 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_642 <= _GEN_1686;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_643 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_643 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_643 <= _GEN_1687;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_644 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_644 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_644 <= _GEN_1688;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_645 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_645 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_645 <= _GEN_1689;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_646 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_646 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_646 <= _GEN_1690;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_647 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_647 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_647 <= _GEN_1691;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_648 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_648 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_648 <= _GEN_1692;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_649 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_649 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_649 <= _GEN_1693;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_650 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_650 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_650 <= _GEN_1694;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_651 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_651 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_651 <= _GEN_1695;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_652 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_652 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_652 <= _GEN_1696;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_653 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_653 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_653 <= _GEN_1697;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_654 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_654 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_654 <= _GEN_1698;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_655 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_655 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_655 <= _GEN_1699;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_656 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_656 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_656 <= _GEN_1700;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_657 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_657 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_657 <= _GEN_1701;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_658 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_658 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_658 <= _GEN_1702;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_659 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_659 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_659 <= _GEN_1703;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_660 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_660 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_660 <= _GEN_1704;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_661 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_661 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_661 <= _GEN_1705;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_662 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_662 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_662 <= _GEN_1706;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_663 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_663 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_663 <= _GEN_1707;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_664 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_664 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_664 <= _GEN_1708;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_665 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_665 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_665 <= _GEN_1709;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_666 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_666 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_666 <= _GEN_1710;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_667 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_667 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_667 <= _GEN_1711;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_668 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_668 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_668 <= _GEN_1712;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_669 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_669 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_669 <= _GEN_1713;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_670 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_670 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_670 <= _GEN_1714;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_671 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_671 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_671 <= _GEN_1715;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_672 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_672 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_672 <= _GEN_1716;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_673 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_673 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_673 <= _GEN_1717;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_674 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_674 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_674 <= _GEN_1718;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_675 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_675 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_675 <= _GEN_1719;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_676 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_676 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_676 <= _GEN_1720;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_677 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_677 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_677 <= _GEN_1721;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_678 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_678 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_678 <= _GEN_1722;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_679 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_679 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_679 <= _GEN_1723;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_680 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_680 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_680 <= _GEN_1724;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_681 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_681 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_681 <= _GEN_1725;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_682 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_682 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_682 <= _GEN_1726;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_683 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_683 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_683 <= _GEN_1727;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_684 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_684 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_684 <= _GEN_1728;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_685 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_685 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_685 <= _GEN_1729;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_686 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_686 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_686 <= _GEN_1730;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_687 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_687 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_687 <= _GEN_1731;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_688 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_688 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_688 <= _GEN_1732;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_689 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_689 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_689 <= _GEN_1733;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_690 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_690 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_690 <= _GEN_1734;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_691 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_691 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_691 <= _GEN_1735;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_692 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_692 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_692 <= _GEN_1736;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_693 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_693 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_693 <= _GEN_1737;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_694 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_694 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_694 <= _GEN_1738;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_695 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_695 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_695 <= _GEN_1739;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_696 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_696 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_696 <= _GEN_1740;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_697 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_697 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_697 <= _GEN_1741;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_698 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_698 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_698 <= _GEN_1742;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_699 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_699 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_699 <= _GEN_1743;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_700 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_700 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_700 <= _GEN_1744;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_701 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_701 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_701 <= _GEN_1745;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_702 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_702 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_702 <= _GEN_1746;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_703 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_703 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_703 <= _GEN_1747;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_704 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_704 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_704 <= _GEN_1748;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_705 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_705 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_705 <= _GEN_1749;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_706 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_706 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_706 <= _GEN_1750;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_707 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_707 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_707 <= _GEN_1751;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_708 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_708 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_708 <= _GEN_1752;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_709 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_709 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_709 <= _GEN_1753;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_710 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_710 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_710 <= _GEN_1754;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_711 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_711 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_711 <= _GEN_1755;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_712 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_712 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_712 <= _GEN_1756;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_713 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_713 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_713 <= _GEN_1757;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_714 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_714 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_714 <= _GEN_1758;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_715 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_715 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_715 <= _GEN_1759;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_716 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_716 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_716 <= _GEN_1760;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_717 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_717 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_717 <= _GEN_1761;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_718 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_718 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_718 <= _GEN_1762;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_719 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_719 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_719 <= _GEN_1763;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_720 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_720 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_720 <= _GEN_1764;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_721 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_721 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_721 <= _GEN_1765;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_722 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_722 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_722 <= _GEN_1766;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_723 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_723 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_723 <= _GEN_1767;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_724 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_724 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_724 <= _GEN_1768;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_725 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_725 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_725 <= _GEN_1769;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_726 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_726 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_726 <= _GEN_1770;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_727 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_727 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_727 <= _GEN_1771;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_728 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_728 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_728 <= _GEN_1772;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_729 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_729 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_729 <= _GEN_1773;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_730 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_730 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_730 <= _GEN_1774;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_731 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_731 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_731 <= _GEN_1775;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_732 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_732 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_732 <= _GEN_1776;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_733 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_733 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_733 <= _GEN_1777;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_734 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_734 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_734 <= _GEN_1778;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_735 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_735 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_735 <= _GEN_1779;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_736 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_736 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_736 <= _GEN_1780;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_737 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_737 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_737 <= _GEN_1781;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_738 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_738 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_738 <= _GEN_1782;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_739 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_739 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_739 <= _GEN_1783;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_740 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_740 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_740 <= _GEN_1784;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_741 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_741 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_741 <= _GEN_1785;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_742 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_742 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_742 <= _GEN_1786;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_743 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_743 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_743 <= _GEN_1787;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_744 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_744 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_744 <= _GEN_1788;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_745 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_745 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_745 <= _GEN_1789;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_746 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_746 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_746 <= _GEN_1790;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_747 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_747 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_747 <= _GEN_1791;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_748 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_748 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_748 <= _GEN_1792;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_749 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_749 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_749 <= _GEN_1793;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_750 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_750 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_750 <= _GEN_1794;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_751 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_751 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_751 <= _GEN_1795;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_752 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_752 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_752 <= _GEN_1796;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_753 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_753 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_753 <= _GEN_1797;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_754 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_754 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_754 <= _GEN_1798;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_755 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_755 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_755 <= _GEN_1799;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_756 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_756 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_756 <= _GEN_1800;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_757 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_757 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_757 <= _GEN_1801;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_758 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_758 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_758 <= _GEN_1802;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_759 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_759 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_759 <= _GEN_1803;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_760 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_760 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_760 <= _GEN_1804;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_761 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_761 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_761 <= _GEN_1805;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_762 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_762 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_762 <= _GEN_1806;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_763 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_763 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_763 <= _GEN_1807;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_764 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_764 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_764 <= _GEN_1808;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_765 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_765 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_765 <= _GEN_1809;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_766 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_766 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_766 <= _GEN_1810;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_767 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_767 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_767 <= _GEN_1811;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_768 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_768 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_768 <= _GEN_1812;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_769 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_769 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_769 <= _GEN_1813;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_770 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_770 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_770 <= _GEN_1814;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_771 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_771 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_771 <= _GEN_1815;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_772 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_772 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_772 <= _GEN_1816;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_773 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_773 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_773 <= _GEN_1817;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_774 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_774 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_774 <= _GEN_1818;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_775 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_775 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_775 <= _GEN_1819;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_776 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_776 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_776 <= _GEN_1820;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_777 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_777 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_777 <= _GEN_1821;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_778 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_778 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_778 <= _GEN_1822;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_779 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_779 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_779 <= _GEN_1823;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_780 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_780 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_780 <= _GEN_1824;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_781 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_781 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_781 <= _GEN_1825;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_782 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_782 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_782 <= _GEN_1826;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_783 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_783 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_783 <= _GEN_1827;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_784 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_784 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_784 <= _GEN_1828;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_785 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_785 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_785 <= _GEN_1829;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_786 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_786 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_786 <= _GEN_1830;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_787 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_787 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_787 <= _GEN_1831;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_788 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_788 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_788 <= _GEN_1832;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_789 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_789 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_789 <= _GEN_1833;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_790 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_790 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_790 <= _GEN_1834;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_791 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_791 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_791 <= _GEN_1835;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_792 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_792 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_792 <= _GEN_1836;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_793 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_793 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_793 <= _GEN_1837;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_794 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_794 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_794 <= _GEN_1838;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_795 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_795 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_795 <= _GEN_1839;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_796 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_796 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_796 <= _GEN_1840;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_797 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_797 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_797 <= _GEN_1841;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_798 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_798 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_798 <= _GEN_1842;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_799 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_799 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_799 <= _GEN_1843;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_800 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_800 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_800 <= _GEN_1844;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_801 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_801 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_801 <= _GEN_1845;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_802 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_802 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_802 <= _GEN_1846;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_803 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_803 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_803 <= _GEN_1847;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_804 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_804 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_804 <= _GEN_1848;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_805 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_805 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_805 <= _GEN_1849;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_806 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_806 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_806 <= _GEN_1850;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_807 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_807 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_807 <= _GEN_1851;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_808 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_808 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_808 <= _GEN_1852;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_809 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_809 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_809 <= _GEN_1853;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_810 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_810 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_810 <= _GEN_1854;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_811 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_811 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_811 <= _GEN_1855;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_812 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_812 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_812 <= _GEN_1856;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_813 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_813 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_813 <= _GEN_1857;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_814 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_814 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_814 <= _GEN_1858;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_815 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_815 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_815 <= _GEN_1859;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_816 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_816 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_816 <= _GEN_1860;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_817 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_817 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_817 <= _GEN_1861;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_818 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_818 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_818 <= _GEN_1862;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_819 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_819 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_819 <= _GEN_1863;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_820 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_820 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_820 <= _GEN_1864;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_821 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_821 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_821 <= _GEN_1865;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_822 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_822 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_822 <= _GEN_1866;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_823 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_823 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_823 <= _GEN_1867;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_824 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_824 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_824 <= _GEN_1868;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_825 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_825 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_825 <= _GEN_1869;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_826 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_826 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_826 <= _GEN_1870;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_827 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_827 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_827 <= _GEN_1871;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_828 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_828 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_828 <= _GEN_1872;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_829 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_829 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_829 <= _GEN_1873;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_830 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_830 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_830 <= _GEN_1874;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_831 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_831 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_831 <= _GEN_1875;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_832 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_832 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_832 <= _GEN_1876;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_833 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_833 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_833 <= _GEN_1877;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_834 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_834 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_834 <= _GEN_1878;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_835 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_835 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_835 <= _GEN_1879;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_836 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_836 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_836 <= _GEN_1880;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_837 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_837 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_837 <= _GEN_1881;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_838 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_838 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_838 <= _GEN_1882;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_839 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_839 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_839 <= _GEN_1883;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_840 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_840 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_840 <= _GEN_1884;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_841 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_841 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_841 <= _GEN_1885;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_842 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_842 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_842 <= _GEN_1886;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_843 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_843 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_843 <= _GEN_1887;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_844 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_844 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_844 <= _GEN_1888;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_845 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_845 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_845 <= _GEN_1889;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_846 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_846 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_846 <= _GEN_1890;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_847 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_847 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_847 <= _GEN_1891;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_848 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_848 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_848 <= _GEN_1892;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_849 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_849 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_849 <= _GEN_1893;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_850 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_850 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_850 <= _GEN_1894;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_851 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_851 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_851 <= _GEN_1895;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_852 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_852 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_852 <= _GEN_1896;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_853 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_853 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_853 <= _GEN_1897;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_854 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_854 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_854 <= _GEN_1898;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_855 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_855 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_855 <= _GEN_1899;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_856 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_856 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_856 <= _GEN_1900;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_857 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_857 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_857 <= _GEN_1901;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_858 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_858 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_858 <= _GEN_1902;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_859 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_859 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_859 <= _GEN_1903;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_860 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_860 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_860 <= _GEN_1904;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_861 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_861 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_861 <= _GEN_1905;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_862 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_862 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_862 <= _GEN_1906;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_863 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_863 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_863 <= _GEN_1907;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_864 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_864 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_864 <= _GEN_1908;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_865 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_865 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_865 <= _GEN_1909;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_866 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_866 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_866 <= _GEN_1910;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_867 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_867 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_867 <= _GEN_1911;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_868 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_868 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_868 <= _GEN_1912;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_869 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_869 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_869 <= _GEN_1913;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_870 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_870 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_870 <= _GEN_1914;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_871 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_871 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_871 <= _GEN_1915;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_872 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_872 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_872 <= _GEN_1916;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_873 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_873 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_873 <= _GEN_1917;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_874 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_874 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_874 <= _GEN_1918;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_875 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_875 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_875 <= _GEN_1919;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_876 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_876 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_876 <= _GEN_1920;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_877 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_877 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_877 <= _GEN_1921;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_878 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_878 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_878 <= _GEN_1922;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_879 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_879 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_879 <= _GEN_1923;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_880 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_880 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_880 <= _GEN_1924;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_881 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_881 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_881 <= _GEN_1925;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_882 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_882 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_882 <= _GEN_1926;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_883 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_883 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_883 <= _GEN_1927;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_884 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_884 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_884 <= _GEN_1928;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_885 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_885 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_885 <= _GEN_1929;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_886 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_886 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_886 <= _GEN_1930;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_887 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_887 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_887 <= _GEN_1931;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_888 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_888 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_888 <= _GEN_1932;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_889 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_889 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_889 <= _GEN_1933;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_890 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_890 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_890 <= _GEN_1934;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_891 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_891 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_891 <= _GEN_1935;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_892 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_892 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_892 <= _GEN_1936;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_893 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_893 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_893 <= _GEN_1937;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_894 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_894 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_894 <= _GEN_1938;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_895 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_895 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_895 <= _GEN_1939;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_896 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_896 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_896 <= _GEN_1940;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_897 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_897 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_897 <= _GEN_1941;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_898 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_898 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_898 <= _GEN_1942;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_899 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_899 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_899 <= _GEN_1943;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_900 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_900 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_900 <= _GEN_1944;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_901 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_901 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_901 <= _GEN_1945;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_902 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_902 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_902 <= _GEN_1946;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_903 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_903 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_903 <= _GEN_1947;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_904 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_904 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_904 <= _GEN_1948;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_905 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_905 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_905 <= _GEN_1949;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_906 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_906 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_906 <= _GEN_1950;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_907 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_907 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_907 <= _GEN_1951;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_908 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_908 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_908 <= _GEN_1952;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_909 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_909 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_909 <= _GEN_1953;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_910 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_910 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_910 <= _GEN_1954;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_911 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_911 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_911 <= _GEN_1955;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_912 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_912 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_912 <= _GEN_1956;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_913 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_913 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_913 <= _GEN_1957;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_914 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_914 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_914 <= _GEN_1958;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_915 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_915 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_915 <= _GEN_1959;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_916 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_916 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_916 <= _GEN_1960;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_917 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_917 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_917 <= _GEN_1961;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_918 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_918 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_918 <= _GEN_1962;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_919 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_919 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_919 <= _GEN_1963;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_920 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_920 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_920 <= _GEN_1964;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_921 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_921 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_921 <= _GEN_1965;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_922 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_922 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_922 <= _GEN_1966;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_923 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_923 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_923 <= _GEN_1967;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_924 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_924 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_924 <= _GEN_1968;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_925 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_925 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_925 <= _GEN_1969;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_926 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_926 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_926 <= _GEN_1970;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_927 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_927 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_927 <= _GEN_1971;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_928 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_928 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_928 <= _GEN_1972;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_929 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_929 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_929 <= _GEN_1973;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_930 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_930 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_930 <= _GEN_1974;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_931 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_931 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_931 <= _GEN_1975;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_932 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_932 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_932 <= _GEN_1976;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_933 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_933 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_933 <= _GEN_1977;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_934 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_934 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_934 <= _GEN_1978;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_935 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_935 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_935 <= _GEN_1979;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_936 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_936 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_936 <= _GEN_1980;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_937 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_937 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_937 <= _GEN_1981;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_938 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_938 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_938 <= _GEN_1982;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_939 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_939 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_939 <= _GEN_1983;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_940 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_940 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_940 <= _GEN_1984;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_941 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_941 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_941 <= _GEN_1985;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_942 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_942 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_942 <= _GEN_1986;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_943 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_943 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_943 <= _GEN_1987;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_944 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_944 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_944 <= _GEN_1988;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_945 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_945 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_945 <= _GEN_1989;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_946 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_946 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_946 <= _GEN_1990;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_947 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_947 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_947 <= _GEN_1991;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_948 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_948 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_948 <= _GEN_1992;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_949 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_949 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_949 <= _GEN_1993;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_950 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_950 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_950 <= _GEN_1994;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_951 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_951 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_951 <= _GEN_1995;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_952 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_952 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_952 <= _GEN_1996;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_953 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_953 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_953 <= _GEN_1997;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_954 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_954 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_954 <= _GEN_1998;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_955 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_955 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_955 <= _GEN_1999;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_956 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_956 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_956 <= _GEN_2000;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_957 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_957 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_957 <= _GEN_2001;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_958 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_958 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_958 <= _GEN_2002;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_959 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_959 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_959 <= _GEN_2003;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_960 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_960 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_960 <= _GEN_2004;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_961 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_961 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_961 <= _GEN_2005;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_962 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_962 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_962 <= _GEN_2006;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_963 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_963 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_963 <= _GEN_2007;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_964 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_964 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_964 <= _GEN_2008;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_965 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_965 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_965 <= _GEN_2009;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_966 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_966 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_966 <= _GEN_2010;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_967 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_967 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_967 <= _GEN_2011;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_968 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_968 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_968 <= _GEN_2012;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_969 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_969 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_969 <= _GEN_2013;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_970 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_970 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_970 <= _GEN_2014;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_971 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_971 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_971 <= _GEN_2015;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_972 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_972 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_972 <= _GEN_2016;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_973 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_973 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_973 <= _GEN_2017;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_974 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_974 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_974 <= _GEN_2018;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_975 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_975 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_975 <= _GEN_2019;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_976 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_976 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_976 <= _GEN_2020;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_977 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_977 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_977 <= _GEN_2021;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_978 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_978 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_978 <= _GEN_2022;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_979 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_979 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_979 <= _GEN_2023;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_980 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_980 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_980 <= _GEN_2024;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_981 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_981 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_981 <= _GEN_2025;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_982 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_982 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_982 <= _GEN_2026;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_983 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_983 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_983 <= _GEN_2027;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_984 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_984 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_984 <= _GEN_2028;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_985 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_985 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_985 <= _GEN_2029;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_986 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_986 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_986 <= _GEN_2030;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_987 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_987 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_987 <= _GEN_2031;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_988 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_988 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_988 <= _GEN_2032;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_989 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_989 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_989 <= _GEN_2033;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_990 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_990 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_990 <= _GEN_2034;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_991 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_991 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_991 <= _GEN_2035;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_992 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_992 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_992 <= _GEN_2036;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_993 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_993 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_993 <= _GEN_2037;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_994 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_994 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_994 <= _GEN_2038;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_995 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_995 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_995 <= _GEN_2039;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_996 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_996 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_996 <= _GEN_2040;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_997 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_997 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_997 <= _GEN_2041;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_998 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_998 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_998 <= _GEN_2042;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_999 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_999 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_999 <= _GEN_2043;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_1000 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_1000 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_1000 <= _GEN_2044;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_1001 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_1001 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_1001 <= _GEN_2045;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_1002 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_1002 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_1002 <= _GEN_2046;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_1003 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_1003 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_1003 <= _GEN_2047;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_1004 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_1004 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_1004 <= _GEN_2048;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_1005 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_1005 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_1005 <= _GEN_2049;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_1006 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_1006 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_1006 <= _GEN_2050;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_1007 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_1007 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_1007 <= _GEN_2051;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_1008 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_1008 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_1008 <= _GEN_2052;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_1009 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_1009 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_1009 <= _GEN_2053;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_1010 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_1010 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_1010 <= _GEN_2054;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_1011 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_1011 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_1011 <= _GEN_2055;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_1012 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_1012 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_1012 <= _GEN_2056;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_1013 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_1013 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_1013 <= _GEN_2057;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_1014 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_1014 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_1014 <= _GEN_2058;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_1015 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_1015 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_1015 <= _GEN_2059;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_1016 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_1016 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_1016 <= _GEN_2060;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_1017 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_1017 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_1017 <= _GEN_2061;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_1018 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_1018 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_1018 <= _GEN_2062;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_1019 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_1019 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_1019 <= _GEN_2063;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_1020 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_1020 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_1020 <= _GEN_2064;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_1021 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_1021 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_1021 <= _GEN_2065;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_1022 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_1022 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_1022 <= _GEN_2066;
    end
    if (reset) begin // @[ICache.scala 51:22]
      valid_1023 <= 1'h0; // @[ICache.scala 51:22]
    end else if (io_fence_i) begin // @[ICache.scala 161:20]
      valid_1023 <= 1'h0; // @[ICache.scala 163:16]
    end else if (_array_io_en_T) begin // @[ICache.scala 124:19]
      valid_1023 <= _GEN_2067;
    end
    if (reset) begin // @[ICache.scala 78:68]
      state <= 3'h4; // @[ICache.scala 78:68]
    end else if (3'h0 == state) begin // @[ICache.scala 80:17]
      if (_state_T & ~_state_T_1) begin // @[ICache.scala 82:19]
        state <= 3'h4;
      end else if (array_hit) begin // @[ICache.scala 82:55]
        state <= 3'h0;
      end else begin
        state <= 3'h1;
      end
    end else if (3'h1 == state) begin // @[ICache.scala 80:17]
      if (_T_2) begin // @[ICache.scala 85:23]
        state <= 3'h2; // @[ICache.scala 86:15]
      end
    end else if (3'h2 == state) begin // @[ICache.scala 80:17]
      state <= _GEN_1034;
    end else begin
      state <= _GEN_1038;
    end
    array_out_REG <= io_cache_req_valid & s2_ready; // @[ICache.scala 56:27]
    if (reset) begin // @[Reg.scala 35:20]
      array_out_r <= 273'h0; // @[Reg.scala 35:20]
    end else if (array_out_REG) begin // @[Utils.scala 50:8]
      array_out_r <= array_io_rdata;
    end
    array_data_REG <= io_cache_req_ready & io_cache_req_valid; // @[Decoupled.scala 51:35]
    if (reset) begin // @[Reg.scala 35:20]
      array_data_r <= 64'h0; // @[Reg.scala 35:20]
    end else if (array_data_REG) begin // @[Reg.scala 36:18]
      if (2'h3 == req_r_addr[4:3]) begin // @[Mux.scala 81:58]
        array_data_r <= array_out_data[255:192];
      end else if (2'h2 == req_r_addr[4:3]) begin // @[Mux.scala 81:58]
        array_data_r <= array_out_data[191:128];
      end else begin
        array_data_r <= _array_data_T_6;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      wdata <= 256'h0; // @[Reg.scala 35:20]
    end else if (_array_io_en_T) begin // @[Reg.scala 36:18]
      wdata <= auto_out_d_bits_data; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Counter.scala 61:40]
      source <= 2'h0; // @[Counter.scala 61:40]
    end else if (_T_2) begin // @[Counter.scala 118:16]
      source <= _source_wrap_value_T_1; // @[Counter.scala 77:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  req_r_addr = _RAND_0[38:0];
  _RAND_1 = {1{`RANDOM}};
  valid_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  valid_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  valid_2 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  valid_3 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  valid_4 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  valid_5 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  valid_6 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  valid_7 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  valid_8 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  valid_9 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  valid_10 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  valid_11 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  valid_12 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  valid_13 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  valid_14 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  valid_15 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  valid_16 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  valid_17 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  valid_18 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  valid_19 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  valid_20 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  valid_21 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  valid_22 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  valid_23 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  valid_24 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  valid_25 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  valid_26 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  valid_27 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  valid_28 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  valid_29 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  valid_30 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  valid_31 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  valid_32 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  valid_33 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  valid_34 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  valid_35 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  valid_36 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  valid_37 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  valid_38 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  valid_39 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  valid_40 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  valid_41 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  valid_42 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  valid_43 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  valid_44 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  valid_45 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  valid_46 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  valid_47 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  valid_48 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  valid_49 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  valid_50 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  valid_51 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  valid_52 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  valid_53 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  valid_54 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  valid_55 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  valid_56 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  valid_57 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  valid_58 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  valid_59 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  valid_60 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  valid_61 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  valid_62 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  valid_63 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  valid_64 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  valid_65 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  valid_66 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  valid_67 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  valid_68 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  valid_69 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  valid_70 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  valid_71 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  valid_72 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  valid_73 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  valid_74 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  valid_75 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  valid_76 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  valid_77 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  valid_78 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  valid_79 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  valid_80 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  valid_81 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  valid_82 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  valid_83 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  valid_84 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  valid_85 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  valid_86 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  valid_87 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  valid_88 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  valid_89 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  valid_90 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  valid_91 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  valid_92 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  valid_93 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  valid_94 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  valid_95 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  valid_96 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  valid_97 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  valid_98 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  valid_99 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  valid_100 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  valid_101 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  valid_102 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  valid_103 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  valid_104 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  valid_105 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  valid_106 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  valid_107 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  valid_108 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  valid_109 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  valid_110 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  valid_111 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  valid_112 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  valid_113 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  valid_114 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  valid_115 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  valid_116 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  valid_117 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  valid_118 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  valid_119 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  valid_120 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  valid_121 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  valid_122 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  valid_123 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  valid_124 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  valid_125 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  valid_126 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  valid_127 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  valid_128 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  valid_129 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  valid_130 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  valid_131 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  valid_132 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  valid_133 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  valid_134 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  valid_135 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  valid_136 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  valid_137 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  valid_138 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  valid_139 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  valid_140 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  valid_141 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  valid_142 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  valid_143 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  valid_144 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  valid_145 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  valid_146 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  valid_147 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  valid_148 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  valid_149 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  valid_150 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  valid_151 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  valid_152 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  valid_153 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  valid_154 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  valid_155 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  valid_156 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  valid_157 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  valid_158 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  valid_159 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  valid_160 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  valid_161 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  valid_162 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  valid_163 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  valid_164 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  valid_165 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  valid_166 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  valid_167 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  valid_168 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  valid_169 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  valid_170 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  valid_171 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  valid_172 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  valid_173 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  valid_174 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  valid_175 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  valid_176 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  valid_177 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  valid_178 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  valid_179 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  valid_180 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  valid_181 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  valid_182 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  valid_183 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  valid_184 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  valid_185 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  valid_186 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  valid_187 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  valid_188 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  valid_189 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  valid_190 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  valid_191 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  valid_192 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  valid_193 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  valid_194 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  valid_195 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  valid_196 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  valid_197 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  valid_198 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  valid_199 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  valid_200 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  valid_201 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  valid_202 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  valid_203 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  valid_204 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  valid_205 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  valid_206 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  valid_207 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  valid_208 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  valid_209 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  valid_210 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  valid_211 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  valid_212 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  valid_213 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  valid_214 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  valid_215 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  valid_216 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  valid_217 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  valid_218 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  valid_219 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  valid_220 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  valid_221 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  valid_222 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  valid_223 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  valid_224 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  valid_225 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  valid_226 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  valid_227 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  valid_228 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  valid_229 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  valid_230 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  valid_231 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  valid_232 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  valid_233 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  valid_234 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  valid_235 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  valid_236 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  valid_237 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  valid_238 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  valid_239 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  valid_240 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  valid_241 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  valid_242 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  valid_243 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  valid_244 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  valid_245 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  valid_246 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  valid_247 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  valid_248 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  valid_249 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  valid_250 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  valid_251 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  valid_252 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  valid_253 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  valid_254 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  valid_255 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  valid_256 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  valid_257 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  valid_258 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  valid_259 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  valid_260 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  valid_261 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  valid_262 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  valid_263 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  valid_264 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  valid_265 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  valid_266 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  valid_267 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  valid_268 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  valid_269 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  valid_270 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  valid_271 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  valid_272 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  valid_273 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  valid_274 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  valid_275 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  valid_276 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  valid_277 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  valid_278 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  valid_279 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  valid_280 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  valid_281 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  valid_282 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  valid_283 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  valid_284 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  valid_285 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  valid_286 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  valid_287 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  valid_288 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  valid_289 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  valid_290 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  valid_291 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  valid_292 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  valid_293 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  valid_294 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  valid_295 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  valid_296 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  valid_297 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  valid_298 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  valid_299 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  valid_300 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  valid_301 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  valid_302 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  valid_303 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  valid_304 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  valid_305 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  valid_306 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  valid_307 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  valid_308 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  valid_309 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  valid_310 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  valid_311 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  valid_312 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  valid_313 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  valid_314 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  valid_315 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  valid_316 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  valid_317 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  valid_318 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  valid_319 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  valid_320 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  valid_321 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  valid_322 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  valid_323 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  valid_324 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  valid_325 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  valid_326 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  valid_327 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  valid_328 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  valid_329 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  valid_330 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  valid_331 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  valid_332 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  valid_333 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  valid_334 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  valid_335 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  valid_336 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  valid_337 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  valid_338 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  valid_339 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  valid_340 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  valid_341 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  valid_342 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  valid_343 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  valid_344 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  valid_345 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  valid_346 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  valid_347 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  valid_348 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  valid_349 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  valid_350 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  valid_351 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  valid_352 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  valid_353 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  valid_354 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  valid_355 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  valid_356 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  valid_357 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  valid_358 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  valid_359 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  valid_360 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  valid_361 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  valid_362 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  valid_363 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  valid_364 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  valid_365 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  valid_366 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  valid_367 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  valid_368 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  valid_369 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  valid_370 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  valid_371 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  valid_372 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  valid_373 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  valid_374 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  valid_375 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  valid_376 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  valid_377 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  valid_378 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  valid_379 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  valid_380 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  valid_381 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  valid_382 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  valid_383 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  valid_384 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  valid_385 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  valid_386 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  valid_387 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  valid_388 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  valid_389 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  valid_390 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  valid_391 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  valid_392 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  valid_393 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  valid_394 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  valid_395 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  valid_396 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  valid_397 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  valid_398 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  valid_399 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  valid_400 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  valid_401 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  valid_402 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  valid_403 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  valid_404 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  valid_405 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  valid_406 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  valid_407 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  valid_408 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  valid_409 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  valid_410 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  valid_411 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  valid_412 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  valid_413 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  valid_414 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  valid_415 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  valid_416 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  valid_417 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  valid_418 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  valid_419 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  valid_420 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  valid_421 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  valid_422 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  valid_423 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  valid_424 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  valid_425 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  valid_426 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  valid_427 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  valid_428 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  valid_429 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  valid_430 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  valid_431 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  valid_432 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  valid_433 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  valid_434 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  valid_435 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  valid_436 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  valid_437 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  valid_438 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  valid_439 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  valid_440 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  valid_441 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  valid_442 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  valid_443 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  valid_444 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  valid_445 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  valid_446 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  valid_447 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  valid_448 = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  valid_449 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  valid_450 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  valid_451 = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  valid_452 = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  valid_453 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  valid_454 = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  valid_455 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  valid_456 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  valid_457 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  valid_458 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  valid_459 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  valid_460 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  valid_461 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  valid_462 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  valid_463 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  valid_464 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  valid_465 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  valid_466 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  valid_467 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  valid_468 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  valid_469 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  valid_470 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  valid_471 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  valid_472 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  valid_473 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  valid_474 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  valid_475 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  valid_476 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  valid_477 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  valid_478 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  valid_479 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  valid_480 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  valid_481 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  valid_482 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  valid_483 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  valid_484 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  valid_485 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  valid_486 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  valid_487 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  valid_488 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  valid_489 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  valid_490 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  valid_491 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  valid_492 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  valid_493 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  valid_494 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  valid_495 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  valid_496 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  valid_497 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  valid_498 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  valid_499 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  valid_500 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  valid_501 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  valid_502 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  valid_503 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  valid_504 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  valid_505 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  valid_506 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  valid_507 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  valid_508 = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  valid_509 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  valid_510 = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  valid_511 = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  valid_512 = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  valid_513 = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  valid_514 = _RAND_515[0:0];
  _RAND_516 = {1{`RANDOM}};
  valid_515 = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  valid_516 = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  valid_517 = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  valid_518 = _RAND_519[0:0];
  _RAND_520 = {1{`RANDOM}};
  valid_519 = _RAND_520[0:0];
  _RAND_521 = {1{`RANDOM}};
  valid_520 = _RAND_521[0:0];
  _RAND_522 = {1{`RANDOM}};
  valid_521 = _RAND_522[0:0];
  _RAND_523 = {1{`RANDOM}};
  valid_522 = _RAND_523[0:0];
  _RAND_524 = {1{`RANDOM}};
  valid_523 = _RAND_524[0:0];
  _RAND_525 = {1{`RANDOM}};
  valid_524 = _RAND_525[0:0];
  _RAND_526 = {1{`RANDOM}};
  valid_525 = _RAND_526[0:0];
  _RAND_527 = {1{`RANDOM}};
  valid_526 = _RAND_527[0:0];
  _RAND_528 = {1{`RANDOM}};
  valid_527 = _RAND_528[0:0];
  _RAND_529 = {1{`RANDOM}};
  valid_528 = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  valid_529 = _RAND_530[0:0];
  _RAND_531 = {1{`RANDOM}};
  valid_530 = _RAND_531[0:0];
  _RAND_532 = {1{`RANDOM}};
  valid_531 = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  valid_532 = _RAND_533[0:0];
  _RAND_534 = {1{`RANDOM}};
  valid_533 = _RAND_534[0:0];
  _RAND_535 = {1{`RANDOM}};
  valid_534 = _RAND_535[0:0];
  _RAND_536 = {1{`RANDOM}};
  valid_535 = _RAND_536[0:0];
  _RAND_537 = {1{`RANDOM}};
  valid_536 = _RAND_537[0:0];
  _RAND_538 = {1{`RANDOM}};
  valid_537 = _RAND_538[0:0];
  _RAND_539 = {1{`RANDOM}};
  valid_538 = _RAND_539[0:0];
  _RAND_540 = {1{`RANDOM}};
  valid_539 = _RAND_540[0:0];
  _RAND_541 = {1{`RANDOM}};
  valid_540 = _RAND_541[0:0];
  _RAND_542 = {1{`RANDOM}};
  valid_541 = _RAND_542[0:0];
  _RAND_543 = {1{`RANDOM}};
  valid_542 = _RAND_543[0:0];
  _RAND_544 = {1{`RANDOM}};
  valid_543 = _RAND_544[0:0];
  _RAND_545 = {1{`RANDOM}};
  valid_544 = _RAND_545[0:0];
  _RAND_546 = {1{`RANDOM}};
  valid_545 = _RAND_546[0:0];
  _RAND_547 = {1{`RANDOM}};
  valid_546 = _RAND_547[0:0];
  _RAND_548 = {1{`RANDOM}};
  valid_547 = _RAND_548[0:0];
  _RAND_549 = {1{`RANDOM}};
  valid_548 = _RAND_549[0:0];
  _RAND_550 = {1{`RANDOM}};
  valid_549 = _RAND_550[0:0];
  _RAND_551 = {1{`RANDOM}};
  valid_550 = _RAND_551[0:0];
  _RAND_552 = {1{`RANDOM}};
  valid_551 = _RAND_552[0:0];
  _RAND_553 = {1{`RANDOM}};
  valid_552 = _RAND_553[0:0];
  _RAND_554 = {1{`RANDOM}};
  valid_553 = _RAND_554[0:0];
  _RAND_555 = {1{`RANDOM}};
  valid_554 = _RAND_555[0:0];
  _RAND_556 = {1{`RANDOM}};
  valid_555 = _RAND_556[0:0];
  _RAND_557 = {1{`RANDOM}};
  valid_556 = _RAND_557[0:0];
  _RAND_558 = {1{`RANDOM}};
  valid_557 = _RAND_558[0:0];
  _RAND_559 = {1{`RANDOM}};
  valid_558 = _RAND_559[0:0];
  _RAND_560 = {1{`RANDOM}};
  valid_559 = _RAND_560[0:0];
  _RAND_561 = {1{`RANDOM}};
  valid_560 = _RAND_561[0:0];
  _RAND_562 = {1{`RANDOM}};
  valid_561 = _RAND_562[0:0];
  _RAND_563 = {1{`RANDOM}};
  valid_562 = _RAND_563[0:0];
  _RAND_564 = {1{`RANDOM}};
  valid_563 = _RAND_564[0:0];
  _RAND_565 = {1{`RANDOM}};
  valid_564 = _RAND_565[0:0];
  _RAND_566 = {1{`RANDOM}};
  valid_565 = _RAND_566[0:0];
  _RAND_567 = {1{`RANDOM}};
  valid_566 = _RAND_567[0:0];
  _RAND_568 = {1{`RANDOM}};
  valid_567 = _RAND_568[0:0];
  _RAND_569 = {1{`RANDOM}};
  valid_568 = _RAND_569[0:0];
  _RAND_570 = {1{`RANDOM}};
  valid_569 = _RAND_570[0:0];
  _RAND_571 = {1{`RANDOM}};
  valid_570 = _RAND_571[0:0];
  _RAND_572 = {1{`RANDOM}};
  valid_571 = _RAND_572[0:0];
  _RAND_573 = {1{`RANDOM}};
  valid_572 = _RAND_573[0:0];
  _RAND_574 = {1{`RANDOM}};
  valid_573 = _RAND_574[0:0];
  _RAND_575 = {1{`RANDOM}};
  valid_574 = _RAND_575[0:0];
  _RAND_576 = {1{`RANDOM}};
  valid_575 = _RAND_576[0:0];
  _RAND_577 = {1{`RANDOM}};
  valid_576 = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  valid_577 = _RAND_578[0:0];
  _RAND_579 = {1{`RANDOM}};
  valid_578 = _RAND_579[0:0];
  _RAND_580 = {1{`RANDOM}};
  valid_579 = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  valid_580 = _RAND_581[0:0];
  _RAND_582 = {1{`RANDOM}};
  valid_581 = _RAND_582[0:0];
  _RAND_583 = {1{`RANDOM}};
  valid_582 = _RAND_583[0:0];
  _RAND_584 = {1{`RANDOM}};
  valid_583 = _RAND_584[0:0];
  _RAND_585 = {1{`RANDOM}};
  valid_584 = _RAND_585[0:0];
  _RAND_586 = {1{`RANDOM}};
  valid_585 = _RAND_586[0:0];
  _RAND_587 = {1{`RANDOM}};
  valid_586 = _RAND_587[0:0];
  _RAND_588 = {1{`RANDOM}};
  valid_587 = _RAND_588[0:0];
  _RAND_589 = {1{`RANDOM}};
  valid_588 = _RAND_589[0:0];
  _RAND_590 = {1{`RANDOM}};
  valid_589 = _RAND_590[0:0];
  _RAND_591 = {1{`RANDOM}};
  valid_590 = _RAND_591[0:0];
  _RAND_592 = {1{`RANDOM}};
  valid_591 = _RAND_592[0:0];
  _RAND_593 = {1{`RANDOM}};
  valid_592 = _RAND_593[0:0];
  _RAND_594 = {1{`RANDOM}};
  valid_593 = _RAND_594[0:0];
  _RAND_595 = {1{`RANDOM}};
  valid_594 = _RAND_595[0:0];
  _RAND_596 = {1{`RANDOM}};
  valid_595 = _RAND_596[0:0];
  _RAND_597 = {1{`RANDOM}};
  valid_596 = _RAND_597[0:0];
  _RAND_598 = {1{`RANDOM}};
  valid_597 = _RAND_598[0:0];
  _RAND_599 = {1{`RANDOM}};
  valid_598 = _RAND_599[0:0];
  _RAND_600 = {1{`RANDOM}};
  valid_599 = _RAND_600[0:0];
  _RAND_601 = {1{`RANDOM}};
  valid_600 = _RAND_601[0:0];
  _RAND_602 = {1{`RANDOM}};
  valid_601 = _RAND_602[0:0];
  _RAND_603 = {1{`RANDOM}};
  valid_602 = _RAND_603[0:0];
  _RAND_604 = {1{`RANDOM}};
  valid_603 = _RAND_604[0:0];
  _RAND_605 = {1{`RANDOM}};
  valid_604 = _RAND_605[0:0];
  _RAND_606 = {1{`RANDOM}};
  valid_605 = _RAND_606[0:0];
  _RAND_607 = {1{`RANDOM}};
  valid_606 = _RAND_607[0:0];
  _RAND_608 = {1{`RANDOM}};
  valid_607 = _RAND_608[0:0];
  _RAND_609 = {1{`RANDOM}};
  valid_608 = _RAND_609[0:0];
  _RAND_610 = {1{`RANDOM}};
  valid_609 = _RAND_610[0:0];
  _RAND_611 = {1{`RANDOM}};
  valid_610 = _RAND_611[0:0];
  _RAND_612 = {1{`RANDOM}};
  valid_611 = _RAND_612[0:0];
  _RAND_613 = {1{`RANDOM}};
  valid_612 = _RAND_613[0:0];
  _RAND_614 = {1{`RANDOM}};
  valid_613 = _RAND_614[0:0];
  _RAND_615 = {1{`RANDOM}};
  valid_614 = _RAND_615[0:0];
  _RAND_616 = {1{`RANDOM}};
  valid_615 = _RAND_616[0:0];
  _RAND_617 = {1{`RANDOM}};
  valid_616 = _RAND_617[0:0];
  _RAND_618 = {1{`RANDOM}};
  valid_617 = _RAND_618[0:0];
  _RAND_619 = {1{`RANDOM}};
  valid_618 = _RAND_619[0:0];
  _RAND_620 = {1{`RANDOM}};
  valid_619 = _RAND_620[0:0];
  _RAND_621 = {1{`RANDOM}};
  valid_620 = _RAND_621[0:0];
  _RAND_622 = {1{`RANDOM}};
  valid_621 = _RAND_622[0:0];
  _RAND_623 = {1{`RANDOM}};
  valid_622 = _RAND_623[0:0];
  _RAND_624 = {1{`RANDOM}};
  valid_623 = _RAND_624[0:0];
  _RAND_625 = {1{`RANDOM}};
  valid_624 = _RAND_625[0:0];
  _RAND_626 = {1{`RANDOM}};
  valid_625 = _RAND_626[0:0];
  _RAND_627 = {1{`RANDOM}};
  valid_626 = _RAND_627[0:0];
  _RAND_628 = {1{`RANDOM}};
  valid_627 = _RAND_628[0:0];
  _RAND_629 = {1{`RANDOM}};
  valid_628 = _RAND_629[0:0];
  _RAND_630 = {1{`RANDOM}};
  valid_629 = _RAND_630[0:0];
  _RAND_631 = {1{`RANDOM}};
  valid_630 = _RAND_631[0:0];
  _RAND_632 = {1{`RANDOM}};
  valid_631 = _RAND_632[0:0];
  _RAND_633 = {1{`RANDOM}};
  valid_632 = _RAND_633[0:0];
  _RAND_634 = {1{`RANDOM}};
  valid_633 = _RAND_634[0:0];
  _RAND_635 = {1{`RANDOM}};
  valid_634 = _RAND_635[0:0];
  _RAND_636 = {1{`RANDOM}};
  valid_635 = _RAND_636[0:0];
  _RAND_637 = {1{`RANDOM}};
  valid_636 = _RAND_637[0:0];
  _RAND_638 = {1{`RANDOM}};
  valid_637 = _RAND_638[0:0];
  _RAND_639 = {1{`RANDOM}};
  valid_638 = _RAND_639[0:0];
  _RAND_640 = {1{`RANDOM}};
  valid_639 = _RAND_640[0:0];
  _RAND_641 = {1{`RANDOM}};
  valid_640 = _RAND_641[0:0];
  _RAND_642 = {1{`RANDOM}};
  valid_641 = _RAND_642[0:0];
  _RAND_643 = {1{`RANDOM}};
  valid_642 = _RAND_643[0:0];
  _RAND_644 = {1{`RANDOM}};
  valid_643 = _RAND_644[0:0];
  _RAND_645 = {1{`RANDOM}};
  valid_644 = _RAND_645[0:0];
  _RAND_646 = {1{`RANDOM}};
  valid_645 = _RAND_646[0:0];
  _RAND_647 = {1{`RANDOM}};
  valid_646 = _RAND_647[0:0];
  _RAND_648 = {1{`RANDOM}};
  valid_647 = _RAND_648[0:0];
  _RAND_649 = {1{`RANDOM}};
  valid_648 = _RAND_649[0:0];
  _RAND_650 = {1{`RANDOM}};
  valid_649 = _RAND_650[0:0];
  _RAND_651 = {1{`RANDOM}};
  valid_650 = _RAND_651[0:0];
  _RAND_652 = {1{`RANDOM}};
  valid_651 = _RAND_652[0:0];
  _RAND_653 = {1{`RANDOM}};
  valid_652 = _RAND_653[0:0];
  _RAND_654 = {1{`RANDOM}};
  valid_653 = _RAND_654[0:0];
  _RAND_655 = {1{`RANDOM}};
  valid_654 = _RAND_655[0:0];
  _RAND_656 = {1{`RANDOM}};
  valid_655 = _RAND_656[0:0];
  _RAND_657 = {1{`RANDOM}};
  valid_656 = _RAND_657[0:0];
  _RAND_658 = {1{`RANDOM}};
  valid_657 = _RAND_658[0:0];
  _RAND_659 = {1{`RANDOM}};
  valid_658 = _RAND_659[0:0];
  _RAND_660 = {1{`RANDOM}};
  valid_659 = _RAND_660[0:0];
  _RAND_661 = {1{`RANDOM}};
  valid_660 = _RAND_661[0:0];
  _RAND_662 = {1{`RANDOM}};
  valid_661 = _RAND_662[0:0];
  _RAND_663 = {1{`RANDOM}};
  valid_662 = _RAND_663[0:0];
  _RAND_664 = {1{`RANDOM}};
  valid_663 = _RAND_664[0:0];
  _RAND_665 = {1{`RANDOM}};
  valid_664 = _RAND_665[0:0];
  _RAND_666 = {1{`RANDOM}};
  valid_665 = _RAND_666[0:0];
  _RAND_667 = {1{`RANDOM}};
  valid_666 = _RAND_667[0:0];
  _RAND_668 = {1{`RANDOM}};
  valid_667 = _RAND_668[0:0];
  _RAND_669 = {1{`RANDOM}};
  valid_668 = _RAND_669[0:0];
  _RAND_670 = {1{`RANDOM}};
  valid_669 = _RAND_670[0:0];
  _RAND_671 = {1{`RANDOM}};
  valid_670 = _RAND_671[0:0];
  _RAND_672 = {1{`RANDOM}};
  valid_671 = _RAND_672[0:0];
  _RAND_673 = {1{`RANDOM}};
  valid_672 = _RAND_673[0:0];
  _RAND_674 = {1{`RANDOM}};
  valid_673 = _RAND_674[0:0];
  _RAND_675 = {1{`RANDOM}};
  valid_674 = _RAND_675[0:0];
  _RAND_676 = {1{`RANDOM}};
  valid_675 = _RAND_676[0:0];
  _RAND_677 = {1{`RANDOM}};
  valid_676 = _RAND_677[0:0];
  _RAND_678 = {1{`RANDOM}};
  valid_677 = _RAND_678[0:0];
  _RAND_679 = {1{`RANDOM}};
  valid_678 = _RAND_679[0:0];
  _RAND_680 = {1{`RANDOM}};
  valid_679 = _RAND_680[0:0];
  _RAND_681 = {1{`RANDOM}};
  valid_680 = _RAND_681[0:0];
  _RAND_682 = {1{`RANDOM}};
  valid_681 = _RAND_682[0:0];
  _RAND_683 = {1{`RANDOM}};
  valid_682 = _RAND_683[0:0];
  _RAND_684 = {1{`RANDOM}};
  valid_683 = _RAND_684[0:0];
  _RAND_685 = {1{`RANDOM}};
  valid_684 = _RAND_685[0:0];
  _RAND_686 = {1{`RANDOM}};
  valid_685 = _RAND_686[0:0];
  _RAND_687 = {1{`RANDOM}};
  valid_686 = _RAND_687[0:0];
  _RAND_688 = {1{`RANDOM}};
  valid_687 = _RAND_688[0:0];
  _RAND_689 = {1{`RANDOM}};
  valid_688 = _RAND_689[0:0];
  _RAND_690 = {1{`RANDOM}};
  valid_689 = _RAND_690[0:0];
  _RAND_691 = {1{`RANDOM}};
  valid_690 = _RAND_691[0:0];
  _RAND_692 = {1{`RANDOM}};
  valid_691 = _RAND_692[0:0];
  _RAND_693 = {1{`RANDOM}};
  valid_692 = _RAND_693[0:0];
  _RAND_694 = {1{`RANDOM}};
  valid_693 = _RAND_694[0:0];
  _RAND_695 = {1{`RANDOM}};
  valid_694 = _RAND_695[0:0];
  _RAND_696 = {1{`RANDOM}};
  valid_695 = _RAND_696[0:0];
  _RAND_697 = {1{`RANDOM}};
  valid_696 = _RAND_697[0:0];
  _RAND_698 = {1{`RANDOM}};
  valid_697 = _RAND_698[0:0];
  _RAND_699 = {1{`RANDOM}};
  valid_698 = _RAND_699[0:0];
  _RAND_700 = {1{`RANDOM}};
  valid_699 = _RAND_700[0:0];
  _RAND_701 = {1{`RANDOM}};
  valid_700 = _RAND_701[0:0];
  _RAND_702 = {1{`RANDOM}};
  valid_701 = _RAND_702[0:0];
  _RAND_703 = {1{`RANDOM}};
  valid_702 = _RAND_703[0:0];
  _RAND_704 = {1{`RANDOM}};
  valid_703 = _RAND_704[0:0];
  _RAND_705 = {1{`RANDOM}};
  valid_704 = _RAND_705[0:0];
  _RAND_706 = {1{`RANDOM}};
  valid_705 = _RAND_706[0:0];
  _RAND_707 = {1{`RANDOM}};
  valid_706 = _RAND_707[0:0];
  _RAND_708 = {1{`RANDOM}};
  valid_707 = _RAND_708[0:0];
  _RAND_709 = {1{`RANDOM}};
  valid_708 = _RAND_709[0:0];
  _RAND_710 = {1{`RANDOM}};
  valid_709 = _RAND_710[0:0];
  _RAND_711 = {1{`RANDOM}};
  valid_710 = _RAND_711[0:0];
  _RAND_712 = {1{`RANDOM}};
  valid_711 = _RAND_712[0:0];
  _RAND_713 = {1{`RANDOM}};
  valid_712 = _RAND_713[0:0];
  _RAND_714 = {1{`RANDOM}};
  valid_713 = _RAND_714[0:0];
  _RAND_715 = {1{`RANDOM}};
  valid_714 = _RAND_715[0:0];
  _RAND_716 = {1{`RANDOM}};
  valid_715 = _RAND_716[0:0];
  _RAND_717 = {1{`RANDOM}};
  valid_716 = _RAND_717[0:0];
  _RAND_718 = {1{`RANDOM}};
  valid_717 = _RAND_718[0:0];
  _RAND_719 = {1{`RANDOM}};
  valid_718 = _RAND_719[0:0];
  _RAND_720 = {1{`RANDOM}};
  valid_719 = _RAND_720[0:0];
  _RAND_721 = {1{`RANDOM}};
  valid_720 = _RAND_721[0:0];
  _RAND_722 = {1{`RANDOM}};
  valid_721 = _RAND_722[0:0];
  _RAND_723 = {1{`RANDOM}};
  valid_722 = _RAND_723[0:0];
  _RAND_724 = {1{`RANDOM}};
  valid_723 = _RAND_724[0:0];
  _RAND_725 = {1{`RANDOM}};
  valid_724 = _RAND_725[0:0];
  _RAND_726 = {1{`RANDOM}};
  valid_725 = _RAND_726[0:0];
  _RAND_727 = {1{`RANDOM}};
  valid_726 = _RAND_727[0:0];
  _RAND_728 = {1{`RANDOM}};
  valid_727 = _RAND_728[0:0];
  _RAND_729 = {1{`RANDOM}};
  valid_728 = _RAND_729[0:0];
  _RAND_730 = {1{`RANDOM}};
  valid_729 = _RAND_730[0:0];
  _RAND_731 = {1{`RANDOM}};
  valid_730 = _RAND_731[0:0];
  _RAND_732 = {1{`RANDOM}};
  valid_731 = _RAND_732[0:0];
  _RAND_733 = {1{`RANDOM}};
  valid_732 = _RAND_733[0:0];
  _RAND_734 = {1{`RANDOM}};
  valid_733 = _RAND_734[0:0];
  _RAND_735 = {1{`RANDOM}};
  valid_734 = _RAND_735[0:0];
  _RAND_736 = {1{`RANDOM}};
  valid_735 = _RAND_736[0:0];
  _RAND_737 = {1{`RANDOM}};
  valid_736 = _RAND_737[0:0];
  _RAND_738 = {1{`RANDOM}};
  valid_737 = _RAND_738[0:0];
  _RAND_739 = {1{`RANDOM}};
  valid_738 = _RAND_739[0:0];
  _RAND_740 = {1{`RANDOM}};
  valid_739 = _RAND_740[0:0];
  _RAND_741 = {1{`RANDOM}};
  valid_740 = _RAND_741[0:0];
  _RAND_742 = {1{`RANDOM}};
  valid_741 = _RAND_742[0:0];
  _RAND_743 = {1{`RANDOM}};
  valid_742 = _RAND_743[0:0];
  _RAND_744 = {1{`RANDOM}};
  valid_743 = _RAND_744[0:0];
  _RAND_745 = {1{`RANDOM}};
  valid_744 = _RAND_745[0:0];
  _RAND_746 = {1{`RANDOM}};
  valid_745 = _RAND_746[0:0];
  _RAND_747 = {1{`RANDOM}};
  valid_746 = _RAND_747[0:0];
  _RAND_748 = {1{`RANDOM}};
  valid_747 = _RAND_748[0:0];
  _RAND_749 = {1{`RANDOM}};
  valid_748 = _RAND_749[0:0];
  _RAND_750 = {1{`RANDOM}};
  valid_749 = _RAND_750[0:0];
  _RAND_751 = {1{`RANDOM}};
  valid_750 = _RAND_751[0:0];
  _RAND_752 = {1{`RANDOM}};
  valid_751 = _RAND_752[0:0];
  _RAND_753 = {1{`RANDOM}};
  valid_752 = _RAND_753[0:0];
  _RAND_754 = {1{`RANDOM}};
  valid_753 = _RAND_754[0:0];
  _RAND_755 = {1{`RANDOM}};
  valid_754 = _RAND_755[0:0];
  _RAND_756 = {1{`RANDOM}};
  valid_755 = _RAND_756[0:0];
  _RAND_757 = {1{`RANDOM}};
  valid_756 = _RAND_757[0:0];
  _RAND_758 = {1{`RANDOM}};
  valid_757 = _RAND_758[0:0];
  _RAND_759 = {1{`RANDOM}};
  valid_758 = _RAND_759[0:0];
  _RAND_760 = {1{`RANDOM}};
  valid_759 = _RAND_760[0:0];
  _RAND_761 = {1{`RANDOM}};
  valid_760 = _RAND_761[0:0];
  _RAND_762 = {1{`RANDOM}};
  valid_761 = _RAND_762[0:0];
  _RAND_763 = {1{`RANDOM}};
  valid_762 = _RAND_763[0:0];
  _RAND_764 = {1{`RANDOM}};
  valid_763 = _RAND_764[0:0];
  _RAND_765 = {1{`RANDOM}};
  valid_764 = _RAND_765[0:0];
  _RAND_766 = {1{`RANDOM}};
  valid_765 = _RAND_766[0:0];
  _RAND_767 = {1{`RANDOM}};
  valid_766 = _RAND_767[0:0];
  _RAND_768 = {1{`RANDOM}};
  valid_767 = _RAND_768[0:0];
  _RAND_769 = {1{`RANDOM}};
  valid_768 = _RAND_769[0:0];
  _RAND_770 = {1{`RANDOM}};
  valid_769 = _RAND_770[0:0];
  _RAND_771 = {1{`RANDOM}};
  valid_770 = _RAND_771[0:0];
  _RAND_772 = {1{`RANDOM}};
  valid_771 = _RAND_772[0:0];
  _RAND_773 = {1{`RANDOM}};
  valid_772 = _RAND_773[0:0];
  _RAND_774 = {1{`RANDOM}};
  valid_773 = _RAND_774[0:0];
  _RAND_775 = {1{`RANDOM}};
  valid_774 = _RAND_775[0:0];
  _RAND_776 = {1{`RANDOM}};
  valid_775 = _RAND_776[0:0];
  _RAND_777 = {1{`RANDOM}};
  valid_776 = _RAND_777[0:0];
  _RAND_778 = {1{`RANDOM}};
  valid_777 = _RAND_778[0:0];
  _RAND_779 = {1{`RANDOM}};
  valid_778 = _RAND_779[0:0];
  _RAND_780 = {1{`RANDOM}};
  valid_779 = _RAND_780[0:0];
  _RAND_781 = {1{`RANDOM}};
  valid_780 = _RAND_781[0:0];
  _RAND_782 = {1{`RANDOM}};
  valid_781 = _RAND_782[0:0];
  _RAND_783 = {1{`RANDOM}};
  valid_782 = _RAND_783[0:0];
  _RAND_784 = {1{`RANDOM}};
  valid_783 = _RAND_784[0:0];
  _RAND_785 = {1{`RANDOM}};
  valid_784 = _RAND_785[0:0];
  _RAND_786 = {1{`RANDOM}};
  valid_785 = _RAND_786[0:0];
  _RAND_787 = {1{`RANDOM}};
  valid_786 = _RAND_787[0:0];
  _RAND_788 = {1{`RANDOM}};
  valid_787 = _RAND_788[0:0];
  _RAND_789 = {1{`RANDOM}};
  valid_788 = _RAND_789[0:0];
  _RAND_790 = {1{`RANDOM}};
  valid_789 = _RAND_790[0:0];
  _RAND_791 = {1{`RANDOM}};
  valid_790 = _RAND_791[0:0];
  _RAND_792 = {1{`RANDOM}};
  valid_791 = _RAND_792[0:0];
  _RAND_793 = {1{`RANDOM}};
  valid_792 = _RAND_793[0:0];
  _RAND_794 = {1{`RANDOM}};
  valid_793 = _RAND_794[0:0];
  _RAND_795 = {1{`RANDOM}};
  valid_794 = _RAND_795[0:0];
  _RAND_796 = {1{`RANDOM}};
  valid_795 = _RAND_796[0:0];
  _RAND_797 = {1{`RANDOM}};
  valid_796 = _RAND_797[0:0];
  _RAND_798 = {1{`RANDOM}};
  valid_797 = _RAND_798[0:0];
  _RAND_799 = {1{`RANDOM}};
  valid_798 = _RAND_799[0:0];
  _RAND_800 = {1{`RANDOM}};
  valid_799 = _RAND_800[0:0];
  _RAND_801 = {1{`RANDOM}};
  valid_800 = _RAND_801[0:0];
  _RAND_802 = {1{`RANDOM}};
  valid_801 = _RAND_802[0:0];
  _RAND_803 = {1{`RANDOM}};
  valid_802 = _RAND_803[0:0];
  _RAND_804 = {1{`RANDOM}};
  valid_803 = _RAND_804[0:0];
  _RAND_805 = {1{`RANDOM}};
  valid_804 = _RAND_805[0:0];
  _RAND_806 = {1{`RANDOM}};
  valid_805 = _RAND_806[0:0];
  _RAND_807 = {1{`RANDOM}};
  valid_806 = _RAND_807[0:0];
  _RAND_808 = {1{`RANDOM}};
  valid_807 = _RAND_808[0:0];
  _RAND_809 = {1{`RANDOM}};
  valid_808 = _RAND_809[0:0];
  _RAND_810 = {1{`RANDOM}};
  valid_809 = _RAND_810[0:0];
  _RAND_811 = {1{`RANDOM}};
  valid_810 = _RAND_811[0:0];
  _RAND_812 = {1{`RANDOM}};
  valid_811 = _RAND_812[0:0];
  _RAND_813 = {1{`RANDOM}};
  valid_812 = _RAND_813[0:0];
  _RAND_814 = {1{`RANDOM}};
  valid_813 = _RAND_814[0:0];
  _RAND_815 = {1{`RANDOM}};
  valid_814 = _RAND_815[0:0];
  _RAND_816 = {1{`RANDOM}};
  valid_815 = _RAND_816[0:0];
  _RAND_817 = {1{`RANDOM}};
  valid_816 = _RAND_817[0:0];
  _RAND_818 = {1{`RANDOM}};
  valid_817 = _RAND_818[0:0];
  _RAND_819 = {1{`RANDOM}};
  valid_818 = _RAND_819[0:0];
  _RAND_820 = {1{`RANDOM}};
  valid_819 = _RAND_820[0:0];
  _RAND_821 = {1{`RANDOM}};
  valid_820 = _RAND_821[0:0];
  _RAND_822 = {1{`RANDOM}};
  valid_821 = _RAND_822[0:0];
  _RAND_823 = {1{`RANDOM}};
  valid_822 = _RAND_823[0:0];
  _RAND_824 = {1{`RANDOM}};
  valid_823 = _RAND_824[0:0];
  _RAND_825 = {1{`RANDOM}};
  valid_824 = _RAND_825[0:0];
  _RAND_826 = {1{`RANDOM}};
  valid_825 = _RAND_826[0:0];
  _RAND_827 = {1{`RANDOM}};
  valid_826 = _RAND_827[0:0];
  _RAND_828 = {1{`RANDOM}};
  valid_827 = _RAND_828[0:0];
  _RAND_829 = {1{`RANDOM}};
  valid_828 = _RAND_829[0:0];
  _RAND_830 = {1{`RANDOM}};
  valid_829 = _RAND_830[0:0];
  _RAND_831 = {1{`RANDOM}};
  valid_830 = _RAND_831[0:0];
  _RAND_832 = {1{`RANDOM}};
  valid_831 = _RAND_832[0:0];
  _RAND_833 = {1{`RANDOM}};
  valid_832 = _RAND_833[0:0];
  _RAND_834 = {1{`RANDOM}};
  valid_833 = _RAND_834[0:0];
  _RAND_835 = {1{`RANDOM}};
  valid_834 = _RAND_835[0:0];
  _RAND_836 = {1{`RANDOM}};
  valid_835 = _RAND_836[0:0];
  _RAND_837 = {1{`RANDOM}};
  valid_836 = _RAND_837[0:0];
  _RAND_838 = {1{`RANDOM}};
  valid_837 = _RAND_838[0:0];
  _RAND_839 = {1{`RANDOM}};
  valid_838 = _RAND_839[0:0];
  _RAND_840 = {1{`RANDOM}};
  valid_839 = _RAND_840[0:0];
  _RAND_841 = {1{`RANDOM}};
  valid_840 = _RAND_841[0:0];
  _RAND_842 = {1{`RANDOM}};
  valid_841 = _RAND_842[0:0];
  _RAND_843 = {1{`RANDOM}};
  valid_842 = _RAND_843[0:0];
  _RAND_844 = {1{`RANDOM}};
  valid_843 = _RAND_844[0:0];
  _RAND_845 = {1{`RANDOM}};
  valid_844 = _RAND_845[0:0];
  _RAND_846 = {1{`RANDOM}};
  valid_845 = _RAND_846[0:0];
  _RAND_847 = {1{`RANDOM}};
  valid_846 = _RAND_847[0:0];
  _RAND_848 = {1{`RANDOM}};
  valid_847 = _RAND_848[0:0];
  _RAND_849 = {1{`RANDOM}};
  valid_848 = _RAND_849[0:0];
  _RAND_850 = {1{`RANDOM}};
  valid_849 = _RAND_850[0:0];
  _RAND_851 = {1{`RANDOM}};
  valid_850 = _RAND_851[0:0];
  _RAND_852 = {1{`RANDOM}};
  valid_851 = _RAND_852[0:0];
  _RAND_853 = {1{`RANDOM}};
  valid_852 = _RAND_853[0:0];
  _RAND_854 = {1{`RANDOM}};
  valid_853 = _RAND_854[0:0];
  _RAND_855 = {1{`RANDOM}};
  valid_854 = _RAND_855[0:0];
  _RAND_856 = {1{`RANDOM}};
  valid_855 = _RAND_856[0:0];
  _RAND_857 = {1{`RANDOM}};
  valid_856 = _RAND_857[0:0];
  _RAND_858 = {1{`RANDOM}};
  valid_857 = _RAND_858[0:0];
  _RAND_859 = {1{`RANDOM}};
  valid_858 = _RAND_859[0:0];
  _RAND_860 = {1{`RANDOM}};
  valid_859 = _RAND_860[0:0];
  _RAND_861 = {1{`RANDOM}};
  valid_860 = _RAND_861[0:0];
  _RAND_862 = {1{`RANDOM}};
  valid_861 = _RAND_862[0:0];
  _RAND_863 = {1{`RANDOM}};
  valid_862 = _RAND_863[0:0];
  _RAND_864 = {1{`RANDOM}};
  valid_863 = _RAND_864[0:0];
  _RAND_865 = {1{`RANDOM}};
  valid_864 = _RAND_865[0:0];
  _RAND_866 = {1{`RANDOM}};
  valid_865 = _RAND_866[0:0];
  _RAND_867 = {1{`RANDOM}};
  valid_866 = _RAND_867[0:0];
  _RAND_868 = {1{`RANDOM}};
  valid_867 = _RAND_868[0:0];
  _RAND_869 = {1{`RANDOM}};
  valid_868 = _RAND_869[0:0];
  _RAND_870 = {1{`RANDOM}};
  valid_869 = _RAND_870[0:0];
  _RAND_871 = {1{`RANDOM}};
  valid_870 = _RAND_871[0:0];
  _RAND_872 = {1{`RANDOM}};
  valid_871 = _RAND_872[0:0];
  _RAND_873 = {1{`RANDOM}};
  valid_872 = _RAND_873[0:0];
  _RAND_874 = {1{`RANDOM}};
  valid_873 = _RAND_874[0:0];
  _RAND_875 = {1{`RANDOM}};
  valid_874 = _RAND_875[0:0];
  _RAND_876 = {1{`RANDOM}};
  valid_875 = _RAND_876[0:0];
  _RAND_877 = {1{`RANDOM}};
  valid_876 = _RAND_877[0:0];
  _RAND_878 = {1{`RANDOM}};
  valid_877 = _RAND_878[0:0];
  _RAND_879 = {1{`RANDOM}};
  valid_878 = _RAND_879[0:0];
  _RAND_880 = {1{`RANDOM}};
  valid_879 = _RAND_880[0:0];
  _RAND_881 = {1{`RANDOM}};
  valid_880 = _RAND_881[0:0];
  _RAND_882 = {1{`RANDOM}};
  valid_881 = _RAND_882[0:0];
  _RAND_883 = {1{`RANDOM}};
  valid_882 = _RAND_883[0:0];
  _RAND_884 = {1{`RANDOM}};
  valid_883 = _RAND_884[0:0];
  _RAND_885 = {1{`RANDOM}};
  valid_884 = _RAND_885[0:0];
  _RAND_886 = {1{`RANDOM}};
  valid_885 = _RAND_886[0:0];
  _RAND_887 = {1{`RANDOM}};
  valid_886 = _RAND_887[0:0];
  _RAND_888 = {1{`RANDOM}};
  valid_887 = _RAND_888[0:0];
  _RAND_889 = {1{`RANDOM}};
  valid_888 = _RAND_889[0:0];
  _RAND_890 = {1{`RANDOM}};
  valid_889 = _RAND_890[0:0];
  _RAND_891 = {1{`RANDOM}};
  valid_890 = _RAND_891[0:0];
  _RAND_892 = {1{`RANDOM}};
  valid_891 = _RAND_892[0:0];
  _RAND_893 = {1{`RANDOM}};
  valid_892 = _RAND_893[0:0];
  _RAND_894 = {1{`RANDOM}};
  valid_893 = _RAND_894[0:0];
  _RAND_895 = {1{`RANDOM}};
  valid_894 = _RAND_895[0:0];
  _RAND_896 = {1{`RANDOM}};
  valid_895 = _RAND_896[0:0];
  _RAND_897 = {1{`RANDOM}};
  valid_896 = _RAND_897[0:0];
  _RAND_898 = {1{`RANDOM}};
  valid_897 = _RAND_898[0:0];
  _RAND_899 = {1{`RANDOM}};
  valid_898 = _RAND_899[0:0];
  _RAND_900 = {1{`RANDOM}};
  valid_899 = _RAND_900[0:0];
  _RAND_901 = {1{`RANDOM}};
  valid_900 = _RAND_901[0:0];
  _RAND_902 = {1{`RANDOM}};
  valid_901 = _RAND_902[0:0];
  _RAND_903 = {1{`RANDOM}};
  valid_902 = _RAND_903[0:0];
  _RAND_904 = {1{`RANDOM}};
  valid_903 = _RAND_904[0:0];
  _RAND_905 = {1{`RANDOM}};
  valid_904 = _RAND_905[0:0];
  _RAND_906 = {1{`RANDOM}};
  valid_905 = _RAND_906[0:0];
  _RAND_907 = {1{`RANDOM}};
  valid_906 = _RAND_907[0:0];
  _RAND_908 = {1{`RANDOM}};
  valid_907 = _RAND_908[0:0];
  _RAND_909 = {1{`RANDOM}};
  valid_908 = _RAND_909[0:0];
  _RAND_910 = {1{`RANDOM}};
  valid_909 = _RAND_910[0:0];
  _RAND_911 = {1{`RANDOM}};
  valid_910 = _RAND_911[0:0];
  _RAND_912 = {1{`RANDOM}};
  valid_911 = _RAND_912[0:0];
  _RAND_913 = {1{`RANDOM}};
  valid_912 = _RAND_913[0:0];
  _RAND_914 = {1{`RANDOM}};
  valid_913 = _RAND_914[0:0];
  _RAND_915 = {1{`RANDOM}};
  valid_914 = _RAND_915[0:0];
  _RAND_916 = {1{`RANDOM}};
  valid_915 = _RAND_916[0:0];
  _RAND_917 = {1{`RANDOM}};
  valid_916 = _RAND_917[0:0];
  _RAND_918 = {1{`RANDOM}};
  valid_917 = _RAND_918[0:0];
  _RAND_919 = {1{`RANDOM}};
  valid_918 = _RAND_919[0:0];
  _RAND_920 = {1{`RANDOM}};
  valid_919 = _RAND_920[0:0];
  _RAND_921 = {1{`RANDOM}};
  valid_920 = _RAND_921[0:0];
  _RAND_922 = {1{`RANDOM}};
  valid_921 = _RAND_922[0:0];
  _RAND_923 = {1{`RANDOM}};
  valid_922 = _RAND_923[0:0];
  _RAND_924 = {1{`RANDOM}};
  valid_923 = _RAND_924[0:0];
  _RAND_925 = {1{`RANDOM}};
  valid_924 = _RAND_925[0:0];
  _RAND_926 = {1{`RANDOM}};
  valid_925 = _RAND_926[0:0];
  _RAND_927 = {1{`RANDOM}};
  valid_926 = _RAND_927[0:0];
  _RAND_928 = {1{`RANDOM}};
  valid_927 = _RAND_928[0:0];
  _RAND_929 = {1{`RANDOM}};
  valid_928 = _RAND_929[0:0];
  _RAND_930 = {1{`RANDOM}};
  valid_929 = _RAND_930[0:0];
  _RAND_931 = {1{`RANDOM}};
  valid_930 = _RAND_931[0:0];
  _RAND_932 = {1{`RANDOM}};
  valid_931 = _RAND_932[0:0];
  _RAND_933 = {1{`RANDOM}};
  valid_932 = _RAND_933[0:0];
  _RAND_934 = {1{`RANDOM}};
  valid_933 = _RAND_934[0:0];
  _RAND_935 = {1{`RANDOM}};
  valid_934 = _RAND_935[0:0];
  _RAND_936 = {1{`RANDOM}};
  valid_935 = _RAND_936[0:0];
  _RAND_937 = {1{`RANDOM}};
  valid_936 = _RAND_937[0:0];
  _RAND_938 = {1{`RANDOM}};
  valid_937 = _RAND_938[0:0];
  _RAND_939 = {1{`RANDOM}};
  valid_938 = _RAND_939[0:0];
  _RAND_940 = {1{`RANDOM}};
  valid_939 = _RAND_940[0:0];
  _RAND_941 = {1{`RANDOM}};
  valid_940 = _RAND_941[0:0];
  _RAND_942 = {1{`RANDOM}};
  valid_941 = _RAND_942[0:0];
  _RAND_943 = {1{`RANDOM}};
  valid_942 = _RAND_943[0:0];
  _RAND_944 = {1{`RANDOM}};
  valid_943 = _RAND_944[0:0];
  _RAND_945 = {1{`RANDOM}};
  valid_944 = _RAND_945[0:0];
  _RAND_946 = {1{`RANDOM}};
  valid_945 = _RAND_946[0:0];
  _RAND_947 = {1{`RANDOM}};
  valid_946 = _RAND_947[0:0];
  _RAND_948 = {1{`RANDOM}};
  valid_947 = _RAND_948[0:0];
  _RAND_949 = {1{`RANDOM}};
  valid_948 = _RAND_949[0:0];
  _RAND_950 = {1{`RANDOM}};
  valid_949 = _RAND_950[0:0];
  _RAND_951 = {1{`RANDOM}};
  valid_950 = _RAND_951[0:0];
  _RAND_952 = {1{`RANDOM}};
  valid_951 = _RAND_952[0:0];
  _RAND_953 = {1{`RANDOM}};
  valid_952 = _RAND_953[0:0];
  _RAND_954 = {1{`RANDOM}};
  valid_953 = _RAND_954[0:0];
  _RAND_955 = {1{`RANDOM}};
  valid_954 = _RAND_955[0:0];
  _RAND_956 = {1{`RANDOM}};
  valid_955 = _RAND_956[0:0];
  _RAND_957 = {1{`RANDOM}};
  valid_956 = _RAND_957[0:0];
  _RAND_958 = {1{`RANDOM}};
  valid_957 = _RAND_958[0:0];
  _RAND_959 = {1{`RANDOM}};
  valid_958 = _RAND_959[0:0];
  _RAND_960 = {1{`RANDOM}};
  valid_959 = _RAND_960[0:0];
  _RAND_961 = {1{`RANDOM}};
  valid_960 = _RAND_961[0:0];
  _RAND_962 = {1{`RANDOM}};
  valid_961 = _RAND_962[0:0];
  _RAND_963 = {1{`RANDOM}};
  valid_962 = _RAND_963[0:0];
  _RAND_964 = {1{`RANDOM}};
  valid_963 = _RAND_964[0:0];
  _RAND_965 = {1{`RANDOM}};
  valid_964 = _RAND_965[0:0];
  _RAND_966 = {1{`RANDOM}};
  valid_965 = _RAND_966[0:0];
  _RAND_967 = {1{`RANDOM}};
  valid_966 = _RAND_967[0:0];
  _RAND_968 = {1{`RANDOM}};
  valid_967 = _RAND_968[0:0];
  _RAND_969 = {1{`RANDOM}};
  valid_968 = _RAND_969[0:0];
  _RAND_970 = {1{`RANDOM}};
  valid_969 = _RAND_970[0:0];
  _RAND_971 = {1{`RANDOM}};
  valid_970 = _RAND_971[0:0];
  _RAND_972 = {1{`RANDOM}};
  valid_971 = _RAND_972[0:0];
  _RAND_973 = {1{`RANDOM}};
  valid_972 = _RAND_973[0:0];
  _RAND_974 = {1{`RANDOM}};
  valid_973 = _RAND_974[0:0];
  _RAND_975 = {1{`RANDOM}};
  valid_974 = _RAND_975[0:0];
  _RAND_976 = {1{`RANDOM}};
  valid_975 = _RAND_976[0:0];
  _RAND_977 = {1{`RANDOM}};
  valid_976 = _RAND_977[0:0];
  _RAND_978 = {1{`RANDOM}};
  valid_977 = _RAND_978[0:0];
  _RAND_979 = {1{`RANDOM}};
  valid_978 = _RAND_979[0:0];
  _RAND_980 = {1{`RANDOM}};
  valid_979 = _RAND_980[0:0];
  _RAND_981 = {1{`RANDOM}};
  valid_980 = _RAND_981[0:0];
  _RAND_982 = {1{`RANDOM}};
  valid_981 = _RAND_982[0:0];
  _RAND_983 = {1{`RANDOM}};
  valid_982 = _RAND_983[0:0];
  _RAND_984 = {1{`RANDOM}};
  valid_983 = _RAND_984[0:0];
  _RAND_985 = {1{`RANDOM}};
  valid_984 = _RAND_985[0:0];
  _RAND_986 = {1{`RANDOM}};
  valid_985 = _RAND_986[0:0];
  _RAND_987 = {1{`RANDOM}};
  valid_986 = _RAND_987[0:0];
  _RAND_988 = {1{`RANDOM}};
  valid_987 = _RAND_988[0:0];
  _RAND_989 = {1{`RANDOM}};
  valid_988 = _RAND_989[0:0];
  _RAND_990 = {1{`RANDOM}};
  valid_989 = _RAND_990[0:0];
  _RAND_991 = {1{`RANDOM}};
  valid_990 = _RAND_991[0:0];
  _RAND_992 = {1{`RANDOM}};
  valid_991 = _RAND_992[0:0];
  _RAND_993 = {1{`RANDOM}};
  valid_992 = _RAND_993[0:0];
  _RAND_994 = {1{`RANDOM}};
  valid_993 = _RAND_994[0:0];
  _RAND_995 = {1{`RANDOM}};
  valid_994 = _RAND_995[0:0];
  _RAND_996 = {1{`RANDOM}};
  valid_995 = _RAND_996[0:0];
  _RAND_997 = {1{`RANDOM}};
  valid_996 = _RAND_997[0:0];
  _RAND_998 = {1{`RANDOM}};
  valid_997 = _RAND_998[0:0];
  _RAND_999 = {1{`RANDOM}};
  valid_998 = _RAND_999[0:0];
  _RAND_1000 = {1{`RANDOM}};
  valid_999 = _RAND_1000[0:0];
  _RAND_1001 = {1{`RANDOM}};
  valid_1000 = _RAND_1001[0:0];
  _RAND_1002 = {1{`RANDOM}};
  valid_1001 = _RAND_1002[0:0];
  _RAND_1003 = {1{`RANDOM}};
  valid_1002 = _RAND_1003[0:0];
  _RAND_1004 = {1{`RANDOM}};
  valid_1003 = _RAND_1004[0:0];
  _RAND_1005 = {1{`RANDOM}};
  valid_1004 = _RAND_1005[0:0];
  _RAND_1006 = {1{`RANDOM}};
  valid_1005 = _RAND_1006[0:0];
  _RAND_1007 = {1{`RANDOM}};
  valid_1006 = _RAND_1007[0:0];
  _RAND_1008 = {1{`RANDOM}};
  valid_1007 = _RAND_1008[0:0];
  _RAND_1009 = {1{`RANDOM}};
  valid_1008 = _RAND_1009[0:0];
  _RAND_1010 = {1{`RANDOM}};
  valid_1009 = _RAND_1010[0:0];
  _RAND_1011 = {1{`RANDOM}};
  valid_1010 = _RAND_1011[0:0];
  _RAND_1012 = {1{`RANDOM}};
  valid_1011 = _RAND_1012[0:0];
  _RAND_1013 = {1{`RANDOM}};
  valid_1012 = _RAND_1013[0:0];
  _RAND_1014 = {1{`RANDOM}};
  valid_1013 = _RAND_1014[0:0];
  _RAND_1015 = {1{`RANDOM}};
  valid_1014 = _RAND_1015[0:0];
  _RAND_1016 = {1{`RANDOM}};
  valid_1015 = _RAND_1016[0:0];
  _RAND_1017 = {1{`RANDOM}};
  valid_1016 = _RAND_1017[0:0];
  _RAND_1018 = {1{`RANDOM}};
  valid_1017 = _RAND_1018[0:0];
  _RAND_1019 = {1{`RANDOM}};
  valid_1018 = _RAND_1019[0:0];
  _RAND_1020 = {1{`RANDOM}};
  valid_1019 = _RAND_1020[0:0];
  _RAND_1021 = {1{`RANDOM}};
  valid_1020 = _RAND_1021[0:0];
  _RAND_1022 = {1{`RANDOM}};
  valid_1021 = _RAND_1022[0:0];
  _RAND_1023 = {1{`RANDOM}};
  valid_1022 = _RAND_1023[0:0];
  _RAND_1024 = {1{`RANDOM}};
  valid_1023 = _RAND_1024[0:0];
  _RAND_1025 = {1{`RANDOM}};
  state = _RAND_1025[2:0];
  _RAND_1026 = {1{`RANDOM}};
  array_out_REG = _RAND_1026[0:0];
  _RAND_1027 = {9{`RANDOM}};
  array_out_r = _RAND_1027[272:0];
  _RAND_1028 = {1{`RANDOM}};
  array_data_REG = _RAND_1028[0:0];
  _RAND_1029 = {2{`RANDOM}};
  array_data_r = _RAND_1029[63:0];
  _RAND_1030 = {8{`RANDOM}};
  wdata = _RAND_1030[255:0];
  _RAND_1031 = {1{`RANDOM}};
  source = _RAND_1031[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DCache(
  input          clock,
  input          reset,
  input          auto_out_a_ready,
  output         auto_out_a_valid,
  output [1:0]   auto_out_a_bits_source,
  output [31:0]  auto_out_a_bits_address,
  output         auto_out_b_ready,
  input          auto_out_b_valid,
  input  [2:0]   auto_out_b_bits_size,
  input  [1:0]   auto_out_b_bits_source,
  input  [31:0]  auto_out_b_bits_address,
  input          auto_out_c_ready,
  output         auto_out_c_valid,
  output [2:0]   auto_out_c_bits_opcode,
  output [2:0]   auto_out_c_bits_param,
  output [2:0]   auto_out_c_bits_size,
  output [1:0]   auto_out_c_bits_source,
  output [31:0]  auto_out_c_bits_address,
  output [255:0] auto_out_c_bits_data,
  output         auto_out_d_ready,
  input          auto_out_d_valid,
  input  [5:0]   auto_out_d_bits_sink,
  input  [255:0] auto_out_d_bits_data,
  input          auto_out_e_ready,
  output         auto_out_e_valid,
  output [5:0]   auto_out_e_bits_sink,
  output         io_cache_req_ready,
  input          io_cache_req_valid,
  input  [38:0]  io_cache_req_bits_addr,
  input  [63:0]  io_cache_req_bits_wdata,
  input  [7:0]   io_cache_req_bits_wmask,
  input          io_cache_req_bits_wen,
  input  [1:0]   io_cache_req_bits_len,
  input          io_cache_req_bits_lrsc,
  input  [4:0]   io_cache_req_bits_amo,
  input          io_cache_resp_ready,
  output         io_cache_resp_valid,
  output [63:0]  io_cache_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [255:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [31:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [31:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
  reg [31:0] _RAND_1034;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
  reg [31:0] _RAND_1038;
  reg [31:0] _RAND_1039;
  reg [31:0] _RAND_1040;
  reg [287:0] _RAND_1041;
  reg [31:0] _RAND_1042;
  reg [31:0] _RAND_1043;
  reg [31:0] _RAND_1044;
  reg [287:0] _RAND_1045;
  reg [31:0] _RAND_1046;
  reg [31:0] _RAND_1047;
`endif // RANDOMIZE_REG_INIT
  wire  array_clock; // @[DCache.scala 55:21]
  wire  array_io_en; // @[DCache.scala 55:21]
  wire [9:0] array_io_addr; // @[DCache.scala 55:21]
  wire [272:0] array_io_wdata; // @[DCache.scala 55:21]
  wire  array_io_wen; // @[DCache.scala 55:21]
  wire [272:0] array_io_rdata; // @[DCache.scala 55:21]
  reg  probing; // @[Utils.scala 36:20]
  wire  _x1_b_ready_T = ~probing; // @[DCache.scala 258:17]
  reg  lrsc_reserved; // @[DCache.scala 127:30]
  wire  _x1_b_ready_T_1 = ~lrsc_reserved; // @[DCache.scala 258:30]
  reg [4:0] lrsc_counter; // @[DCache.scala 129:30]
  wire  lrsc_backoff = lrsc_counter[4]; // @[DCache.scala 130:35]
  wire  tl_b_ready = ~probing & (~lrsc_reserved | lrsc_backoff); // @[DCache.scala 258:26]
  wire  _tl_b_bits_r_T = tl_b_ready & auto_out_b_valid; // @[Decoupled.scala 51:35]
  reg [2:0] tl_b_bits_r_size; // @[Reg.scala 35:20]
  reg [1:0] tl_b_bits_r_source; // @[Reg.scala 35:20]
  reg [31:0] tl_b_bits_r_address; // @[Reg.scala 35:20]
  wire [31:0] _GEN_4 = _tl_b_bits_r_T ? auto_out_b_bits_address : tl_b_bits_r_address; // @[Reg.scala 36:18 35:20 36:22]
  reg [2:0] state; // @[DCache.scala 60:118]
  wire  tl_d_ready = state == 3'h3 | state == 3'h5; // @[DCache.scala 261:43]
  wire  _tl_d_bits_r_T = tl_d_ready & auto_out_d_valid; // @[Decoupled.scala 51:35]
  reg [5:0] tl_d_bits_r_sink; // @[Reg.scala 35:20]
  reg [255:0] tl_d_bits_r_data; // @[Reg.scala 35:20]
  wire  _req_r_T = io_cache_req_ready & io_cache_req_valid; // @[Decoupled.scala 51:35]
  reg [38:0] req_r_addr; // @[Reg.scala 35:20]
  reg [63:0] req_r_wdata; // @[Reg.scala 35:20]
  reg [7:0] req_r_wmask; // @[Reg.scala 35:20]
  reg  req_r_wen; // @[Reg.scala 35:20]
  reg [1:0] req_r_len; // @[Reg.scala 35:20]
  reg  req_r_lrsc; // @[Reg.scala 35:20]
  reg [4:0] req_r_amo; // @[Reg.scala 35:20]
  wire [38:0] _GEN_16 = _req_r_T ? io_cache_req_bits_addr : req_r_addr; // @[Reg.scala 36:18 35:20 36:22]
  reg  valid_0; // @[DCache.scala 56:22]
  reg  valid_1; // @[DCache.scala 56:22]
  reg  valid_2; // @[DCache.scala 56:22]
  reg  valid_3; // @[DCache.scala 56:22]
  reg  valid_4; // @[DCache.scala 56:22]
  reg  valid_5; // @[DCache.scala 56:22]
  reg  valid_6; // @[DCache.scala 56:22]
  reg  valid_7; // @[DCache.scala 56:22]
  reg  valid_8; // @[DCache.scala 56:22]
  reg  valid_9; // @[DCache.scala 56:22]
  reg  valid_10; // @[DCache.scala 56:22]
  reg  valid_11; // @[DCache.scala 56:22]
  reg  valid_12; // @[DCache.scala 56:22]
  reg  valid_13; // @[DCache.scala 56:22]
  reg  valid_14; // @[DCache.scala 56:22]
  reg  valid_15; // @[DCache.scala 56:22]
  reg  valid_16; // @[DCache.scala 56:22]
  reg  valid_17; // @[DCache.scala 56:22]
  reg  valid_18; // @[DCache.scala 56:22]
  reg  valid_19; // @[DCache.scala 56:22]
  reg  valid_20; // @[DCache.scala 56:22]
  reg  valid_21; // @[DCache.scala 56:22]
  reg  valid_22; // @[DCache.scala 56:22]
  reg  valid_23; // @[DCache.scala 56:22]
  reg  valid_24; // @[DCache.scala 56:22]
  reg  valid_25; // @[DCache.scala 56:22]
  reg  valid_26; // @[DCache.scala 56:22]
  reg  valid_27; // @[DCache.scala 56:22]
  reg  valid_28; // @[DCache.scala 56:22]
  reg  valid_29; // @[DCache.scala 56:22]
  reg  valid_30; // @[DCache.scala 56:22]
  reg  valid_31; // @[DCache.scala 56:22]
  reg  valid_32; // @[DCache.scala 56:22]
  reg  valid_33; // @[DCache.scala 56:22]
  reg  valid_34; // @[DCache.scala 56:22]
  reg  valid_35; // @[DCache.scala 56:22]
  reg  valid_36; // @[DCache.scala 56:22]
  reg  valid_37; // @[DCache.scala 56:22]
  reg  valid_38; // @[DCache.scala 56:22]
  reg  valid_39; // @[DCache.scala 56:22]
  reg  valid_40; // @[DCache.scala 56:22]
  reg  valid_41; // @[DCache.scala 56:22]
  reg  valid_42; // @[DCache.scala 56:22]
  reg  valid_43; // @[DCache.scala 56:22]
  reg  valid_44; // @[DCache.scala 56:22]
  reg  valid_45; // @[DCache.scala 56:22]
  reg  valid_46; // @[DCache.scala 56:22]
  reg  valid_47; // @[DCache.scala 56:22]
  reg  valid_48; // @[DCache.scala 56:22]
  reg  valid_49; // @[DCache.scala 56:22]
  reg  valid_50; // @[DCache.scala 56:22]
  reg  valid_51; // @[DCache.scala 56:22]
  reg  valid_52; // @[DCache.scala 56:22]
  reg  valid_53; // @[DCache.scala 56:22]
  reg  valid_54; // @[DCache.scala 56:22]
  reg  valid_55; // @[DCache.scala 56:22]
  reg  valid_56; // @[DCache.scala 56:22]
  reg  valid_57; // @[DCache.scala 56:22]
  reg  valid_58; // @[DCache.scala 56:22]
  reg  valid_59; // @[DCache.scala 56:22]
  reg  valid_60; // @[DCache.scala 56:22]
  reg  valid_61; // @[DCache.scala 56:22]
  reg  valid_62; // @[DCache.scala 56:22]
  reg  valid_63; // @[DCache.scala 56:22]
  reg  valid_64; // @[DCache.scala 56:22]
  reg  valid_65; // @[DCache.scala 56:22]
  reg  valid_66; // @[DCache.scala 56:22]
  reg  valid_67; // @[DCache.scala 56:22]
  reg  valid_68; // @[DCache.scala 56:22]
  reg  valid_69; // @[DCache.scala 56:22]
  reg  valid_70; // @[DCache.scala 56:22]
  reg  valid_71; // @[DCache.scala 56:22]
  reg  valid_72; // @[DCache.scala 56:22]
  reg  valid_73; // @[DCache.scala 56:22]
  reg  valid_74; // @[DCache.scala 56:22]
  reg  valid_75; // @[DCache.scala 56:22]
  reg  valid_76; // @[DCache.scala 56:22]
  reg  valid_77; // @[DCache.scala 56:22]
  reg  valid_78; // @[DCache.scala 56:22]
  reg  valid_79; // @[DCache.scala 56:22]
  reg  valid_80; // @[DCache.scala 56:22]
  reg  valid_81; // @[DCache.scala 56:22]
  reg  valid_82; // @[DCache.scala 56:22]
  reg  valid_83; // @[DCache.scala 56:22]
  reg  valid_84; // @[DCache.scala 56:22]
  reg  valid_85; // @[DCache.scala 56:22]
  reg  valid_86; // @[DCache.scala 56:22]
  reg  valid_87; // @[DCache.scala 56:22]
  reg  valid_88; // @[DCache.scala 56:22]
  reg  valid_89; // @[DCache.scala 56:22]
  reg  valid_90; // @[DCache.scala 56:22]
  reg  valid_91; // @[DCache.scala 56:22]
  reg  valid_92; // @[DCache.scala 56:22]
  reg  valid_93; // @[DCache.scala 56:22]
  reg  valid_94; // @[DCache.scala 56:22]
  reg  valid_95; // @[DCache.scala 56:22]
  reg  valid_96; // @[DCache.scala 56:22]
  reg  valid_97; // @[DCache.scala 56:22]
  reg  valid_98; // @[DCache.scala 56:22]
  reg  valid_99; // @[DCache.scala 56:22]
  reg  valid_100; // @[DCache.scala 56:22]
  reg  valid_101; // @[DCache.scala 56:22]
  reg  valid_102; // @[DCache.scala 56:22]
  reg  valid_103; // @[DCache.scala 56:22]
  reg  valid_104; // @[DCache.scala 56:22]
  reg  valid_105; // @[DCache.scala 56:22]
  reg  valid_106; // @[DCache.scala 56:22]
  reg  valid_107; // @[DCache.scala 56:22]
  reg  valid_108; // @[DCache.scala 56:22]
  reg  valid_109; // @[DCache.scala 56:22]
  reg  valid_110; // @[DCache.scala 56:22]
  reg  valid_111; // @[DCache.scala 56:22]
  reg  valid_112; // @[DCache.scala 56:22]
  reg  valid_113; // @[DCache.scala 56:22]
  reg  valid_114; // @[DCache.scala 56:22]
  reg  valid_115; // @[DCache.scala 56:22]
  reg  valid_116; // @[DCache.scala 56:22]
  reg  valid_117; // @[DCache.scala 56:22]
  reg  valid_118; // @[DCache.scala 56:22]
  reg  valid_119; // @[DCache.scala 56:22]
  reg  valid_120; // @[DCache.scala 56:22]
  reg  valid_121; // @[DCache.scala 56:22]
  reg  valid_122; // @[DCache.scala 56:22]
  reg  valid_123; // @[DCache.scala 56:22]
  reg  valid_124; // @[DCache.scala 56:22]
  reg  valid_125; // @[DCache.scala 56:22]
  reg  valid_126; // @[DCache.scala 56:22]
  reg  valid_127; // @[DCache.scala 56:22]
  reg  valid_128; // @[DCache.scala 56:22]
  reg  valid_129; // @[DCache.scala 56:22]
  reg  valid_130; // @[DCache.scala 56:22]
  reg  valid_131; // @[DCache.scala 56:22]
  reg  valid_132; // @[DCache.scala 56:22]
  reg  valid_133; // @[DCache.scala 56:22]
  reg  valid_134; // @[DCache.scala 56:22]
  reg  valid_135; // @[DCache.scala 56:22]
  reg  valid_136; // @[DCache.scala 56:22]
  reg  valid_137; // @[DCache.scala 56:22]
  reg  valid_138; // @[DCache.scala 56:22]
  reg  valid_139; // @[DCache.scala 56:22]
  reg  valid_140; // @[DCache.scala 56:22]
  reg  valid_141; // @[DCache.scala 56:22]
  reg  valid_142; // @[DCache.scala 56:22]
  reg  valid_143; // @[DCache.scala 56:22]
  reg  valid_144; // @[DCache.scala 56:22]
  reg  valid_145; // @[DCache.scala 56:22]
  reg  valid_146; // @[DCache.scala 56:22]
  reg  valid_147; // @[DCache.scala 56:22]
  reg  valid_148; // @[DCache.scala 56:22]
  reg  valid_149; // @[DCache.scala 56:22]
  reg  valid_150; // @[DCache.scala 56:22]
  reg  valid_151; // @[DCache.scala 56:22]
  reg  valid_152; // @[DCache.scala 56:22]
  reg  valid_153; // @[DCache.scala 56:22]
  reg  valid_154; // @[DCache.scala 56:22]
  reg  valid_155; // @[DCache.scala 56:22]
  reg  valid_156; // @[DCache.scala 56:22]
  reg  valid_157; // @[DCache.scala 56:22]
  reg  valid_158; // @[DCache.scala 56:22]
  reg  valid_159; // @[DCache.scala 56:22]
  reg  valid_160; // @[DCache.scala 56:22]
  reg  valid_161; // @[DCache.scala 56:22]
  reg  valid_162; // @[DCache.scala 56:22]
  reg  valid_163; // @[DCache.scala 56:22]
  reg  valid_164; // @[DCache.scala 56:22]
  reg  valid_165; // @[DCache.scala 56:22]
  reg  valid_166; // @[DCache.scala 56:22]
  reg  valid_167; // @[DCache.scala 56:22]
  reg  valid_168; // @[DCache.scala 56:22]
  reg  valid_169; // @[DCache.scala 56:22]
  reg  valid_170; // @[DCache.scala 56:22]
  reg  valid_171; // @[DCache.scala 56:22]
  reg  valid_172; // @[DCache.scala 56:22]
  reg  valid_173; // @[DCache.scala 56:22]
  reg  valid_174; // @[DCache.scala 56:22]
  reg  valid_175; // @[DCache.scala 56:22]
  reg  valid_176; // @[DCache.scala 56:22]
  reg  valid_177; // @[DCache.scala 56:22]
  reg  valid_178; // @[DCache.scala 56:22]
  reg  valid_179; // @[DCache.scala 56:22]
  reg  valid_180; // @[DCache.scala 56:22]
  reg  valid_181; // @[DCache.scala 56:22]
  reg  valid_182; // @[DCache.scala 56:22]
  reg  valid_183; // @[DCache.scala 56:22]
  reg  valid_184; // @[DCache.scala 56:22]
  reg  valid_185; // @[DCache.scala 56:22]
  reg  valid_186; // @[DCache.scala 56:22]
  reg  valid_187; // @[DCache.scala 56:22]
  reg  valid_188; // @[DCache.scala 56:22]
  reg  valid_189; // @[DCache.scala 56:22]
  reg  valid_190; // @[DCache.scala 56:22]
  reg  valid_191; // @[DCache.scala 56:22]
  reg  valid_192; // @[DCache.scala 56:22]
  reg  valid_193; // @[DCache.scala 56:22]
  reg  valid_194; // @[DCache.scala 56:22]
  reg  valid_195; // @[DCache.scala 56:22]
  reg  valid_196; // @[DCache.scala 56:22]
  reg  valid_197; // @[DCache.scala 56:22]
  reg  valid_198; // @[DCache.scala 56:22]
  reg  valid_199; // @[DCache.scala 56:22]
  reg  valid_200; // @[DCache.scala 56:22]
  reg  valid_201; // @[DCache.scala 56:22]
  reg  valid_202; // @[DCache.scala 56:22]
  reg  valid_203; // @[DCache.scala 56:22]
  reg  valid_204; // @[DCache.scala 56:22]
  reg  valid_205; // @[DCache.scala 56:22]
  reg  valid_206; // @[DCache.scala 56:22]
  reg  valid_207; // @[DCache.scala 56:22]
  reg  valid_208; // @[DCache.scala 56:22]
  reg  valid_209; // @[DCache.scala 56:22]
  reg  valid_210; // @[DCache.scala 56:22]
  reg  valid_211; // @[DCache.scala 56:22]
  reg  valid_212; // @[DCache.scala 56:22]
  reg  valid_213; // @[DCache.scala 56:22]
  reg  valid_214; // @[DCache.scala 56:22]
  reg  valid_215; // @[DCache.scala 56:22]
  reg  valid_216; // @[DCache.scala 56:22]
  reg  valid_217; // @[DCache.scala 56:22]
  reg  valid_218; // @[DCache.scala 56:22]
  reg  valid_219; // @[DCache.scala 56:22]
  reg  valid_220; // @[DCache.scala 56:22]
  reg  valid_221; // @[DCache.scala 56:22]
  reg  valid_222; // @[DCache.scala 56:22]
  reg  valid_223; // @[DCache.scala 56:22]
  reg  valid_224; // @[DCache.scala 56:22]
  reg  valid_225; // @[DCache.scala 56:22]
  reg  valid_226; // @[DCache.scala 56:22]
  reg  valid_227; // @[DCache.scala 56:22]
  reg  valid_228; // @[DCache.scala 56:22]
  reg  valid_229; // @[DCache.scala 56:22]
  reg  valid_230; // @[DCache.scala 56:22]
  reg  valid_231; // @[DCache.scala 56:22]
  reg  valid_232; // @[DCache.scala 56:22]
  reg  valid_233; // @[DCache.scala 56:22]
  reg  valid_234; // @[DCache.scala 56:22]
  reg  valid_235; // @[DCache.scala 56:22]
  reg  valid_236; // @[DCache.scala 56:22]
  reg  valid_237; // @[DCache.scala 56:22]
  reg  valid_238; // @[DCache.scala 56:22]
  reg  valid_239; // @[DCache.scala 56:22]
  reg  valid_240; // @[DCache.scala 56:22]
  reg  valid_241; // @[DCache.scala 56:22]
  reg  valid_242; // @[DCache.scala 56:22]
  reg  valid_243; // @[DCache.scala 56:22]
  reg  valid_244; // @[DCache.scala 56:22]
  reg  valid_245; // @[DCache.scala 56:22]
  reg  valid_246; // @[DCache.scala 56:22]
  reg  valid_247; // @[DCache.scala 56:22]
  reg  valid_248; // @[DCache.scala 56:22]
  reg  valid_249; // @[DCache.scala 56:22]
  reg  valid_250; // @[DCache.scala 56:22]
  reg  valid_251; // @[DCache.scala 56:22]
  reg  valid_252; // @[DCache.scala 56:22]
  reg  valid_253; // @[DCache.scala 56:22]
  reg  valid_254; // @[DCache.scala 56:22]
  reg  valid_255; // @[DCache.scala 56:22]
  reg  valid_256; // @[DCache.scala 56:22]
  reg  valid_257; // @[DCache.scala 56:22]
  reg  valid_258; // @[DCache.scala 56:22]
  reg  valid_259; // @[DCache.scala 56:22]
  reg  valid_260; // @[DCache.scala 56:22]
  reg  valid_261; // @[DCache.scala 56:22]
  reg  valid_262; // @[DCache.scala 56:22]
  reg  valid_263; // @[DCache.scala 56:22]
  reg  valid_264; // @[DCache.scala 56:22]
  reg  valid_265; // @[DCache.scala 56:22]
  reg  valid_266; // @[DCache.scala 56:22]
  reg  valid_267; // @[DCache.scala 56:22]
  reg  valid_268; // @[DCache.scala 56:22]
  reg  valid_269; // @[DCache.scala 56:22]
  reg  valid_270; // @[DCache.scala 56:22]
  reg  valid_271; // @[DCache.scala 56:22]
  reg  valid_272; // @[DCache.scala 56:22]
  reg  valid_273; // @[DCache.scala 56:22]
  reg  valid_274; // @[DCache.scala 56:22]
  reg  valid_275; // @[DCache.scala 56:22]
  reg  valid_276; // @[DCache.scala 56:22]
  reg  valid_277; // @[DCache.scala 56:22]
  reg  valid_278; // @[DCache.scala 56:22]
  reg  valid_279; // @[DCache.scala 56:22]
  reg  valid_280; // @[DCache.scala 56:22]
  reg  valid_281; // @[DCache.scala 56:22]
  reg  valid_282; // @[DCache.scala 56:22]
  reg  valid_283; // @[DCache.scala 56:22]
  reg  valid_284; // @[DCache.scala 56:22]
  reg  valid_285; // @[DCache.scala 56:22]
  reg  valid_286; // @[DCache.scala 56:22]
  reg  valid_287; // @[DCache.scala 56:22]
  reg  valid_288; // @[DCache.scala 56:22]
  reg  valid_289; // @[DCache.scala 56:22]
  reg  valid_290; // @[DCache.scala 56:22]
  reg  valid_291; // @[DCache.scala 56:22]
  reg  valid_292; // @[DCache.scala 56:22]
  reg  valid_293; // @[DCache.scala 56:22]
  reg  valid_294; // @[DCache.scala 56:22]
  reg  valid_295; // @[DCache.scala 56:22]
  reg  valid_296; // @[DCache.scala 56:22]
  reg  valid_297; // @[DCache.scala 56:22]
  reg  valid_298; // @[DCache.scala 56:22]
  reg  valid_299; // @[DCache.scala 56:22]
  reg  valid_300; // @[DCache.scala 56:22]
  reg  valid_301; // @[DCache.scala 56:22]
  reg  valid_302; // @[DCache.scala 56:22]
  reg  valid_303; // @[DCache.scala 56:22]
  reg  valid_304; // @[DCache.scala 56:22]
  reg  valid_305; // @[DCache.scala 56:22]
  reg  valid_306; // @[DCache.scala 56:22]
  reg  valid_307; // @[DCache.scala 56:22]
  reg  valid_308; // @[DCache.scala 56:22]
  reg  valid_309; // @[DCache.scala 56:22]
  reg  valid_310; // @[DCache.scala 56:22]
  reg  valid_311; // @[DCache.scala 56:22]
  reg  valid_312; // @[DCache.scala 56:22]
  reg  valid_313; // @[DCache.scala 56:22]
  reg  valid_314; // @[DCache.scala 56:22]
  reg  valid_315; // @[DCache.scala 56:22]
  reg  valid_316; // @[DCache.scala 56:22]
  reg  valid_317; // @[DCache.scala 56:22]
  reg  valid_318; // @[DCache.scala 56:22]
  reg  valid_319; // @[DCache.scala 56:22]
  reg  valid_320; // @[DCache.scala 56:22]
  reg  valid_321; // @[DCache.scala 56:22]
  reg  valid_322; // @[DCache.scala 56:22]
  reg  valid_323; // @[DCache.scala 56:22]
  reg  valid_324; // @[DCache.scala 56:22]
  reg  valid_325; // @[DCache.scala 56:22]
  reg  valid_326; // @[DCache.scala 56:22]
  reg  valid_327; // @[DCache.scala 56:22]
  reg  valid_328; // @[DCache.scala 56:22]
  reg  valid_329; // @[DCache.scala 56:22]
  reg  valid_330; // @[DCache.scala 56:22]
  reg  valid_331; // @[DCache.scala 56:22]
  reg  valid_332; // @[DCache.scala 56:22]
  reg  valid_333; // @[DCache.scala 56:22]
  reg  valid_334; // @[DCache.scala 56:22]
  reg  valid_335; // @[DCache.scala 56:22]
  reg  valid_336; // @[DCache.scala 56:22]
  reg  valid_337; // @[DCache.scala 56:22]
  reg  valid_338; // @[DCache.scala 56:22]
  reg  valid_339; // @[DCache.scala 56:22]
  reg  valid_340; // @[DCache.scala 56:22]
  reg  valid_341; // @[DCache.scala 56:22]
  reg  valid_342; // @[DCache.scala 56:22]
  reg  valid_343; // @[DCache.scala 56:22]
  reg  valid_344; // @[DCache.scala 56:22]
  reg  valid_345; // @[DCache.scala 56:22]
  reg  valid_346; // @[DCache.scala 56:22]
  reg  valid_347; // @[DCache.scala 56:22]
  reg  valid_348; // @[DCache.scala 56:22]
  reg  valid_349; // @[DCache.scala 56:22]
  reg  valid_350; // @[DCache.scala 56:22]
  reg  valid_351; // @[DCache.scala 56:22]
  reg  valid_352; // @[DCache.scala 56:22]
  reg  valid_353; // @[DCache.scala 56:22]
  reg  valid_354; // @[DCache.scala 56:22]
  reg  valid_355; // @[DCache.scala 56:22]
  reg  valid_356; // @[DCache.scala 56:22]
  reg  valid_357; // @[DCache.scala 56:22]
  reg  valid_358; // @[DCache.scala 56:22]
  reg  valid_359; // @[DCache.scala 56:22]
  reg  valid_360; // @[DCache.scala 56:22]
  reg  valid_361; // @[DCache.scala 56:22]
  reg  valid_362; // @[DCache.scala 56:22]
  reg  valid_363; // @[DCache.scala 56:22]
  reg  valid_364; // @[DCache.scala 56:22]
  reg  valid_365; // @[DCache.scala 56:22]
  reg  valid_366; // @[DCache.scala 56:22]
  reg  valid_367; // @[DCache.scala 56:22]
  reg  valid_368; // @[DCache.scala 56:22]
  reg  valid_369; // @[DCache.scala 56:22]
  reg  valid_370; // @[DCache.scala 56:22]
  reg  valid_371; // @[DCache.scala 56:22]
  reg  valid_372; // @[DCache.scala 56:22]
  reg  valid_373; // @[DCache.scala 56:22]
  reg  valid_374; // @[DCache.scala 56:22]
  reg  valid_375; // @[DCache.scala 56:22]
  reg  valid_376; // @[DCache.scala 56:22]
  reg  valid_377; // @[DCache.scala 56:22]
  reg  valid_378; // @[DCache.scala 56:22]
  reg  valid_379; // @[DCache.scala 56:22]
  reg  valid_380; // @[DCache.scala 56:22]
  reg  valid_381; // @[DCache.scala 56:22]
  reg  valid_382; // @[DCache.scala 56:22]
  reg  valid_383; // @[DCache.scala 56:22]
  reg  valid_384; // @[DCache.scala 56:22]
  reg  valid_385; // @[DCache.scala 56:22]
  reg  valid_386; // @[DCache.scala 56:22]
  reg  valid_387; // @[DCache.scala 56:22]
  reg  valid_388; // @[DCache.scala 56:22]
  reg  valid_389; // @[DCache.scala 56:22]
  reg  valid_390; // @[DCache.scala 56:22]
  reg  valid_391; // @[DCache.scala 56:22]
  reg  valid_392; // @[DCache.scala 56:22]
  reg  valid_393; // @[DCache.scala 56:22]
  reg  valid_394; // @[DCache.scala 56:22]
  reg  valid_395; // @[DCache.scala 56:22]
  reg  valid_396; // @[DCache.scala 56:22]
  reg  valid_397; // @[DCache.scala 56:22]
  reg  valid_398; // @[DCache.scala 56:22]
  reg  valid_399; // @[DCache.scala 56:22]
  reg  valid_400; // @[DCache.scala 56:22]
  reg  valid_401; // @[DCache.scala 56:22]
  reg  valid_402; // @[DCache.scala 56:22]
  reg  valid_403; // @[DCache.scala 56:22]
  reg  valid_404; // @[DCache.scala 56:22]
  reg  valid_405; // @[DCache.scala 56:22]
  reg  valid_406; // @[DCache.scala 56:22]
  reg  valid_407; // @[DCache.scala 56:22]
  reg  valid_408; // @[DCache.scala 56:22]
  reg  valid_409; // @[DCache.scala 56:22]
  reg  valid_410; // @[DCache.scala 56:22]
  reg  valid_411; // @[DCache.scala 56:22]
  reg  valid_412; // @[DCache.scala 56:22]
  reg  valid_413; // @[DCache.scala 56:22]
  reg  valid_414; // @[DCache.scala 56:22]
  reg  valid_415; // @[DCache.scala 56:22]
  reg  valid_416; // @[DCache.scala 56:22]
  reg  valid_417; // @[DCache.scala 56:22]
  reg  valid_418; // @[DCache.scala 56:22]
  reg  valid_419; // @[DCache.scala 56:22]
  reg  valid_420; // @[DCache.scala 56:22]
  reg  valid_421; // @[DCache.scala 56:22]
  reg  valid_422; // @[DCache.scala 56:22]
  reg  valid_423; // @[DCache.scala 56:22]
  reg  valid_424; // @[DCache.scala 56:22]
  reg  valid_425; // @[DCache.scala 56:22]
  reg  valid_426; // @[DCache.scala 56:22]
  reg  valid_427; // @[DCache.scala 56:22]
  reg  valid_428; // @[DCache.scala 56:22]
  reg  valid_429; // @[DCache.scala 56:22]
  reg  valid_430; // @[DCache.scala 56:22]
  reg  valid_431; // @[DCache.scala 56:22]
  reg  valid_432; // @[DCache.scala 56:22]
  reg  valid_433; // @[DCache.scala 56:22]
  reg  valid_434; // @[DCache.scala 56:22]
  reg  valid_435; // @[DCache.scala 56:22]
  reg  valid_436; // @[DCache.scala 56:22]
  reg  valid_437; // @[DCache.scala 56:22]
  reg  valid_438; // @[DCache.scala 56:22]
  reg  valid_439; // @[DCache.scala 56:22]
  reg  valid_440; // @[DCache.scala 56:22]
  reg  valid_441; // @[DCache.scala 56:22]
  reg  valid_442; // @[DCache.scala 56:22]
  reg  valid_443; // @[DCache.scala 56:22]
  reg  valid_444; // @[DCache.scala 56:22]
  reg  valid_445; // @[DCache.scala 56:22]
  reg  valid_446; // @[DCache.scala 56:22]
  reg  valid_447; // @[DCache.scala 56:22]
  reg  valid_448; // @[DCache.scala 56:22]
  reg  valid_449; // @[DCache.scala 56:22]
  reg  valid_450; // @[DCache.scala 56:22]
  reg  valid_451; // @[DCache.scala 56:22]
  reg  valid_452; // @[DCache.scala 56:22]
  reg  valid_453; // @[DCache.scala 56:22]
  reg  valid_454; // @[DCache.scala 56:22]
  reg  valid_455; // @[DCache.scala 56:22]
  reg  valid_456; // @[DCache.scala 56:22]
  reg  valid_457; // @[DCache.scala 56:22]
  reg  valid_458; // @[DCache.scala 56:22]
  reg  valid_459; // @[DCache.scala 56:22]
  reg  valid_460; // @[DCache.scala 56:22]
  reg  valid_461; // @[DCache.scala 56:22]
  reg  valid_462; // @[DCache.scala 56:22]
  reg  valid_463; // @[DCache.scala 56:22]
  reg  valid_464; // @[DCache.scala 56:22]
  reg  valid_465; // @[DCache.scala 56:22]
  reg  valid_466; // @[DCache.scala 56:22]
  reg  valid_467; // @[DCache.scala 56:22]
  reg  valid_468; // @[DCache.scala 56:22]
  reg  valid_469; // @[DCache.scala 56:22]
  reg  valid_470; // @[DCache.scala 56:22]
  reg  valid_471; // @[DCache.scala 56:22]
  reg  valid_472; // @[DCache.scala 56:22]
  reg  valid_473; // @[DCache.scala 56:22]
  reg  valid_474; // @[DCache.scala 56:22]
  reg  valid_475; // @[DCache.scala 56:22]
  reg  valid_476; // @[DCache.scala 56:22]
  reg  valid_477; // @[DCache.scala 56:22]
  reg  valid_478; // @[DCache.scala 56:22]
  reg  valid_479; // @[DCache.scala 56:22]
  reg  valid_480; // @[DCache.scala 56:22]
  reg  valid_481; // @[DCache.scala 56:22]
  reg  valid_482; // @[DCache.scala 56:22]
  reg  valid_483; // @[DCache.scala 56:22]
  reg  valid_484; // @[DCache.scala 56:22]
  reg  valid_485; // @[DCache.scala 56:22]
  reg  valid_486; // @[DCache.scala 56:22]
  reg  valid_487; // @[DCache.scala 56:22]
  reg  valid_488; // @[DCache.scala 56:22]
  reg  valid_489; // @[DCache.scala 56:22]
  reg  valid_490; // @[DCache.scala 56:22]
  reg  valid_491; // @[DCache.scala 56:22]
  reg  valid_492; // @[DCache.scala 56:22]
  reg  valid_493; // @[DCache.scala 56:22]
  reg  valid_494; // @[DCache.scala 56:22]
  reg  valid_495; // @[DCache.scala 56:22]
  reg  valid_496; // @[DCache.scala 56:22]
  reg  valid_497; // @[DCache.scala 56:22]
  reg  valid_498; // @[DCache.scala 56:22]
  reg  valid_499; // @[DCache.scala 56:22]
  reg  valid_500; // @[DCache.scala 56:22]
  reg  valid_501; // @[DCache.scala 56:22]
  reg  valid_502; // @[DCache.scala 56:22]
  reg  valid_503; // @[DCache.scala 56:22]
  reg  valid_504; // @[DCache.scala 56:22]
  reg  valid_505; // @[DCache.scala 56:22]
  reg  valid_506; // @[DCache.scala 56:22]
  reg  valid_507; // @[DCache.scala 56:22]
  reg  valid_508; // @[DCache.scala 56:22]
  reg  valid_509; // @[DCache.scala 56:22]
  reg  valid_510; // @[DCache.scala 56:22]
  reg  valid_511; // @[DCache.scala 56:22]
  reg  valid_512; // @[DCache.scala 56:22]
  reg  valid_513; // @[DCache.scala 56:22]
  reg  valid_514; // @[DCache.scala 56:22]
  reg  valid_515; // @[DCache.scala 56:22]
  reg  valid_516; // @[DCache.scala 56:22]
  reg  valid_517; // @[DCache.scala 56:22]
  reg  valid_518; // @[DCache.scala 56:22]
  reg  valid_519; // @[DCache.scala 56:22]
  reg  valid_520; // @[DCache.scala 56:22]
  reg  valid_521; // @[DCache.scala 56:22]
  reg  valid_522; // @[DCache.scala 56:22]
  reg  valid_523; // @[DCache.scala 56:22]
  reg  valid_524; // @[DCache.scala 56:22]
  reg  valid_525; // @[DCache.scala 56:22]
  reg  valid_526; // @[DCache.scala 56:22]
  reg  valid_527; // @[DCache.scala 56:22]
  reg  valid_528; // @[DCache.scala 56:22]
  reg  valid_529; // @[DCache.scala 56:22]
  reg  valid_530; // @[DCache.scala 56:22]
  reg  valid_531; // @[DCache.scala 56:22]
  reg  valid_532; // @[DCache.scala 56:22]
  reg  valid_533; // @[DCache.scala 56:22]
  reg  valid_534; // @[DCache.scala 56:22]
  reg  valid_535; // @[DCache.scala 56:22]
  reg  valid_536; // @[DCache.scala 56:22]
  reg  valid_537; // @[DCache.scala 56:22]
  reg  valid_538; // @[DCache.scala 56:22]
  reg  valid_539; // @[DCache.scala 56:22]
  reg  valid_540; // @[DCache.scala 56:22]
  reg  valid_541; // @[DCache.scala 56:22]
  reg  valid_542; // @[DCache.scala 56:22]
  reg  valid_543; // @[DCache.scala 56:22]
  reg  valid_544; // @[DCache.scala 56:22]
  reg  valid_545; // @[DCache.scala 56:22]
  reg  valid_546; // @[DCache.scala 56:22]
  reg  valid_547; // @[DCache.scala 56:22]
  reg  valid_548; // @[DCache.scala 56:22]
  reg  valid_549; // @[DCache.scala 56:22]
  reg  valid_550; // @[DCache.scala 56:22]
  reg  valid_551; // @[DCache.scala 56:22]
  reg  valid_552; // @[DCache.scala 56:22]
  reg  valid_553; // @[DCache.scala 56:22]
  reg  valid_554; // @[DCache.scala 56:22]
  reg  valid_555; // @[DCache.scala 56:22]
  reg  valid_556; // @[DCache.scala 56:22]
  reg  valid_557; // @[DCache.scala 56:22]
  reg  valid_558; // @[DCache.scala 56:22]
  reg  valid_559; // @[DCache.scala 56:22]
  reg  valid_560; // @[DCache.scala 56:22]
  reg  valid_561; // @[DCache.scala 56:22]
  reg  valid_562; // @[DCache.scala 56:22]
  reg  valid_563; // @[DCache.scala 56:22]
  reg  valid_564; // @[DCache.scala 56:22]
  reg  valid_565; // @[DCache.scala 56:22]
  reg  valid_566; // @[DCache.scala 56:22]
  reg  valid_567; // @[DCache.scala 56:22]
  reg  valid_568; // @[DCache.scala 56:22]
  reg  valid_569; // @[DCache.scala 56:22]
  reg  valid_570; // @[DCache.scala 56:22]
  reg  valid_571; // @[DCache.scala 56:22]
  reg  valid_572; // @[DCache.scala 56:22]
  reg  valid_573; // @[DCache.scala 56:22]
  reg  valid_574; // @[DCache.scala 56:22]
  reg  valid_575; // @[DCache.scala 56:22]
  reg  valid_576; // @[DCache.scala 56:22]
  reg  valid_577; // @[DCache.scala 56:22]
  reg  valid_578; // @[DCache.scala 56:22]
  reg  valid_579; // @[DCache.scala 56:22]
  reg  valid_580; // @[DCache.scala 56:22]
  reg  valid_581; // @[DCache.scala 56:22]
  reg  valid_582; // @[DCache.scala 56:22]
  reg  valid_583; // @[DCache.scala 56:22]
  reg  valid_584; // @[DCache.scala 56:22]
  reg  valid_585; // @[DCache.scala 56:22]
  reg  valid_586; // @[DCache.scala 56:22]
  reg  valid_587; // @[DCache.scala 56:22]
  reg  valid_588; // @[DCache.scala 56:22]
  reg  valid_589; // @[DCache.scala 56:22]
  reg  valid_590; // @[DCache.scala 56:22]
  reg  valid_591; // @[DCache.scala 56:22]
  reg  valid_592; // @[DCache.scala 56:22]
  reg  valid_593; // @[DCache.scala 56:22]
  reg  valid_594; // @[DCache.scala 56:22]
  reg  valid_595; // @[DCache.scala 56:22]
  reg  valid_596; // @[DCache.scala 56:22]
  reg  valid_597; // @[DCache.scala 56:22]
  reg  valid_598; // @[DCache.scala 56:22]
  reg  valid_599; // @[DCache.scala 56:22]
  reg  valid_600; // @[DCache.scala 56:22]
  reg  valid_601; // @[DCache.scala 56:22]
  reg  valid_602; // @[DCache.scala 56:22]
  reg  valid_603; // @[DCache.scala 56:22]
  reg  valid_604; // @[DCache.scala 56:22]
  reg  valid_605; // @[DCache.scala 56:22]
  reg  valid_606; // @[DCache.scala 56:22]
  reg  valid_607; // @[DCache.scala 56:22]
  reg  valid_608; // @[DCache.scala 56:22]
  reg  valid_609; // @[DCache.scala 56:22]
  reg  valid_610; // @[DCache.scala 56:22]
  reg  valid_611; // @[DCache.scala 56:22]
  reg  valid_612; // @[DCache.scala 56:22]
  reg  valid_613; // @[DCache.scala 56:22]
  reg  valid_614; // @[DCache.scala 56:22]
  reg  valid_615; // @[DCache.scala 56:22]
  reg  valid_616; // @[DCache.scala 56:22]
  reg  valid_617; // @[DCache.scala 56:22]
  reg  valid_618; // @[DCache.scala 56:22]
  reg  valid_619; // @[DCache.scala 56:22]
  reg  valid_620; // @[DCache.scala 56:22]
  reg  valid_621; // @[DCache.scala 56:22]
  reg  valid_622; // @[DCache.scala 56:22]
  reg  valid_623; // @[DCache.scala 56:22]
  reg  valid_624; // @[DCache.scala 56:22]
  reg  valid_625; // @[DCache.scala 56:22]
  reg  valid_626; // @[DCache.scala 56:22]
  reg  valid_627; // @[DCache.scala 56:22]
  reg  valid_628; // @[DCache.scala 56:22]
  reg  valid_629; // @[DCache.scala 56:22]
  reg  valid_630; // @[DCache.scala 56:22]
  reg  valid_631; // @[DCache.scala 56:22]
  reg  valid_632; // @[DCache.scala 56:22]
  reg  valid_633; // @[DCache.scala 56:22]
  reg  valid_634; // @[DCache.scala 56:22]
  reg  valid_635; // @[DCache.scala 56:22]
  reg  valid_636; // @[DCache.scala 56:22]
  reg  valid_637; // @[DCache.scala 56:22]
  reg  valid_638; // @[DCache.scala 56:22]
  reg  valid_639; // @[DCache.scala 56:22]
  reg  valid_640; // @[DCache.scala 56:22]
  reg  valid_641; // @[DCache.scala 56:22]
  reg  valid_642; // @[DCache.scala 56:22]
  reg  valid_643; // @[DCache.scala 56:22]
  reg  valid_644; // @[DCache.scala 56:22]
  reg  valid_645; // @[DCache.scala 56:22]
  reg  valid_646; // @[DCache.scala 56:22]
  reg  valid_647; // @[DCache.scala 56:22]
  reg  valid_648; // @[DCache.scala 56:22]
  reg  valid_649; // @[DCache.scala 56:22]
  reg  valid_650; // @[DCache.scala 56:22]
  reg  valid_651; // @[DCache.scala 56:22]
  reg  valid_652; // @[DCache.scala 56:22]
  reg  valid_653; // @[DCache.scala 56:22]
  reg  valid_654; // @[DCache.scala 56:22]
  reg  valid_655; // @[DCache.scala 56:22]
  reg  valid_656; // @[DCache.scala 56:22]
  reg  valid_657; // @[DCache.scala 56:22]
  reg  valid_658; // @[DCache.scala 56:22]
  reg  valid_659; // @[DCache.scala 56:22]
  reg  valid_660; // @[DCache.scala 56:22]
  reg  valid_661; // @[DCache.scala 56:22]
  reg  valid_662; // @[DCache.scala 56:22]
  reg  valid_663; // @[DCache.scala 56:22]
  reg  valid_664; // @[DCache.scala 56:22]
  reg  valid_665; // @[DCache.scala 56:22]
  reg  valid_666; // @[DCache.scala 56:22]
  reg  valid_667; // @[DCache.scala 56:22]
  reg  valid_668; // @[DCache.scala 56:22]
  reg  valid_669; // @[DCache.scala 56:22]
  reg  valid_670; // @[DCache.scala 56:22]
  reg  valid_671; // @[DCache.scala 56:22]
  reg  valid_672; // @[DCache.scala 56:22]
  reg  valid_673; // @[DCache.scala 56:22]
  reg  valid_674; // @[DCache.scala 56:22]
  reg  valid_675; // @[DCache.scala 56:22]
  reg  valid_676; // @[DCache.scala 56:22]
  reg  valid_677; // @[DCache.scala 56:22]
  reg  valid_678; // @[DCache.scala 56:22]
  reg  valid_679; // @[DCache.scala 56:22]
  reg  valid_680; // @[DCache.scala 56:22]
  reg  valid_681; // @[DCache.scala 56:22]
  reg  valid_682; // @[DCache.scala 56:22]
  reg  valid_683; // @[DCache.scala 56:22]
  reg  valid_684; // @[DCache.scala 56:22]
  reg  valid_685; // @[DCache.scala 56:22]
  reg  valid_686; // @[DCache.scala 56:22]
  reg  valid_687; // @[DCache.scala 56:22]
  reg  valid_688; // @[DCache.scala 56:22]
  reg  valid_689; // @[DCache.scala 56:22]
  reg  valid_690; // @[DCache.scala 56:22]
  reg  valid_691; // @[DCache.scala 56:22]
  reg  valid_692; // @[DCache.scala 56:22]
  reg  valid_693; // @[DCache.scala 56:22]
  reg  valid_694; // @[DCache.scala 56:22]
  reg  valid_695; // @[DCache.scala 56:22]
  reg  valid_696; // @[DCache.scala 56:22]
  reg  valid_697; // @[DCache.scala 56:22]
  reg  valid_698; // @[DCache.scala 56:22]
  reg  valid_699; // @[DCache.scala 56:22]
  reg  valid_700; // @[DCache.scala 56:22]
  reg  valid_701; // @[DCache.scala 56:22]
  reg  valid_702; // @[DCache.scala 56:22]
  reg  valid_703; // @[DCache.scala 56:22]
  reg  valid_704; // @[DCache.scala 56:22]
  reg  valid_705; // @[DCache.scala 56:22]
  reg  valid_706; // @[DCache.scala 56:22]
  reg  valid_707; // @[DCache.scala 56:22]
  reg  valid_708; // @[DCache.scala 56:22]
  reg  valid_709; // @[DCache.scala 56:22]
  reg  valid_710; // @[DCache.scala 56:22]
  reg  valid_711; // @[DCache.scala 56:22]
  reg  valid_712; // @[DCache.scala 56:22]
  reg  valid_713; // @[DCache.scala 56:22]
  reg  valid_714; // @[DCache.scala 56:22]
  reg  valid_715; // @[DCache.scala 56:22]
  reg  valid_716; // @[DCache.scala 56:22]
  reg  valid_717; // @[DCache.scala 56:22]
  reg  valid_718; // @[DCache.scala 56:22]
  reg  valid_719; // @[DCache.scala 56:22]
  reg  valid_720; // @[DCache.scala 56:22]
  reg  valid_721; // @[DCache.scala 56:22]
  reg  valid_722; // @[DCache.scala 56:22]
  reg  valid_723; // @[DCache.scala 56:22]
  reg  valid_724; // @[DCache.scala 56:22]
  reg  valid_725; // @[DCache.scala 56:22]
  reg  valid_726; // @[DCache.scala 56:22]
  reg  valid_727; // @[DCache.scala 56:22]
  reg  valid_728; // @[DCache.scala 56:22]
  reg  valid_729; // @[DCache.scala 56:22]
  reg  valid_730; // @[DCache.scala 56:22]
  reg  valid_731; // @[DCache.scala 56:22]
  reg  valid_732; // @[DCache.scala 56:22]
  reg  valid_733; // @[DCache.scala 56:22]
  reg  valid_734; // @[DCache.scala 56:22]
  reg  valid_735; // @[DCache.scala 56:22]
  reg  valid_736; // @[DCache.scala 56:22]
  reg  valid_737; // @[DCache.scala 56:22]
  reg  valid_738; // @[DCache.scala 56:22]
  reg  valid_739; // @[DCache.scala 56:22]
  reg  valid_740; // @[DCache.scala 56:22]
  reg  valid_741; // @[DCache.scala 56:22]
  reg  valid_742; // @[DCache.scala 56:22]
  reg  valid_743; // @[DCache.scala 56:22]
  reg  valid_744; // @[DCache.scala 56:22]
  reg  valid_745; // @[DCache.scala 56:22]
  reg  valid_746; // @[DCache.scala 56:22]
  reg  valid_747; // @[DCache.scala 56:22]
  reg  valid_748; // @[DCache.scala 56:22]
  reg  valid_749; // @[DCache.scala 56:22]
  reg  valid_750; // @[DCache.scala 56:22]
  reg  valid_751; // @[DCache.scala 56:22]
  reg  valid_752; // @[DCache.scala 56:22]
  reg  valid_753; // @[DCache.scala 56:22]
  reg  valid_754; // @[DCache.scala 56:22]
  reg  valid_755; // @[DCache.scala 56:22]
  reg  valid_756; // @[DCache.scala 56:22]
  reg  valid_757; // @[DCache.scala 56:22]
  reg  valid_758; // @[DCache.scala 56:22]
  reg  valid_759; // @[DCache.scala 56:22]
  reg  valid_760; // @[DCache.scala 56:22]
  reg  valid_761; // @[DCache.scala 56:22]
  reg  valid_762; // @[DCache.scala 56:22]
  reg  valid_763; // @[DCache.scala 56:22]
  reg  valid_764; // @[DCache.scala 56:22]
  reg  valid_765; // @[DCache.scala 56:22]
  reg  valid_766; // @[DCache.scala 56:22]
  reg  valid_767; // @[DCache.scala 56:22]
  reg  valid_768; // @[DCache.scala 56:22]
  reg  valid_769; // @[DCache.scala 56:22]
  reg  valid_770; // @[DCache.scala 56:22]
  reg  valid_771; // @[DCache.scala 56:22]
  reg  valid_772; // @[DCache.scala 56:22]
  reg  valid_773; // @[DCache.scala 56:22]
  reg  valid_774; // @[DCache.scala 56:22]
  reg  valid_775; // @[DCache.scala 56:22]
  reg  valid_776; // @[DCache.scala 56:22]
  reg  valid_777; // @[DCache.scala 56:22]
  reg  valid_778; // @[DCache.scala 56:22]
  reg  valid_779; // @[DCache.scala 56:22]
  reg  valid_780; // @[DCache.scala 56:22]
  reg  valid_781; // @[DCache.scala 56:22]
  reg  valid_782; // @[DCache.scala 56:22]
  reg  valid_783; // @[DCache.scala 56:22]
  reg  valid_784; // @[DCache.scala 56:22]
  reg  valid_785; // @[DCache.scala 56:22]
  reg  valid_786; // @[DCache.scala 56:22]
  reg  valid_787; // @[DCache.scala 56:22]
  reg  valid_788; // @[DCache.scala 56:22]
  reg  valid_789; // @[DCache.scala 56:22]
  reg  valid_790; // @[DCache.scala 56:22]
  reg  valid_791; // @[DCache.scala 56:22]
  reg  valid_792; // @[DCache.scala 56:22]
  reg  valid_793; // @[DCache.scala 56:22]
  reg  valid_794; // @[DCache.scala 56:22]
  reg  valid_795; // @[DCache.scala 56:22]
  reg  valid_796; // @[DCache.scala 56:22]
  reg  valid_797; // @[DCache.scala 56:22]
  reg  valid_798; // @[DCache.scala 56:22]
  reg  valid_799; // @[DCache.scala 56:22]
  reg  valid_800; // @[DCache.scala 56:22]
  reg  valid_801; // @[DCache.scala 56:22]
  reg  valid_802; // @[DCache.scala 56:22]
  reg  valid_803; // @[DCache.scala 56:22]
  reg  valid_804; // @[DCache.scala 56:22]
  reg  valid_805; // @[DCache.scala 56:22]
  reg  valid_806; // @[DCache.scala 56:22]
  reg  valid_807; // @[DCache.scala 56:22]
  reg  valid_808; // @[DCache.scala 56:22]
  reg  valid_809; // @[DCache.scala 56:22]
  reg  valid_810; // @[DCache.scala 56:22]
  reg  valid_811; // @[DCache.scala 56:22]
  reg  valid_812; // @[DCache.scala 56:22]
  reg  valid_813; // @[DCache.scala 56:22]
  reg  valid_814; // @[DCache.scala 56:22]
  reg  valid_815; // @[DCache.scala 56:22]
  reg  valid_816; // @[DCache.scala 56:22]
  reg  valid_817; // @[DCache.scala 56:22]
  reg  valid_818; // @[DCache.scala 56:22]
  reg  valid_819; // @[DCache.scala 56:22]
  reg  valid_820; // @[DCache.scala 56:22]
  reg  valid_821; // @[DCache.scala 56:22]
  reg  valid_822; // @[DCache.scala 56:22]
  reg  valid_823; // @[DCache.scala 56:22]
  reg  valid_824; // @[DCache.scala 56:22]
  reg  valid_825; // @[DCache.scala 56:22]
  reg  valid_826; // @[DCache.scala 56:22]
  reg  valid_827; // @[DCache.scala 56:22]
  reg  valid_828; // @[DCache.scala 56:22]
  reg  valid_829; // @[DCache.scala 56:22]
  reg  valid_830; // @[DCache.scala 56:22]
  reg  valid_831; // @[DCache.scala 56:22]
  reg  valid_832; // @[DCache.scala 56:22]
  reg  valid_833; // @[DCache.scala 56:22]
  reg  valid_834; // @[DCache.scala 56:22]
  reg  valid_835; // @[DCache.scala 56:22]
  reg  valid_836; // @[DCache.scala 56:22]
  reg  valid_837; // @[DCache.scala 56:22]
  reg  valid_838; // @[DCache.scala 56:22]
  reg  valid_839; // @[DCache.scala 56:22]
  reg  valid_840; // @[DCache.scala 56:22]
  reg  valid_841; // @[DCache.scala 56:22]
  reg  valid_842; // @[DCache.scala 56:22]
  reg  valid_843; // @[DCache.scala 56:22]
  reg  valid_844; // @[DCache.scala 56:22]
  reg  valid_845; // @[DCache.scala 56:22]
  reg  valid_846; // @[DCache.scala 56:22]
  reg  valid_847; // @[DCache.scala 56:22]
  reg  valid_848; // @[DCache.scala 56:22]
  reg  valid_849; // @[DCache.scala 56:22]
  reg  valid_850; // @[DCache.scala 56:22]
  reg  valid_851; // @[DCache.scala 56:22]
  reg  valid_852; // @[DCache.scala 56:22]
  reg  valid_853; // @[DCache.scala 56:22]
  reg  valid_854; // @[DCache.scala 56:22]
  reg  valid_855; // @[DCache.scala 56:22]
  reg  valid_856; // @[DCache.scala 56:22]
  reg  valid_857; // @[DCache.scala 56:22]
  reg  valid_858; // @[DCache.scala 56:22]
  reg  valid_859; // @[DCache.scala 56:22]
  reg  valid_860; // @[DCache.scala 56:22]
  reg  valid_861; // @[DCache.scala 56:22]
  reg  valid_862; // @[DCache.scala 56:22]
  reg  valid_863; // @[DCache.scala 56:22]
  reg  valid_864; // @[DCache.scala 56:22]
  reg  valid_865; // @[DCache.scala 56:22]
  reg  valid_866; // @[DCache.scala 56:22]
  reg  valid_867; // @[DCache.scala 56:22]
  reg  valid_868; // @[DCache.scala 56:22]
  reg  valid_869; // @[DCache.scala 56:22]
  reg  valid_870; // @[DCache.scala 56:22]
  reg  valid_871; // @[DCache.scala 56:22]
  reg  valid_872; // @[DCache.scala 56:22]
  reg  valid_873; // @[DCache.scala 56:22]
  reg  valid_874; // @[DCache.scala 56:22]
  reg  valid_875; // @[DCache.scala 56:22]
  reg  valid_876; // @[DCache.scala 56:22]
  reg  valid_877; // @[DCache.scala 56:22]
  reg  valid_878; // @[DCache.scala 56:22]
  reg  valid_879; // @[DCache.scala 56:22]
  reg  valid_880; // @[DCache.scala 56:22]
  reg  valid_881; // @[DCache.scala 56:22]
  reg  valid_882; // @[DCache.scala 56:22]
  reg  valid_883; // @[DCache.scala 56:22]
  reg  valid_884; // @[DCache.scala 56:22]
  reg  valid_885; // @[DCache.scala 56:22]
  reg  valid_886; // @[DCache.scala 56:22]
  reg  valid_887; // @[DCache.scala 56:22]
  reg  valid_888; // @[DCache.scala 56:22]
  reg  valid_889; // @[DCache.scala 56:22]
  reg  valid_890; // @[DCache.scala 56:22]
  reg  valid_891; // @[DCache.scala 56:22]
  reg  valid_892; // @[DCache.scala 56:22]
  reg  valid_893; // @[DCache.scala 56:22]
  reg  valid_894; // @[DCache.scala 56:22]
  reg  valid_895; // @[DCache.scala 56:22]
  reg  valid_896; // @[DCache.scala 56:22]
  reg  valid_897; // @[DCache.scala 56:22]
  reg  valid_898; // @[DCache.scala 56:22]
  reg  valid_899; // @[DCache.scala 56:22]
  reg  valid_900; // @[DCache.scala 56:22]
  reg  valid_901; // @[DCache.scala 56:22]
  reg  valid_902; // @[DCache.scala 56:22]
  reg  valid_903; // @[DCache.scala 56:22]
  reg  valid_904; // @[DCache.scala 56:22]
  reg  valid_905; // @[DCache.scala 56:22]
  reg  valid_906; // @[DCache.scala 56:22]
  reg  valid_907; // @[DCache.scala 56:22]
  reg  valid_908; // @[DCache.scala 56:22]
  reg  valid_909; // @[DCache.scala 56:22]
  reg  valid_910; // @[DCache.scala 56:22]
  reg  valid_911; // @[DCache.scala 56:22]
  reg  valid_912; // @[DCache.scala 56:22]
  reg  valid_913; // @[DCache.scala 56:22]
  reg  valid_914; // @[DCache.scala 56:22]
  reg  valid_915; // @[DCache.scala 56:22]
  reg  valid_916; // @[DCache.scala 56:22]
  reg  valid_917; // @[DCache.scala 56:22]
  reg  valid_918; // @[DCache.scala 56:22]
  reg  valid_919; // @[DCache.scala 56:22]
  reg  valid_920; // @[DCache.scala 56:22]
  reg  valid_921; // @[DCache.scala 56:22]
  reg  valid_922; // @[DCache.scala 56:22]
  reg  valid_923; // @[DCache.scala 56:22]
  reg  valid_924; // @[DCache.scala 56:22]
  reg  valid_925; // @[DCache.scala 56:22]
  reg  valid_926; // @[DCache.scala 56:22]
  reg  valid_927; // @[DCache.scala 56:22]
  reg  valid_928; // @[DCache.scala 56:22]
  reg  valid_929; // @[DCache.scala 56:22]
  reg  valid_930; // @[DCache.scala 56:22]
  reg  valid_931; // @[DCache.scala 56:22]
  reg  valid_932; // @[DCache.scala 56:22]
  reg  valid_933; // @[DCache.scala 56:22]
  reg  valid_934; // @[DCache.scala 56:22]
  reg  valid_935; // @[DCache.scala 56:22]
  reg  valid_936; // @[DCache.scala 56:22]
  reg  valid_937; // @[DCache.scala 56:22]
  reg  valid_938; // @[DCache.scala 56:22]
  reg  valid_939; // @[DCache.scala 56:22]
  reg  valid_940; // @[DCache.scala 56:22]
  reg  valid_941; // @[DCache.scala 56:22]
  reg  valid_942; // @[DCache.scala 56:22]
  reg  valid_943; // @[DCache.scala 56:22]
  reg  valid_944; // @[DCache.scala 56:22]
  reg  valid_945; // @[DCache.scala 56:22]
  reg  valid_946; // @[DCache.scala 56:22]
  reg  valid_947; // @[DCache.scala 56:22]
  reg  valid_948; // @[DCache.scala 56:22]
  reg  valid_949; // @[DCache.scala 56:22]
  reg  valid_950; // @[DCache.scala 56:22]
  reg  valid_951; // @[DCache.scala 56:22]
  reg  valid_952; // @[DCache.scala 56:22]
  reg  valid_953; // @[DCache.scala 56:22]
  reg  valid_954; // @[DCache.scala 56:22]
  reg  valid_955; // @[DCache.scala 56:22]
  reg  valid_956; // @[DCache.scala 56:22]
  reg  valid_957; // @[DCache.scala 56:22]
  reg  valid_958; // @[DCache.scala 56:22]
  reg  valid_959; // @[DCache.scala 56:22]
  reg  valid_960; // @[DCache.scala 56:22]
  reg  valid_961; // @[DCache.scala 56:22]
  reg  valid_962; // @[DCache.scala 56:22]
  reg  valid_963; // @[DCache.scala 56:22]
  reg  valid_964; // @[DCache.scala 56:22]
  reg  valid_965; // @[DCache.scala 56:22]
  reg  valid_966; // @[DCache.scala 56:22]
  reg  valid_967; // @[DCache.scala 56:22]
  reg  valid_968; // @[DCache.scala 56:22]
  reg  valid_969; // @[DCache.scala 56:22]
  reg  valid_970; // @[DCache.scala 56:22]
  reg  valid_971; // @[DCache.scala 56:22]
  reg  valid_972; // @[DCache.scala 56:22]
  reg  valid_973; // @[DCache.scala 56:22]
  reg  valid_974; // @[DCache.scala 56:22]
  reg  valid_975; // @[DCache.scala 56:22]
  reg  valid_976; // @[DCache.scala 56:22]
  reg  valid_977; // @[DCache.scala 56:22]
  reg  valid_978; // @[DCache.scala 56:22]
  reg  valid_979; // @[DCache.scala 56:22]
  reg  valid_980; // @[DCache.scala 56:22]
  reg  valid_981; // @[DCache.scala 56:22]
  reg  valid_982; // @[DCache.scala 56:22]
  reg  valid_983; // @[DCache.scala 56:22]
  reg  valid_984; // @[DCache.scala 56:22]
  reg  valid_985; // @[DCache.scala 56:22]
  reg  valid_986; // @[DCache.scala 56:22]
  reg  valid_987; // @[DCache.scala 56:22]
  reg  valid_988; // @[DCache.scala 56:22]
  reg  valid_989; // @[DCache.scala 56:22]
  reg  valid_990; // @[DCache.scala 56:22]
  reg  valid_991; // @[DCache.scala 56:22]
  reg  valid_992; // @[DCache.scala 56:22]
  reg  valid_993; // @[DCache.scala 56:22]
  reg  valid_994; // @[DCache.scala 56:22]
  reg  valid_995; // @[DCache.scala 56:22]
  reg  valid_996; // @[DCache.scala 56:22]
  reg  valid_997; // @[DCache.scala 56:22]
  reg  valid_998; // @[DCache.scala 56:22]
  reg  valid_999; // @[DCache.scala 56:22]
  reg  valid_1000; // @[DCache.scala 56:22]
  reg  valid_1001; // @[DCache.scala 56:22]
  reg  valid_1002; // @[DCache.scala 56:22]
  reg  valid_1003; // @[DCache.scala 56:22]
  reg  valid_1004; // @[DCache.scala 56:22]
  reg  valid_1005; // @[DCache.scala 56:22]
  reg  valid_1006; // @[DCache.scala 56:22]
  reg  valid_1007; // @[DCache.scala 56:22]
  reg  valid_1008; // @[DCache.scala 56:22]
  reg  valid_1009; // @[DCache.scala 56:22]
  reg  valid_1010; // @[DCache.scala 56:22]
  reg  valid_1011; // @[DCache.scala 56:22]
  reg  valid_1012; // @[DCache.scala 56:22]
  reg  valid_1013; // @[DCache.scala 56:22]
  reg  valid_1014; // @[DCache.scala 56:22]
  reg  valid_1015; // @[DCache.scala 56:22]
  reg  valid_1016; // @[DCache.scala 56:22]
  reg  valid_1017; // @[DCache.scala 56:22]
  reg  valid_1018; // @[DCache.scala 56:22]
  reg  valid_1019; // @[DCache.scala 56:22]
  reg  valid_1020; // @[DCache.scala 56:22]
  reg  valid_1021; // @[DCache.scala 56:22]
  reg  valid_1022; // @[DCache.scala 56:22]
  reg  valid_1023; // @[DCache.scala 56:22]
  wire [31:0] array_addr = _GEN_16[31:0]; // @[DCache.scala 63:24 64:14]
  wire [16:0] array_wdata_tag = array_addr[31:15]; // @[DCache.scala 53:29]
  wire  _array_io_en_T_1 = io_cache_resp_ready & io_cache_resp_valid; // @[Decoupled.scala 51:35]
  wire  _T_11 = state == 3'h7; // @[DCache.scala 165:16]
  wire  amo_w = req_r_len == 2'h2; // @[DCache.scala 98:37]
  wire [31:0] _amo_wdata_raw_64_T_4 = req_r_addr[2] ? req_r_wdata[63:32] : req_r_wdata[31:0]; // @[DCache.scala 106:21]
  wire [31:0] _amo_wdata_raw_64_T_7 = _amo_wdata_raw_64_T_4[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _amo_wdata_raw_64_T_8 = {_amo_wdata_raw_64_T_7,_amo_wdata_raw_64_T_4}; // @[Cat.scala 33:92]
  wire [63:0] amo_wdata_raw_64 = amo_w ? _amo_wdata_raw_64_T_8 : req_r_wdata; // @[DCache.scala 104:26]
  reg  array_out_REG; // @[DCache.scala 76:55]
  reg [272:0] array_out_r; // @[Reg.scala 35:20]
  wire [272:0] _array_out_T_1 = array_out_REG ? array_io_rdata : array_out_r; // @[Utils.scala 50:8]
  wire [255:0] array_out_data = _array_out_T_1[255:0]; // @[DCache.scala 76:75]
  wire [255:0] rdata_256 = _T_11 ? tl_d_bits_r_data : array_out_data; // @[DCache.scala 81:22]
  wire [63:0] _rdata_64_T_6 = 2'h1 == array_addr[4:3] ? rdata_256[127:64] : rdata_256[63:0]; // @[Mux.scala 81:58]
  wire [63:0] _rdata_64_T_8 = 2'h2 == array_addr[4:3] ? rdata_256[191:128] : _rdata_64_T_6; // @[Mux.scala 81:58]
  wire [63:0] rdata_64 = 2'h3 == array_addr[4:3] ? rdata_256[255:192] : _rdata_64_T_8; // @[Mux.scala 81:58]
  wire [31:0] _amo_rdata_raw_64_T_4 = req_r_addr[2] ? rdata_64[63:32] : rdata_64[31:0]; // @[DCache.scala 101:21]
  wire [31:0] _amo_rdata_raw_64_T_7 = _amo_rdata_raw_64_T_4[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _amo_rdata_raw_64_T_8 = {_amo_rdata_raw_64_T_7,_amo_rdata_raw_64_T_4}; // @[Cat.scala 33:92]
  wire [63:0] amo_rdata_raw_64 = amo_w ? _amo_rdata_raw_64_T_8 : rdata_64; // @[DCache.scala 99:26]
  wire [63:0] _amo_result_64_T_16 = amo_wdata_raw_64 < amo_rdata_raw_64 ? amo_wdata_raw_64 : amo_rdata_raw_64; // @[DCache.scala 121:32]
  wire [63:0] _amo_result_64_T_11 = amo_w ? _amo_wdata_raw_64_T_8 : req_r_wdata; // @[DCache.scala 120:50]
  wire [63:0] _amo_result_64_T_12 = amo_w ? _amo_rdata_raw_64_T_8 : rdata_64; // @[DCache.scala 120:76]
  wire [63:0] _amo_result_64_T_14 = $signed(_amo_result_64_T_11) < $signed(_amo_result_64_T_12) ? amo_wdata_raw_64 :
    amo_rdata_raw_64; // @[DCache.scala 120:32]
  wire [63:0] _amo_result_64_T_10 = amo_wdata_raw_64 > amo_rdata_raw_64 ? amo_wdata_raw_64 : amo_rdata_raw_64; // @[DCache.scala 119:32]
  wire [63:0] _amo_result_64_T_8 = $signed(_amo_result_64_T_11) > $signed(_amo_result_64_T_12) ? amo_wdata_raw_64 :
    amo_rdata_raw_64; // @[DCache.scala 118:32]
  wire [63:0] _amo_result_64_T_4 = amo_wdata_raw_64 ^ amo_rdata_raw_64; // @[DCache.scala 117:47]
  wire [63:0] _amo_result_64_T_3 = amo_wdata_raw_64 | amo_rdata_raw_64; // @[DCache.scala 116:47]
  wire [63:0] _amo_result_64_T_2 = amo_wdata_raw_64 & amo_rdata_raw_64; // @[DCache.scala 115:47]
  wire [63:0] _amo_result_64_T_1 = amo_wdata_raw_64 + amo_rdata_raw_64; // @[DCache.scala 114:47]
  wire [63:0] _amo_result_64_T_18 = 5'h1b == req_r_amo ? amo_wdata_raw_64 : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _amo_result_64_T_20 = 5'h14 == req_r_amo ? _amo_result_64_T_1 : _amo_result_64_T_18; // @[Mux.scala 81:58]
  wire [63:0] _amo_result_64_T_22 = 5'h1a == req_r_amo ? _amo_result_64_T_2 : _amo_result_64_T_20; // @[Mux.scala 81:58]
  wire [63:0] _amo_result_64_T_24 = 5'h19 == req_r_amo ? _amo_result_64_T_3 : _amo_result_64_T_22; // @[Mux.scala 81:58]
  wire [63:0] _amo_result_64_T_26 = 5'h18 == req_r_amo ? _amo_result_64_T_4 : _amo_result_64_T_24; // @[Mux.scala 81:58]
  wire [63:0] _amo_result_64_T_28 = 5'h11 == req_r_amo ? _amo_result_64_T_8 : _amo_result_64_T_26; // @[Mux.scala 81:58]
  wire [63:0] _amo_result_64_T_30 = 5'h13 == req_r_amo ? _amo_result_64_T_10 : _amo_result_64_T_28; // @[Mux.scala 81:58]
  wire [63:0] _amo_result_64_T_32 = 5'h10 == req_r_amo ? _amo_result_64_T_14 : _amo_result_64_T_30; // @[Mux.scala 81:58]
  wire [63:0] amo_result_64 = 5'h12 == req_r_amo ? _amo_result_64_T_16 : _amo_result_64_T_32; // @[Mux.scala 81:58]
  wire [63:0] _amo_wdata_64_T_4 = {amo_result_64[31:0],32'h0}; // @[Cat.scala 33:92]
  wire [63:0] amo_wdata_64 = amo_w & req_r_addr[2] ? _amo_wdata_64_T_4 : amo_result_64; // @[DCache.scala 124:22]
  wire [63:0] wdata_64 = req_r_amo[4] ? amo_wdata_64 : req_r_wdata; // @[DCache.scala 157:22]
  wire [7:0] _wdata_256_T_1 = {req_r_addr[4:3], 6'h0}; // @[DCache.scala 160:51]
  wire [318:0] _GEN_0 = {{255'd0}, wdata_64}; // @[DCache.scala 160:25]
  wire [318:0] _wdata_256_T_2 = _GEN_0 << _wdata_256_T_1; // @[DCache.scala 160:25]
  wire [255:0] wdata_256 = _wdata_256_T_2[255:0]; // @[DCache.scala 158:23 160:13]
  wire [7:0] _wmask_256_T_23 = req_r_wmask[7] ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _wmask_256_T_21 = req_r_wmask[6] ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _wmask_256_T_19 = req_r_wmask[5] ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _wmask_256_T_17 = req_r_wmask[4] ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _wmask_256_T_15 = req_r_wmask[3] ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _wmask_256_T_13 = req_r_wmask[2] ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _wmask_256_T_11 = req_r_wmask[1] ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _wmask_256_T_9 = req_r_wmask[0] ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _wmask_256_T_24 = {_wmask_256_T_23,_wmask_256_T_21,_wmask_256_T_19,_wmask_256_T_17,_wmask_256_T_15,
    _wmask_256_T_13,_wmask_256_T_11,_wmask_256_T_9}; // @[Cat.scala 33:92]
  wire [318:0] _GEN_1 = {{255'd0}, _wmask_256_T_24}; // @[DCache.scala 161:40]
  wire [318:0] _wmask_256_T_27 = _GEN_1 << _wdata_256_T_1; // @[DCache.scala 161:40]
  wire [255:0] wmask_256 = _wmask_256_T_27[255:0]; // @[DCache.scala 159:23 161:13]
  wire [255:0] _array_wdata_data_T = wdata_256 & wmask_256; // @[Utils.scala 18:15]
  wire [255:0] _array_wdata_data_T_1 = ~wmask_256; // @[Utils.scala 18:38]
  wire [255:0] _array_wdata_data_T_2 = tl_d_bits_r_data & _array_wdata_data_T_1; // @[Utils.scala 18:35]
  wire [255:0] _array_wdata_data_T_3 = _array_wdata_data_T | _array_wdata_data_T_2; // @[Utils.scala 18:23]
  wire [255:0] _array_wdata_data_T_4 = req_r_wen ? _array_wdata_data_T_3 : tl_d_bits_r_data; // @[DCache.scala 166:30]
  wire [255:0] _array_wdata_data_T_7 = array_out_data & _array_wdata_data_T_1; // @[Utils.scala 18:35]
  wire [255:0] _array_wdata_data_T_8 = _array_wdata_data_T | _array_wdata_data_T_7; // @[Utils.scala 18:23]
  wire [255:0] _GEN_3106 = state == 3'h7 ? _array_wdata_data_T_4 : _array_wdata_data_T_8; // @[DCache.scala 165:26 166:24 176:24]
  wire [255:0] array_wdata_data = _array_io_en_T_1 ? _GEN_3106 : 256'h0; // @[DCache.scala 164:19 69:20]
  wire [16:0] array_out_tag = _array_out_T_1[272:256]; // @[DCache.scala 76:75]
  wire  _GEN_25 = 10'h1 == array_addr[14:5] ? valid_1 : valid_0; // @[DCache.scala 78:{33,33}]
  wire  _GEN_26 = 10'h2 == array_addr[14:5] ? valid_2 : _GEN_25; // @[DCache.scala 78:{33,33}]
  wire  _GEN_27 = 10'h3 == array_addr[14:5] ? valid_3 : _GEN_26; // @[DCache.scala 78:{33,33}]
  wire  _GEN_28 = 10'h4 == array_addr[14:5] ? valid_4 : _GEN_27; // @[DCache.scala 78:{33,33}]
  wire  _GEN_29 = 10'h5 == array_addr[14:5] ? valid_5 : _GEN_28; // @[DCache.scala 78:{33,33}]
  wire  _GEN_30 = 10'h6 == array_addr[14:5] ? valid_6 : _GEN_29; // @[DCache.scala 78:{33,33}]
  wire  _GEN_31 = 10'h7 == array_addr[14:5] ? valid_7 : _GEN_30; // @[DCache.scala 78:{33,33}]
  wire  _GEN_32 = 10'h8 == array_addr[14:5] ? valid_8 : _GEN_31; // @[DCache.scala 78:{33,33}]
  wire  _GEN_33 = 10'h9 == array_addr[14:5] ? valid_9 : _GEN_32; // @[DCache.scala 78:{33,33}]
  wire  _GEN_34 = 10'ha == array_addr[14:5] ? valid_10 : _GEN_33; // @[DCache.scala 78:{33,33}]
  wire  _GEN_35 = 10'hb == array_addr[14:5] ? valid_11 : _GEN_34; // @[DCache.scala 78:{33,33}]
  wire  _GEN_36 = 10'hc == array_addr[14:5] ? valid_12 : _GEN_35; // @[DCache.scala 78:{33,33}]
  wire  _GEN_37 = 10'hd == array_addr[14:5] ? valid_13 : _GEN_36; // @[DCache.scala 78:{33,33}]
  wire  _GEN_38 = 10'he == array_addr[14:5] ? valid_14 : _GEN_37; // @[DCache.scala 78:{33,33}]
  wire  _GEN_39 = 10'hf == array_addr[14:5] ? valid_15 : _GEN_38; // @[DCache.scala 78:{33,33}]
  wire  _GEN_40 = 10'h10 == array_addr[14:5] ? valid_16 : _GEN_39; // @[DCache.scala 78:{33,33}]
  wire  _GEN_41 = 10'h11 == array_addr[14:5] ? valid_17 : _GEN_40; // @[DCache.scala 78:{33,33}]
  wire  _GEN_42 = 10'h12 == array_addr[14:5] ? valid_18 : _GEN_41; // @[DCache.scala 78:{33,33}]
  wire  _GEN_43 = 10'h13 == array_addr[14:5] ? valid_19 : _GEN_42; // @[DCache.scala 78:{33,33}]
  wire  _GEN_44 = 10'h14 == array_addr[14:5] ? valid_20 : _GEN_43; // @[DCache.scala 78:{33,33}]
  wire  _GEN_45 = 10'h15 == array_addr[14:5] ? valid_21 : _GEN_44; // @[DCache.scala 78:{33,33}]
  wire  _GEN_46 = 10'h16 == array_addr[14:5] ? valid_22 : _GEN_45; // @[DCache.scala 78:{33,33}]
  wire  _GEN_47 = 10'h17 == array_addr[14:5] ? valid_23 : _GEN_46; // @[DCache.scala 78:{33,33}]
  wire  _GEN_48 = 10'h18 == array_addr[14:5] ? valid_24 : _GEN_47; // @[DCache.scala 78:{33,33}]
  wire  _GEN_49 = 10'h19 == array_addr[14:5] ? valid_25 : _GEN_48; // @[DCache.scala 78:{33,33}]
  wire  _GEN_50 = 10'h1a == array_addr[14:5] ? valid_26 : _GEN_49; // @[DCache.scala 78:{33,33}]
  wire  _GEN_51 = 10'h1b == array_addr[14:5] ? valid_27 : _GEN_50; // @[DCache.scala 78:{33,33}]
  wire  _GEN_52 = 10'h1c == array_addr[14:5] ? valid_28 : _GEN_51; // @[DCache.scala 78:{33,33}]
  wire  _GEN_53 = 10'h1d == array_addr[14:5] ? valid_29 : _GEN_52; // @[DCache.scala 78:{33,33}]
  wire  _GEN_54 = 10'h1e == array_addr[14:5] ? valid_30 : _GEN_53; // @[DCache.scala 78:{33,33}]
  wire  _GEN_55 = 10'h1f == array_addr[14:5] ? valid_31 : _GEN_54; // @[DCache.scala 78:{33,33}]
  wire  _GEN_56 = 10'h20 == array_addr[14:5] ? valid_32 : _GEN_55; // @[DCache.scala 78:{33,33}]
  wire  _GEN_57 = 10'h21 == array_addr[14:5] ? valid_33 : _GEN_56; // @[DCache.scala 78:{33,33}]
  wire  _GEN_58 = 10'h22 == array_addr[14:5] ? valid_34 : _GEN_57; // @[DCache.scala 78:{33,33}]
  wire  _GEN_59 = 10'h23 == array_addr[14:5] ? valid_35 : _GEN_58; // @[DCache.scala 78:{33,33}]
  wire  _GEN_60 = 10'h24 == array_addr[14:5] ? valid_36 : _GEN_59; // @[DCache.scala 78:{33,33}]
  wire  _GEN_61 = 10'h25 == array_addr[14:5] ? valid_37 : _GEN_60; // @[DCache.scala 78:{33,33}]
  wire  _GEN_62 = 10'h26 == array_addr[14:5] ? valid_38 : _GEN_61; // @[DCache.scala 78:{33,33}]
  wire  _GEN_63 = 10'h27 == array_addr[14:5] ? valid_39 : _GEN_62; // @[DCache.scala 78:{33,33}]
  wire  _GEN_64 = 10'h28 == array_addr[14:5] ? valid_40 : _GEN_63; // @[DCache.scala 78:{33,33}]
  wire  _GEN_65 = 10'h29 == array_addr[14:5] ? valid_41 : _GEN_64; // @[DCache.scala 78:{33,33}]
  wire  _GEN_66 = 10'h2a == array_addr[14:5] ? valid_42 : _GEN_65; // @[DCache.scala 78:{33,33}]
  wire  _GEN_67 = 10'h2b == array_addr[14:5] ? valid_43 : _GEN_66; // @[DCache.scala 78:{33,33}]
  wire  _GEN_68 = 10'h2c == array_addr[14:5] ? valid_44 : _GEN_67; // @[DCache.scala 78:{33,33}]
  wire  _GEN_69 = 10'h2d == array_addr[14:5] ? valid_45 : _GEN_68; // @[DCache.scala 78:{33,33}]
  wire  _GEN_70 = 10'h2e == array_addr[14:5] ? valid_46 : _GEN_69; // @[DCache.scala 78:{33,33}]
  wire  _GEN_71 = 10'h2f == array_addr[14:5] ? valid_47 : _GEN_70; // @[DCache.scala 78:{33,33}]
  wire  _GEN_72 = 10'h30 == array_addr[14:5] ? valid_48 : _GEN_71; // @[DCache.scala 78:{33,33}]
  wire  _GEN_73 = 10'h31 == array_addr[14:5] ? valid_49 : _GEN_72; // @[DCache.scala 78:{33,33}]
  wire  _GEN_74 = 10'h32 == array_addr[14:5] ? valid_50 : _GEN_73; // @[DCache.scala 78:{33,33}]
  wire  _GEN_75 = 10'h33 == array_addr[14:5] ? valid_51 : _GEN_74; // @[DCache.scala 78:{33,33}]
  wire  _GEN_76 = 10'h34 == array_addr[14:5] ? valid_52 : _GEN_75; // @[DCache.scala 78:{33,33}]
  wire  _GEN_77 = 10'h35 == array_addr[14:5] ? valid_53 : _GEN_76; // @[DCache.scala 78:{33,33}]
  wire  _GEN_78 = 10'h36 == array_addr[14:5] ? valid_54 : _GEN_77; // @[DCache.scala 78:{33,33}]
  wire  _GEN_79 = 10'h37 == array_addr[14:5] ? valid_55 : _GEN_78; // @[DCache.scala 78:{33,33}]
  wire  _GEN_80 = 10'h38 == array_addr[14:5] ? valid_56 : _GEN_79; // @[DCache.scala 78:{33,33}]
  wire  _GEN_81 = 10'h39 == array_addr[14:5] ? valid_57 : _GEN_80; // @[DCache.scala 78:{33,33}]
  wire  _GEN_82 = 10'h3a == array_addr[14:5] ? valid_58 : _GEN_81; // @[DCache.scala 78:{33,33}]
  wire  _GEN_83 = 10'h3b == array_addr[14:5] ? valid_59 : _GEN_82; // @[DCache.scala 78:{33,33}]
  wire  _GEN_84 = 10'h3c == array_addr[14:5] ? valid_60 : _GEN_83; // @[DCache.scala 78:{33,33}]
  wire  _GEN_85 = 10'h3d == array_addr[14:5] ? valid_61 : _GEN_84; // @[DCache.scala 78:{33,33}]
  wire  _GEN_86 = 10'h3e == array_addr[14:5] ? valid_62 : _GEN_85; // @[DCache.scala 78:{33,33}]
  wire  _GEN_87 = 10'h3f == array_addr[14:5] ? valid_63 : _GEN_86; // @[DCache.scala 78:{33,33}]
  wire  _GEN_88 = 10'h40 == array_addr[14:5] ? valid_64 : _GEN_87; // @[DCache.scala 78:{33,33}]
  wire  _GEN_89 = 10'h41 == array_addr[14:5] ? valid_65 : _GEN_88; // @[DCache.scala 78:{33,33}]
  wire  _GEN_90 = 10'h42 == array_addr[14:5] ? valid_66 : _GEN_89; // @[DCache.scala 78:{33,33}]
  wire  _GEN_91 = 10'h43 == array_addr[14:5] ? valid_67 : _GEN_90; // @[DCache.scala 78:{33,33}]
  wire  _GEN_92 = 10'h44 == array_addr[14:5] ? valid_68 : _GEN_91; // @[DCache.scala 78:{33,33}]
  wire  _GEN_93 = 10'h45 == array_addr[14:5] ? valid_69 : _GEN_92; // @[DCache.scala 78:{33,33}]
  wire  _GEN_94 = 10'h46 == array_addr[14:5] ? valid_70 : _GEN_93; // @[DCache.scala 78:{33,33}]
  wire  _GEN_95 = 10'h47 == array_addr[14:5] ? valid_71 : _GEN_94; // @[DCache.scala 78:{33,33}]
  wire  _GEN_96 = 10'h48 == array_addr[14:5] ? valid_72 : _GEN_95; // @[DCache.scala 78:{33,33}]
  wire  _GEN_97 = 10'h49 == array_addr[14:5] ? valid_73 : _GEN_96; // @[DCache.scala 78:{33,33}]
  wire  _GEN_98 = 10'h4a == array_addr[14:5] ? valid_74 : _GEN_97; // @[DCache.scala 78:{33,33}]
  wire  _GEN_99 = 10'h4b == array_addr[14:5] ? valid_75 : _GEN_98; // @[DCache.scala 78:{33,33}]
  wire  _GEN_100 = 10'h4c == array_addr[14:5] ? valid_76 : _GEN_99; // @[DCache.scala 78:{33,33}]
  wire  _GEN_101 = 10'h4d == array_addr[14:5] ? valid_77 : _GEN_100; // @[DCache.scala 78:{33,33}]
  wire  _GEN_102 = 10'h4e == array_addr[14:5] ? valid_78 : _GEN_101; // @[DCache.scala 78:{33,33}]
  wire  _GEN_103 = 10'h4f == array_addr[14:5] ? valid_79 : _GEN_102; // @[DCache.scala 78:{33,33}]
  wire  _GEN_104 = 10'h50 == array_addr[14:5] ? valid_80 : _GEN_103; // @[DCache.scala 78:{33,33}]
  wire  _GEN_105 = 10'h51 == array_addr[14:5] ? valid_81 : _GEN_104; // @[DCache.scala 78:{33,33}]
  wire  _GEN_106 = 10'h52 == array_addr[14:5] ? valid_82 : _GEN_105; // @[DCache.scala 78:{33,33}]
  wire  _GEN_107 = 10'h53 == array_addr[14:5] ? valid_83 : _GEN_106; // @[DCache.scala 78:{33,33}]
  wire  _GEN_108 = 10'h54 == array_addr[14:5] ? valid_84 : _GEN_107; // @[DCache.scala 78:{33,33}]
  wire  _GEN_109 = 10'h55 == array_addr[14:5] ? valid_85 : _GEN_108; // @[DCache.scala 78:{33,33}]
  wire  _GEN_110 = 10'h56 == array_addr[14:5] ? valid_86 : _GEN_109; // @[DCache.scala 78:{33,33}]
  wire  _GEN_111 = 10'h57 == array_addr[14:5] ? valid_87 : _GEN_110; // @[DCache.scala 78:{33,33}]
  wire  _GEN_112 = 10'h58 == array_addr[14:5] ? valid_88 : _GEN_111; // @[DCache.scala 78:{33,33}]
  wire  _GEN_113 = 10'h59 == array_addr[14:5] ? valid_89 : _GEN_112; // @[DCache.scala 78:{33,33}]
  wire  _GEN_114 = 10'h5a == array_addr[14:5] ? valid_90 : _GEN_113; // @[DCache.scala 78:{33,33}]
  wire  _GEN_115 = 10'h5b == array_addr[14:5] ? valid_91 : _GEN_114; // @[DCache.scala 78:{33,33}]
  wire  _GEN_116 = 10'h5c == array_addr[14:5] ? valid_92 : _GEN_115; // @[DCache.scala 78:{33,33}]
  wire  _GEN_117 = 10'h5d == array_addr[14:5] ? valid_93 : _GEN_116; // @[DCache.scala 78:{33,33}]
  wire  _GEN_118 = 10'h5e == array_addr[14:5] ? valid_94 : _GEN_117; // @[DCache.scala 78:{33,33}]
  wire  _GEN_119 = 10'h5f == array_addr[14:5] ? valid_95 : _GEN_118; // @[DCache.scala 78:{33,33}]
  wire  _GEN_120 = 10'h60 == array_addr[14:5] ? valid_96 : _GEN_119; // @[DCache.scala 78:{33,33}]
  wire  _GEN_121 = 10'h61 == array_addr[14:5] ? valid_97 : _GEN_120; // @[DCache.scala 78:{33,33}]
  wire  _GEN_122 = 10'h62 == array_addr[14:5] ? valid_98 : _GEN_121; // @[DCache.scala 78:{33,33}]
  wire  _GEN_123 = 10'h63 == array_addr[14:5] ? valid_99 : _GEN_122; // @[DCache.scala 78:{33,33}]
  wire  _GEN_124 = 10'h64 == array_addr[14:5] ? valid_100 : _GEN_123; // @[DCache.scala 78:{33,33}]
  wire  _GEN_125 = 10'h65 == array_addr[14:5] ? valid_101 : _GEN_124; // @[DCache.scala 78:{33,33}]
  wire  _GEN_126 = 10'h66 == array_addr[14:5] ? valid_102 : _GEN_125; // @[DCache.scala 78:{33,33}]
  wire  _GEN_127 = 10'h67 == array_addr[14:5] ? valid_103 : _GEN_126; // @[DCache.scala 78:{33,33}]
  wire  _GEN_128 = 10'h68 == array_addr[14:5] ? valid_104 : _GEN_127; // @[DCache.scala 78:{33,33}]
  wire  _GEN_129 = 10'h69 == array_addr[14:5] ? valid_105 : _GEN_128; // @[DCache.scala 78:{33,33}]
  wire  _GEN_130 = 10'h6a == array_addr[14:5] ? valid_106 : _GEN_129; // @[DCache.scala 78:{33,33}]
  wire  _GEN_131 = 10'h6b == array_addr[14:5] ? valid_107 : _GEN_130; // @[DCache.scala 78:{33,33}]
  wire  _GEN_132 = 10'h6c == array_addr[14:5] ? valid_108 : _GEN_131; // @[DCache.scala 78:{33,33}]
  wire  _GEN_133 = 10'h6d == array_addr[14:5] ? valid_109 : _GEN_132; // @[DCache.scala 78:{33,33}]
  wire  _GEN_134 = 10'h6e == array_addr[14:5] ? valid_110 : _GEN_133; // @[DCache.scala 78:{33,33}]
  wire  _GEN_135 = 10'h6f == array_addr[14:5] ? valid_111 : _GEN_134; // @[DCache.scala 78:{33,33}]
  wire  _GEN_136 = 10'h70 == array_addr[14:5] ? valid_112 : _GEN_135; // @[DCache.scala 78:{33,33}]
  wire  _GEN_137 = 10'h71 == array_addr[14:5] ? valid_113 : _GEN_136; // @[DCache.scala 78:{33,33}]
  wire  _GEN_138 = 10'h72 == array_addr[14:5] ? valid_114 : _GEN_137; // @[DCache.scala 78:{33,33}]
  wire  _GEN_139 = 10'h73 == array_addr[14:5] ? valid_115 : _GEN_138; // @[DCache.scala 78:{33,33}]
  wire  _GEN_140 = 10'h74 == array_addr[14:5] ? valid_116 : _GEN_139; // @[DCache.scala 78:{33,33}]
  wire  _GEN_141 = 10'h75 == array_addr[14:5] ? valid_117 : _GEN_140; // @[DCache.scala 78:{33,33}]
  wire  _GEN_142 = 10'h76 == array_addr[14:5] ? valid_118 : _GEN_141; // @[DCache.scala 78:{33,33}]
  wire  _GEN_143 = 10'h77 == array_addr[14:5] ? valid_119 : _GEN_142; // @[DCache.scala 78:{33,33}]
  wire  _GEN_144 = 10'h78 == array_addr[14:5] ? valid_120 : _GEN_143; // @[DCache.scala 78:{33,33}]
  wire  _GEN_145 = 10'h79 == array_addr[14:5] ? valid_121 : _GEN_144; // @[DCache.scala 78:{33,33}]
  wire  _GEN_146 = 10'h7a == array_addr[14:5] ? valid_122 : _GEN_145; // @[DCache.scala 78:{33,33}]
  wire  _GEN_147 = 10'h7b == array_addr[14:5] ? valid_123 : _GEN_146; // @[DCache.scala 78:{33,33}]
  wire  _GEN_148 = 10'h7c == array_addr[14:5] ? valid_124 : _GEN_147; // @[DCache.scala 78:{33,33}]
  wire  _GEN_149 = 10'h7d == array_addr[14:5] ? valid_125 : _GEN_148; // @[DCache.scala 78:{33,33}]
  wire  _GEN_150 = 10'h7e == array_addr[14:5] ? valid_126 : _GEN_149; // @[DCache.scala 78:{33,33}]
  wire  _GEN_151 = 10'h7f == array_addr[14:5] ? valid_127 : _GEN_150; // @[DCache.scala 78:{33,33}]
  wire  _GEN_152 = 10'h80 == array_addr[14:5] ? valid_128 : _GEN_151; // @[DCache.scala 78:{33,33}]
  wire  _GEN_153 = 10'h81 == array_addr[14:5] ? valid_129 : _GEN_152; // @[DCache.scala 78:{33,33}]
  wire  _GEN_154 = 10'h82 == array_addr[14:5] ? valid_130 : _GEN_153; // @[DCache.scala 78:{33,33}]
  wire  _GEN_155 = 10'h83 == array_addr[14:5] ? valid_131 : _GEN_154; // @[DCache.scala 78:{33,33}]
  wire  _GEN_156 = 10'h84 == array_addr[14:5] ? valid_132 : _GEN_155; // @[DCache.scala 78:{33,33}]
  wire  _GEN_157 = 10'h85 == array_addr[14:5] ? valid_133 : _GEN_156; // @[DCache.scala 78:{33,33}]
  wire  _GEN_158 = 10'h86 == array_addr[14:5] ? valid_134 : _GEN_157; // @[DCache.scala 78:{33,33}]
  wire  _GEN_159 = 10'h87 == array_addr[14:5] ? valid_135 : _GEN_158; // @[DCache.scala 78:{33,33}]
  wire  _GEN_160 = 10'h88 == array_addr[14:5] ? valid_136 : _GEN_159; // @[DCache.scala 78:{33,33}]
  wire  _GEN_161 = 10'h89 == array_addr[14:5] ? valid_137 : _GEN_160; // @[DCache.scala 78:{33,33}]
  wire  _GEN_162 = 10'h8a == array_addr[14:5] ? valid_138 : _GEN_161; // @[DCache.scala 78:{33,33}]
  wire  _GEN_163 = 10'h8b == array_addr[14:5] ? valid_139 : _GEN_162; // @[DCache.scala 78:{33,33}]
  wire  _GEN_164 = 10'h8c == array_addr[14:5] ? valid_140 : _GEN_163; // @[DCache.scala 78:{33,33}]
  wire  _GEN_165 = 10'h8d == array_addr[14:5] ? valid_141 : _GEN_164; // @[DCache.scala 78:{33,33}]
  wire  _GEN_166 = 10'h8e == array_addr[14:5] ? valid_142 : _GEN_165; // @[DCache.scala 78:{33,33}]
  wire  _GEN_167 = 10'h8f == array_addr[14:5] ? valid_143 : _GEN_166; // @[DCache.scala 78:{33,33}]
  wire  _GEN_168 = 10'h90 == array_addr[14:5] ? valid_144 : _GEN_167; // @[DCache.scala 78:{33,33}]
  wire  _GEN_169 = 10'h91 == array_addr[14:5] ? valid_145 : _GEN_168; // @[DCache.scala 78:{33,33}]
  wire  _GEN_170 = 10'h92 == array_addr[14:5] ? valid_146 : _GEN_169; // @[DCache.scala 78:{33,33}]
  wire  _GEN_171 = 10'h93 == array_addr[14:5] ? valid_147 : _GEN_170; // @[DCache.scala 78:{33,33}]
  wire  _GEN_172 = 10'h94 == array_addr[14:5] ? valid_148 : _GEN_171; // @[DCache.scala 78:{33,33}]
  wire  _GEN_173 = 10'h95 == array_addr[14:5] ? valid_149 : _GEN_172; // @[DCache.scala 78:{33,33}]
  wire  _GEN_174 = 10'h96 == array_addr[14:5] ? valid_150 : _GEN_173; // @[DCache.scala 78:{33,33}]
  wire  _GEN_175 = 10'h97 == array_addr[14:5] ? valid_151 : _GEN_174; // @[DCache.scala 78:{33,33}]
  wire  _GEN_176 = 10'h98 == array_addr[14:5] ? valid_152 : _GEN_175; // @[DCache.scala 78:{33,33}]
  wire  _GEN_177 = 10'h99 == array_addr[14:5] ? valid_153 : _GEN_176; // @[DCache.scala 78:{33,33}]
  wire  _GEN_178 = 10'h9a == array_addr[14:5] ? valid_154 : _GEN_177; // @[DCache.scala 78:{33,33}]
  wire  _GEN_179 = 10'h9b == array_addr[14:5] ? valid_155 : _GEN_178; // @[DCache.scala 78:{33,33}]
  wire  _GEN_180 = 10'h9c == array_addr[14:5] ? valid_156 : _GEN_179; // @[DCache.scala 78:{33,33}]
  wire  _GEN_181 = 10'h9d == array_addr[14:5] ? valid_157 : _GEN_180; // @[DCache.scala 78:{33,33}]
  wire  _GEN_182 = 10'h9e == array_addr[14:5] ? valid_158 : _GEN_181; // @[DCache.scala 78:{33,33}]
  wire  _GEN_183 = 10'h9f == array_addr[14:5] ? valid_159 : _GEN_182; // @[DCache.scala 78:{33,33}]
  wire  _GEN_184 = 10'ha0 == array_addr[14:5] ? valid_160 : _GEN_183; // @[DCache.scala 78:{33,33}]
  wire  _GEN_185 = 10'ha1 == array_addr[14:5] ? valid_161 : _GEN_184; // @[DCache.scala 78:{33,33}]
  wire  _GEN_186 = 10'ha2 == array_addr[14:5] ? valid_162 : _GEN_185; // @[DCache.scala 78:{33,33}]
  wire  _GEN_187 = 10'ha3 == array_addr[14:5] ? valid_163 : _GEN_186; // @[DCache.scala 78:{33,33}]
  wire  _GEN_188 = 10'ha4 == array_addr[14:5] ? valid_164 : _GEN_187; // @[DCache.scala 78:{33,33}]
  wire  _GEN_189 = 10'ha5 == array_addr[14:5] ? valid_165 : _GEN_188; // @[DCache.scala 78:{33,33}]
  wire  _GEN_190 = 10'ha6 == array_addr[14:5] ? valid_166 : _GEN_189; // @[DCache.scala 78:{33,33}]
  wire  _GEN_191 = 10'ha7 == array_addr[14:5] ? valid_167 : _GEN_190; // @[DCache.scala 78:{33,33}]
  wire  _GEN_192 = 10'ha8 == array_addr[14:5] ? valid_168 : _GEN_191; // @[DCache.scala 78:{33,33}]
  wire  _GEN_193 = 10'ha9 == array_addr[14:5] ? valid_169 : _GEN_192; // @[DCache.scala 78:{33,33}]
  wire  _GEN_194 = 10'haa == array_addr[14:5] ? valid_170 : _GEN_193; // @[DCache.scala 78:{33,33}]
  wire  _GEN_195 = 10'hab == array_addr[14:5] ? valid_171 : _GEN_194; // @[DCache.scala 78:{33,33}]
  wire  _GEN_196 = 10'hac == array_addr[14:5] ? valid_172 : _GEN_195; // @[DCache.scala 78:{33,33}]
  wire  _GEN_197 = 10'had == array_addr[14:5] ? valid_173 : _GEN_196; // @[DCache.scala 78:{33,33}]
  wire  _GEN_198 = 10'hae == array_addr[14:5] ? valid_174 : _GEN_197; // @[DCache.scala 78:{33,33}]
  wire  _GEN_199 = 10'haf == array_addr[14:5] ? valid_175 : _GEN_198; // @[DCache.scala 78:{33,33}]
  wire  _GEN_200 = 10'hb0 == array_addr[14:5] ? valid_176 : _GEN_199; // @[DCache.scala 78:{33,33}]
  wire  _GEN_201 = 10'hb1 == array_addr[14:5] ? valid_177 : _GEN_200; // @[DCache.scala 78:{33,33}]
  wire  _GEN_202 = 10'hb2 == array_addr[14:5] ? valid_178 : _GEN_201; // @[DCache.scala 78:{33,33}]
  wire  _GEN_203 = 10'hb3 == array_addr[14:5] ? valid_179 : _GEN_202; // @[DCache.scala 78:{33,33}]
  wire  _GEN_204 = 10'hb4 == array_addr[14:5] ? valid_180 : _GEN_203; // @[DCache.scala 78:{33,33}]
  wire  _GEN_205 = 10'hb5 == array_addr[14:5] ? valid_181 : _GEN_204; // @[DCache.scala 78:{33,33}]
  wire  _GEN_206 = 10'hb6 == array_addr[14:5] ? valid_182 : _GEN_205; // @[DCache.scala 78:{33,33}]
  wire  _GEN_207 = 10'hb7 == array_addr[14:5] ? valid_183 : _GEN_206; // @[DCache.scala 78:{33,33}]
  wire  _GEN_208 = 10'hb8 == array_addr[14:5] ? valid_184 : _GEN_207; // @[DCache.scala 78:{33,33}]
  wire  _GEN_209 = 10'hb9 == array_addr[14:5] ? valid_185 : _GEN_208; // @[DCache.scala 78:{33,33}]
  wire  _GEN_210 = 10'hba == array_addr[14:5] ? valid_186 : _GEN_209; // @[DCache.scala 78:{33,33}]
  wire  _GEN_211 = 10'hbb == array_addr[14:5] ? valid_187 : _GEN_210; // @[DCache.scala 78:{33,33}]
  wire  _GEN_212 = 10'hbc == array_addr[14:5] ? valid_188 : _GEN_211; // @[DCache.scala 78:{33,33}]
  wire  _GEN_213 = 10'hbd == array_addr[14:5] ? valid_189 : _GEN_212; // @[DCache.scala 78:{33,33}]
  wire  _GEN_214 = 10'hbe == array_addr[14:5] ? valid_190 : _GEN_213; // @[DCache.scala 78:{33,33}]
  wire  _GEN_215 = 10'hbf == array_addr[14:5] ? valid_191 : _GEN_214; // @[DCache.scala 78:{33,33}]
  wire  _GEN_216 = 10'hc0 == array_addr[14:5] ? valid_192 : _GEN_215; // @[DCache.scala 78:{33,33}]
  wire  _GEN_217 = 10'hc1 == array_addr[14:5] ? valid_193 : _GEN_216; // @[DCache.scala 78:{33,33}]
  wire  _GEN_218 = 10'hc2 == array_addr[14:5] ? valid_194 : _GEN_217; // @[DCache.scala 78:{33,33}]
  wire  _GEN_219 = 10'hc3 == array_addr[14:5] ? valid_195 : _GEN_218; // @[DCache.scala 78:{33,33}]
  wire  _GEN_220 = 10'hc4 == array_addr[14:5] ? valid_196 : _GEN_219; // @[DCache.scala 78:{33,33}]
  wire  _GEN_221 = 10'hc5 == array_addr[14:5] ? valid_197 : _GEN_220; // @[DCache.scala 78:{33,33}]
  wire  _GEN_222 = 10'hc6 == array_addr[14:5] ? valid_198 : _GEN_221; // @[DCache.scala 78:{33,33}]
  wire  _GEN_223 = 10'hc7 == array_addr[14:5] ? valid_199 : _GEN_222; // @[DCache.scala 78:{33,33}]
  wire  _GEN_224 = 10'hc8 == array_addr[14:5] ? valid_200 : _GEN_223; // @[DCache.scala 78:{33,33}]
  wire  _GEN_225 = 10'hc9 == array_addr[14:5] ? valid_201 : _GEN_224; // @[DCache.scala 78:{33,33}]
  wire  _GEN_226 = 10'hca == array_addr[14:5] ? valid_202 : _GEN_225; // @[DCache.scala 78:{33,33}]
  wire  _GEN_227 = 10'hcb == array_addr[14:5] ? valid_203 : _GEN_226; // @[DCache.scala 78:{33,33}]
  wire  _GEN_228 = 10'hcc == array_addr[14:5] ? valid_204 : _GEN_227; // @[DCache.scala 78:{33,33}]
  wire  _GEN_229 = 10'hcd == array_addr[14:5] ? valid_205 : _GEN_228; // @[DCache.scala 78:{33,33}]
  wire  _GEN_230 = 10'hce == array_addr[14:5] ? valid_206 : _GEN_229; // @[DCache.scala 78:{33,33}]
  wire  _GEN_231 = 10'hcf == array_addr[14:5] ? valid_207 : _GEN_230; // @[DCache.scala 78:{33,33}]
  wire  _GEN_232 = 10'hd0 == array_addr[14:5] ? valid_208 : _GEN_231; // @[DCache.scala 78:{33,33}]
  wire  _GEN_233 = 10'hd1 == array_addr[14:5] ? valid_209 : _GEN_232; // @[DCache.scala 78:{33,33}]
  wire  _GEN_234 = 10'hd2 == array_addr[14:5] ? valid_210 : _GEN_233; // @[DCache.scala 78:{33,33}]
  wire  _GEN_235 = 10'hd3 == array_addr[14:5] ? valid_211 : _GEN_234; // @[DCache.scala 78:{33,33}]
  wire  _GEN_236 = 10'hd4 == array_addr[14:5] ? valid_212 : _GEN_235; // @[DCache.scala 78:{33,33}]
  wire  _GEN_237 = 10'hd5 == array_addr[14:5] ? valid_213 : _GEN_236; // @[DCache.scala 78:{33,33}]
  wire  _GEN_238 = 10'hd6 == array_addr[14:5] ? valid_214 : _GEN_237; // @[DCache.scala 78:{33,33}]
  wire  _GEN_239 = 10'hd7 == array_addr[14:5] ? valid_215 : _GEN_238; // @[DCache.scala 78:{33,33}]
  wire  _GEN_240 = 10'hd8 == array_addr[14:5] ? valid_216 : _GEN_239; // @[DCache.scala 78:{33,33}]
  wire  _GEN_241 = 10'hd9 == array_addr[14:5] ? valid_217 : _GEN_240; // @[DCache.scala 78:{33,33}]
  wire  _GEN_242 = 10'hda == array_addr[14:5] ? valid_218 : _GEN_241; // @[DCache.scala 78:{33,33}]
  wire  _GEN_243 = 10'hdb == array_addr[14:5] ? valid_219 : _GEN_242; // @[DCache.scala 78:{33,33}]
  wire  _GEN_244 = 10'hdc == array_addr[14:5] ? valid_220 : _GEN_243; // @[DCache.scala 78:{33,33}]
  wire  _GEN_245 = 10'hdd == array_addr[14:5] ? valid_221 : _GEN_244; // @[DCache.scala 78:{33,33}]
  wire  _GEN_246 = 10'hde == array_addr[14:5] ? valid_222 : _GEN_245; // @[DCache.scala 78:{33,33}]
  wire  _GEN_247 = 10'hdf == array_addr[14:5] ? valid_223 : _GEN_246; // @[DCache.scala 78:{33,33}]
  wire  _GEN_248 = 10'he0 == array_addr[14:5] ? valid_224 : _GEN_247; // @[DCache.scala 78:{33,33}]
  wire  _GEN_249 = 10'he1 == array_addr[14:5] ? valid_225 : _GEN_248; // @[DCache.scala 78:{33,33}]
  wire  _GEN_250 = 10'he2 == array_addr[14:5] ? valid_226 : _GEN_249; // @[DCache.scala 78:{33,33}]
  wire  _GEN_251 = 10'he3 == array_addr[14:5] ? valid_227 : _GEN_250; // @[DCache.scala 78:{33,33}]
  wire  _GEN_252 = 10'he4 == array_addr[14:5] ? valid_228 : _GEN_251; // @[DCache.scala 78:{33,33}]
  wire  _GEN_253 = 10'he5 == array_addr[14:5] ? valid_229 : _GEN_252; // @[DCache.scala 78:{33,33}]
  wire  _GEN_254 = 10'he6 == array_addr[14:5] ? valid_230 : _GEN_253; // @[DCache.scala 78:{33,33}]
  wire  _GEN_255 = 10'he7 == array_addr[14:5] ? valid_231 : _GEN_254; // @[DCache.scala 78:{33,33}]
  wire  _GEN_256 = 10'he8 == array_addr[14:5] ? valid_232 : _GEN_255; // @[DCache.scala 78:{33,33}]
  wire  _GEN_257 = 10'he9 == array_addr[14:5] ? valid_233 : _GEN_256; // @[DCache.scala 78:{33,33}]
  wire  _GEN_258 = 10'hea == array_addr[14:5] ? valid_234 : _GEN_257; // @[DCache.scala 78:{33,33}]
  wire  _GEN_259 = 10'heb == array_addr[14:5] ? valid_235 : _GEN_258; // @[DCache.scala 78:{33,33}]
  wire  _GEN_260 = 10'hec == array_addr[14:5] ? valid_236 : _GEN_259; // @[DCache.scala 78:{33,33}]
  wire  _GEN_261 = 10'hed == array_addr[14:5] ? valid_237 : _GEN_260; // @[DCache.scala 78:{33,33}]
  wire  _GEN_262 = 10'hee == array_addr[14:5] ? valid_238 : _GEN_261; // @[DCache.scala 78:{33,33}]
  wire  _GEN_263 = 10'hef == array_addr[14:5] ? valid_239 : _GEN_262; // @[DCache.scala 78:{33,33}]
  wire  _GEN_264 = 10'hf0 == array_addr[14:5] ? valid_240 : _GEN_263; // @[DCache.scala 78:{33,33}]
  wire  _GEN_265 = 10'hf1 == array_addr[14:5] ? valid_241 : _GEN_264; // @[DCache.scala 78:{33,33}]
  wire  _GEN_266 = 10'hf2 == array_addr[14:5] ? valid_242 : _GEN_265; // @[DCache.scala 78:{33,33}]
  wire  _GEN_267 = 10'hf3 == array_addr[14:5] ? valid_243 : _GEN_266; // @[DCache.scala 78:{33,33}]
  wire  _GEN_268 = 10'hf4 == array_addr[14:5] ? valid_244 : _GEN_267; // @[DCache.scala 78:{33,33}]
  wire  _GEN_269 = 10'hf5 == array_addr[14:5] ? valid_245 : _GEN_268; // @[DCache.scala 78:{33,33}]
  wire  _GEN_270 = 10'hf6 == array_addr[14:5] ? valid_246 : _GEN_269; // @[DCache.scala 78:{33,33}]
  wire  _GEN_271 = 10'hf7 == array_addr[14:5] ? valid_247 : _GEN_270; // @[DCache.scala 78:{33,33}]
  wire  _GEN_272 = 10'hf8 == array_addr[14:5] ? valid_248 : _GEN_271; // @[DCache.scala 78:{33,33}]
  wire  _GEN_273 = 10'hf9 == array_addr[14:5] ? valid_249 : _GEN_272; // @[DCache.scala 78:{33,33}]
  wire  _GEN_274 = 10'hfa == array_addr[14:5] ? valid_250 : _GEN_273; // @[DCache.scala 78:{33,33}]
  wire  _GEN_275 = 10'hfb == array_addr[14:5] ? valid_251 : _GEN_274; // @[DCache.scala 78:{33,33}]
  wire  _GEN_276 = 10'hfc == array_addr[14:5] ? valid_252 : _GEN_275; // @[DCache.scala 78:{33,33}]
  wire  _GEN_277 = 10'hfd == array_addr[14:5] ? valid_253 : _GEN_276; // @[DCache.scala 78:{33,33}]
  wire  _GEN_278 = 10'hfe == array_addr[14:5] ? valid_254 : _GEN_277; // @[DCache.scala 78:{33,33}]
  wire  _GEN_279 = 10'hff == array_addr[14:5] ? valid_255 : _GEN_278; // @[DCache.scala 78:{33,33}]
  wire  _GEN_280 = 10'h100 == array_addr[14:5] ? valid_256 : _GEN_279; // @[DCache.scala 78:{33,33}]
  wire  _GEN_281 = 10'h101 == array_addr[14:5] ? valid_257 : _GEN_280; // @[DCache.scala 78:{33,33}]
  wire  _GEN_282 = 10'h102 == array_addr[14:5] ? valid_258 : _GEN_281; // @[DCache.scala 78:{33,33}]
  wire  _GEN_283 = 10'h103 == array_addr[14:5] ? valid_259 : _GEN_282; // @[DCache.scala 78:{33,33}]
  wire  _GEN_284 = 10'h104 == array_addr[14:5] ? valid_260 : _GEN_283; // @[DCache.scala 78:{33,33}]
  wire  _GEN_285 = 10'h105 == array_addr[14:5] ? valid_261 : _GEN_284; // @[DCache.scala 78:{33,33}]
  wire  _GEN_286 = 10'h106 == array_addr[14:5] ? valid_262 : _GEN_285; // @[DCache.scala 78:{33,33}]
  wire  _GEN_287 = 10'h107 == array_addr[14:5] ? valid_263 : _GEN_286; // @[DCache.scala 78:{33,33}]
  wire  _GEN_288 = 10'h108 == array_addr[14:5] ? valid_264 : _GEN_287; // @[DCache.scala 78:{33,33}]
  wire  _GEN_289 = 10'h109 == array_addr[14:5] ? valid_265 : _GEN_288; // @[DCache.scala 78:{33,33}]
  wire  _GEN_290 = 10'h10a == array_addr[14:5] ? valid_266 : _GEN_289; // @[DCache.scala 78:{33,33}]
  wire  _GEN_291 = 10'h10b == array_addr[14:5] ? valid_267 : _GEN_290; // @[DCache.scala 78:{33,33}]
  wire  _GEN_292 = 10'h10c == array_addr[14:5] ? valid_268 : _GEN_291; // @[DCache.scala 78:{33,33}]
  wire  _GEN_293 = 10'h10d == array_addr[14:5] ? valid_269 : _GEN_292; // @[DCache.scala 78:{33,33}]
  wire  _GEN_294 = 10'h10e == array_addr[14:5] ? valid_270 : _GEN_293; // @[DCache.scala 78:{33,33}]
  wire  _GEN_295 = 10'h10f == array_addr[14:5] ? valid_271 : _GEN_294; // @[DCache.scala 78:{33,33}]
  wire  _GEN_296 = 10'h110 == array_addr[14:5] ? valid_272 : _GEN_295; // @[DCache.scala 78:{33,33}]
  wire  _GEN_297 = 10'h111 == array_addr[14:5] ? valid_273 : _GEN_296; // @[DCache.scala 78:{33,33}]
  wire  _GEN_298 = 10'h112 == array_addr[14:5] ? valid_274 : _GEN_297; // @[DCache.scala 78:{33,33}]
  wire  _GEN_299 = 10'h113 == array_addr[14:5] ? valid_275 : _GEN_298; // @[DCache.scala 78:{33,33}]
  wire  _GEN_300 = 10'h114 == array_addr[14:5] ? valid_276 : _GEN_299; // @[DCache.scala 78:{33,33}]
  wire  _GEN_301 = 10'h115 == array_addr[14:5] ? valid_277 : _GEN_300; // @[DCache.scala 78:{33,33}]
  wire  _GEN_302 = 10'h116 == array_addr[14:5] ? valid_278 : _GEN_301; // @[DCache.scala 78:{33,33}]
  wire  _GEN_303 = 10'h117 == array_addr[14:5] ? valid_279 : _GEN_302; // @[DCache.scala 78:{33,33}]
  wire  _GEN_304 = 10'h118 == array_addr[14:5] ? valid_280 : _GEN_303; // @[DCache.scala 78:{33,33}]
  wire  _GEN_305 = 10'h119 == array_addr[14:5] ? valid_281 : _GEN_304; // @[DCache.scala 78:{33,33}]
  wire  _GEN_306 = 10'h11a == array_addr[14:5] ? valid_282 : _GEN_305; // @[DCache.scala 78:{33,33}]
  wire  _GEN_307 = 10'h11b == array_addr[14:5] ? valid_283 : _GEN_306; // @[DCache.scala 78:{33,33}]
  wire  _GEN_308 = 10'h11c == array_addr[14:5] ? valid_284 : _GEN_307; // @[DCache.scala 78:{33,33}]
  wire  _GEN_309 = 10'h11d == array_addr[14:5] ? valid_285 : _GEN_308; // @[DCache.scala 78:{33,33}]
  wire  _GEN_310 = 10'h11e == array_addr[14:5] ? valid_286 : _GEN_309; // @[DCache.scala 78:{33,33}]
  wire  _GEN_311 = 10'h11f == array_addr[14:5] ? valid_287 : _GEN_310; // @[DCache.scala 78:{33,33}]
  wire  _GEN_312 = 10'h120 == array_addr[14:5] ? valid_288 : _GEN_311; // @[DCache.scala 78:{33,33}]
  wire  _GEN_313 = 10'h121 == array_addr[14:5] ? valid_289 : _GEN_312; // @[DCache.scala 78:{33,33}]
  wire  _GEN_314 = 10'h122 == array_addr[14:5] ? valid_290 : _GEN_313; // @[DCache.scala 78:{33,33}]
  wire  _GEN_315 = 10'h123 == array_addr[14:5] ? valid_291 : _GEN_314; // @[DCache.scala 78:{33,33}]
  wire  _GEN_316 = 10'h124 == array_addr[14:5] ? valid_292 : _GEN_315; // @[DCache.scala 78:{33,33}]
  wire  _GEN_317 = 10'h125 == array_addr[14:5] ? valid_293 : _GEN_316; // @[DCache.scala 78:{33,33}]
  wire  _GEN_318 = 10'h126 == array_addr[14:5] ? valid_294 : _GEN_317; // @[DCache.scala 78:{33,33}]
  wire  _GEN_319 = 10'h127 == array_addr[14:5] ? valid_295 : _GEN_318; // @[DCache.scala 78:{33,33}]
  wire  _GEN_320 = 10'h128 == array_addr[14:5] ? valid_296 : _GEN_319; // @[DCache.scala 78:{33,33}]
  wire  _GEN_321 = 10'h129 == array_addr[14:5] ? valid_297 : _GEN_320; // @[DCache.scala 78:{33,33}]
  wire  _GEN_322 = 10'h12a == array_addr[14:5] ? valid_298 : _GEN_321; // @[DCache.scala 78:{33,33}]
  wire  _GEN_323 = 10'h12b == array_addr[14:5] ? valid_299 : _GEN_322; // @[DCache.scala 78:{33,33}]
  wire  _GEN_324 = 10'h12c == array_addr[14:5] ? valid_300 : _GEN_323; // @[DCache.scala 78:{33,33}]
  wire  _GEN_325 = 10'h12d == array_addr[14:5] ? valid_301 : _GEN_324; // @[DCache.scala 78:{33,33}]
  wire  _GEN_326 = 10'h12e == array_addr[14:5] ? valid_302 : _GEN_325; // @[DCache.scala 78:{33,33}]
  wire  _GEN_327 = 10'h12f == array_addr[14:5] ? valid_303 : _GEN_326; // @[DCache.scala 78:{33,33}]
  wire  _GEN_328 = 10'h130 == array_addr[14:5] ? valid_304 : _GEN_327; // @[DCache.scala 78:{33,33}]
  wire  _GEN_329 = 10'h131 == array_addr[14:5] ? valid_305 : _GEN_328; // @[DCache.scala 78:{33,33}]
  wire  _GEN_330 = 10'h132 == array_addr[14:5] ? valid_306 : _GEN_329; // @[DCache.scala 78:{33,33}]
  wire  _GEN_331 = 10'h133 == array_addr[14:5] ? valid_307 : _GEN_330; // @[DCache.scala 78:{33,33}]
  wire  _GEN_332 = 10'h134 == array_addr[14:5] ? valid_308 : _GEN_331; // @[DCache.scala 78:{33,33}]
  wire  _GEN_333 = 10'h135 == array_addr[14:5] ? valid_309 : _GEN_332; // @[DCache.scala 78:{33,33}]
  wire  _GEN_334 = 10'h136 == array_addr[14:5] ? valid_310 : _GEN_333; // @[DCache.scala 78:{33,33}]
  wire  _GEN_335 = 10'h137 == array_addr[14:5] ? valid_311 : _GEN_334; // @[DCache.scala 78:{33,33}]
  wire  _GEN_336 = 10'h138 == array_addr[14:5] ? valid_312 : _GEN_335; // @[DCache.scala 78:{33,33}]
  wire  _GEN_337 = 10'h139 == array_addr[14:5] ? valid_313 : _GEN_336; // @[DCache.scala 78:{33,33}]
  wire  _GEN_338 = 10'h13a == array_addr[14:5] ? valid_314 : _GEN_337; // @[DCache.scala 78:{33,33}]
  wire  _GEN_339 = 10'h13b == array_addr[14:5] ? valid_315 : _GEN_338; // @[DCache.scala 78:{33,33}]
  wire  _GEN_340 = 10'h13c == array_addr[14:5] ? valid_316 : _GEN_339; // @[DCache.scala 78:{33,33}]
  wire  _GEN_341 = 10'h13d == array_addr[14:5] ? valid_317 : _GEN_340; // @[DCache.scala 78:{33,33}]
  wire  _GEN_342 = 10'h13e == array_addr[14:5] ? valid_318 : _GEN_341; // @[DCache.scala 78:{33,33}]
  wire  _GEN_343 = 10'h13f == array_addr[14:5] ? valid_319 : _GEN_342; // @[DCache.scala 78:{33,33}]
  wire  _GEN_344 = 10'h140 == array_addr[14:5] ? valid_320 : _GEN_343; // @[DCache.scala 78:{33,33}]
  wire  _GEN_345 = 10'h141 == array_addr[14:5] ? valid_321 : _GEN_344; // @[DCache.scala 78:{33,33}]
  wire  _GEN_346 = 10'h142 == array_addr[14:5] ? valid_322 : _GEN_345; // @[DCache.scala 78:{33,33}]
  wire  _GEN_347 = 10'h143 == array_addr[14:5] ? valid_323 : _GEN_346; // @[DCache.scala 78:{33,33}]
  wire  _GEN_348 = 10'h144 == array_addr[14:5] ? valid_324 : _GEN_347; // @[DCache.scala 78:{33,33}]
  wire  _GEN_349 = 10'h145 == array_addr[14:5] ? valid_325 : _GEN_348; // @[DCache.scala 78:{33,33}]
  wire  _GEN_350 = 10'h146 == array_addr[14:5] ? valid_326 : _GEN_349; // @[DCache.scala 78:{33,33}]
  wire  _GEN_351 = 10'h147 == array_addr[14:5] ? valid_327 : _GEN_350; // @[DCache.scala 78:{33,33}]
  wire  _GEN_352 = 10'h148 == array_addr[14:5] ? valid_328 : _GEN_351; // @[DCache.scala 78:{33,33}]
  wire  _GEN_353 = 10'h149 == array_addr[14:5] ? valid_329 : _GEN_352; // @[DCache.scala 78:{33,33}]
  wire  _GEN_354 = 10'h14a == array_addr[14:5] ? valid_330 : _GEN_353; // @[DCache.scala 78:{33,33}]
  wire  _GEN_355 = 10'h14b == array_addr[14:5] ? valid_331 : _GEN_354; // @[DCache.scala 78:{33,33}]
  wire  _GEN_356 = 10'h14c == array_addr[14:5] ? valid_332 : _GEN_355; // @[DCache.scala 78:{33,33}]
  wire  _GEN_357 = 10'h14d == array_addr[14:5] ? valid_333 : _GEN_356; // @[DCache.scala 78:{33,33}]
  wire  _GEN_358 = 10'h14e == array_addr[14:5] ? valid_334 : _GEN_357; // @[DCache.scala 78:{33,33}]
  wire  _GEN_359 = 10'h14f == array_addr[14:5] ? valid_335 : _GEN_358; // @[DCache.scala 78:{33,33}]
  wire  _GEN_360 = 10'h150 == array_addr[14:5] ? valid_336 : _GEN_359; // @[DCache.scala 78:{33,33}]
  wire  _GEN_361 = 10'h151 == array_addr[14:5] ? valid_337 : _GEN_360; // @[DCache.scala 78:{33,33}]
  wire  _GEN_362 = 10'h152 == array_addr[14:5] ? valid_338 : _GEN_361; // @[DCache.scala 78:{33,33}]
  wire  _GEN_363 = 10'h153 == array_addr[14:5] ? valid_339 : _GEN_362; // @[DCache.scala 78:{33,33}]
  wire  _GEN_364 = 10'h154 == array_addr[14:5] ? valid_340 : _GEN_363; // @[DCache.scala 78:{33,33}]
  wire  _GEN_365 = 10'h155 == array_addr[14:5] ? valid_341 : _GEN_364; // @[DCache.scala 78:{33,33}]
  wire  _GEN_366 = 10'h156 == array_addr[14:5] ? valid_342 : _GEN_365; // @[DCache.scala 78:{33,33}]
  wire  _GEN_367 = 10'h157 == array_addr[14:5] ? valid_343 : _GEN_366; // @[DCache.scala 78:{33,33}]
  wire  _GEN_368 = 10'h158 == array_addr[14:5] ? valid_344 : _GEN_367; // @[DCache.scala 78:{33,33}]
  wire  _GEN_369 = 10'h159 == array_addr[14:5] ? valid_345 : _GEN_368; // @[DCache.scala 78:{33,33}]
  wire  _GEN_370 = 10'h15a == array_addr[14:5] ? valid_346 : _GEN_369; // @[DCache.scala 78:{33,33}]
  wire  _GEN_371 = 10'h15b == array_addr[14:5] ? valid_347 : _GEN_370; // @[DCache.scala 78:{33,33}]
  wire  _GEN_372 = 10'h15c == array_addr[14:5] ? valid_348 : _GEN_371; // @[DCache.scala 78:{33,33}]
  wire  _GEN_373 = 10'h15d == array_addr[14:5] ? valid_349 : _GEN_372; // @[DCache.scala 78:{33,33}]
  wire  _GEN_374 = 10'h15e == array_addr[14:5] ? valid_350 : _GEN_373; // @[DCache.scala 78:{33,33}]
  wire  _GEN_375 = 10'h15f == array_addr[14:5] ? valid_351 : _GEN_374; // @[DCache.scala 78:{33,33}]
  wire  _GEN_376 = 10'h160 == array_addr[14:5] ? valid_352 : _GEN_375; // @[DCache.scala 78:{33,33}]
  wire  _GEN_377 = 10'h161 == array_addr[14:5] ? valid_353 : _GEN_376; // @[DCache.scala 78:{33,33}]
  wire  _GEN_378 = 10'h162 == array_addr[14:5] ? valid_354 : _GEN_377; // @[DCache.scala 78:{33,33}]
  wire  _GEN_379 = 10'h163 == array_addr[14:5] ? valid_355 : _GEN_378; // @[DCache.scala 78:{33,33}]
  wire  _GEN_380 = 10'h164 == array_addr[14:5] ? valid_356 : _GEN_379; // @[DCache.scala 78:{33,33}]
  wire  _GEN_381 = 10'h165 == array_addr[14:5] ? valid_357 : _GEN_380; // @[DCache.scala 78:{33,33}]
  wire  _GEN_382 = 10'h166 == array_addr[14:5] ? valid_358 : _GEN_381; // @[DCache.scala 78:{33,33}]
  wire  _GEN_383 = 10'h167 == array_addr[14:5] ? valid_359 : _GEN_382; // @[DCache.scala 78:{33,33}]
  wire  _GEN_384 = 10'h168 == array_addr[14:5] ? valid_360 : _GEN_383; // @[DCache.scala 78:{33,33}]
  wire  _GEN_385 = 10'h169 == array_addr[14:5] ? valid_361 : _GEN_384; // @[DCache.scala 78:{33,33}]
  wire  _GEN_386 = 10'h16a == array_addr[14:5] ? valid_362 : _GEN_385; // @[DCache.scala 78:{33,33}]
  wire  _GEN_387 = 10'h16b == array_addr[14:5] ? valid_363 : _GEN_386; // @[DCache.scala 78:{33,33}]
  wire  _GEN_388 = 10'h16c == array_addr[14:5] ? valid_364 : _GEN_387; // @[DCache.scala 78:{33,33}]
  wire  _GEN_389 = 10'h16d == array_addr[14:5] ? valid_365 : _GEN_388; // @[DCache.scala 78:{33,33}]
  wire  _GEN_390 = 10'h16e == array_addr[14:5] ? valid_366 : _GEN_389; // @[DCache.scala 78:{33,33}]
  wire  _GEN_391 = 10'h16f == array_addr[14:5] ? valid_367 : _GEN_390; // @[DCache.scala 78:{33,33}]
  wire  _GEN_392 = 10'h170 == array_addr[14:5] ? valid_368 : _GEN_391; // @[DCache.scala 78:{33,33}]
  wire  _GEN_393 = 10'h171 == array_addr[14:5] ? valid_369 : _GEN_392; // @[DCache.scala 78:{33,33}]
  wire  _GEN_394 = 10'h172 == array_addr[14:5] ? valid_370 : _GEN_393; // @[DCache.scala 78:{33,33}]
  wire  _GEN_395 = 10'h173 == array_addr[14:5] ? valid_371 : _GEN_394; // @[DCache.scala 78:{33,33}]
  wire  _GEN_396 = 10'h174 == array_addr[14:5] ? valid_372 : _GEN_395; // @[DCache.scala 78:{33,33}]
  wire  _GEN_397 = 10'h175 == array_addr[14:5] ? valid_373 : _GEN_396; // @[DCache.scala 78:{33,33}]
  wire  _GEN_398 = 10'h176 == array_addr[14:5] ? valid_374 : _GEN_397; // @[DCache.scala 78:{33,33}]
  wire  _GEN_399 = 10'h177 == array_addr[14:5] ? valid_375 : _GEN_398; // @[DCache.scala 78:{33,33}]
  wire  _GEN_400 = 10'h178 == array_addr[14:5] ? valid_376 : _GEN_399; // @[DCache.scala 78:{33,33}]
  wire  _GEN_401 = 10'h179 == array_addr[14:5] ? valid_377 : _GEN_400; // @[DCache.scala 78:{33,33}]
  wire  _GEN_402 = 10'h17a == array_addr[14:5] ? valid_378 : _GEN_401; // @[DCache.scala 78:{33,33}]
  wire  _GEN_403 = 10'h17b == array_addr[14:5] ? valid_379 : _GEN_402; // @[DCache.scala 78:{33,33}]
  wire  _GEN_404 = 10'h17c == array_addr[14:5] ? valid_380 : _GEN_403; // @[DCache.scala 78:{33,33}]
  wire  _GEN_405 = 10'h17d == array_addr[14:5] ? valid_381 : _GEN_404; // @[DCache.scala 78:{33,33}]
  wire  _GEN_406 = 10'h17e == array_addr[14:5] ? valid_382 : _GEN_405; // @[DCache.scala 78:{33,33}]
  wire  _GEN_407 = 10'h17f == array_addr[14:5] ? valid_383 : _GEN_406; // @[DCache.scala 78:{33,33}]
  wire  _GEN_408 = 10'h180 == array_addr[14:5] ? valid_384 : _GEN_407; // @[DCache.scala 78:{33,33}]
  wire  _GEN_409 = 10'h181 == array_addr[14:5] ? valid_385 : _GEN_408; // @[DCache.scala 78:{33,33}]
  wire  _GEN_410 = 10'h182 == array_addr[14:5] ? valid_386 : _GEN_409; // @[DCache.scala 78:{33,33}]
  wire  _GEN_411 = 10'h183 == array_addr[14:5] ? valid_387 : _GEN_410; // @[DCache.scala 78:{33,33}]
  wire  _GEN_412 = 10'h184 == array_addr[14:5] ? valid_388 : _GEN_411; // @[DCache.scala 78:{33,33}]
  wire  _GEN_413 = 10'h185 == array_addr[14:5] ? valid_389 : _GEN_412; // @[DCache.scala 78:{33,33}]
  wire  _GEN_414 = 10'h186 == array_addr[14:5] ? valid_390 : _GEN_413; // @[DCache.scala 78:{33,33}]
  wire  _GEN_415 = 10'h187 == array_addr[14:5] ? valid_391 : _GEN_414; // @[DCache.scala 78:{33,33}]
  wire  _GEN_416 = 10'h188 == array_addr[14:5] ? valid_392 : _GEN_415; // @[DCache.scala 78:{33,33}]
  wire  _GEN_417 = 10'h189 == array_addr[14:5] ? valid_393 : _GEN_416; // @[DCache.scala 78:{33,33}]
  wire  _GEN_418 = 10'h18a == array_addr[14:5] ? valid_394 : _GEN_417; // @[DCache.scala 78:{33,33}]
  wire  _GEN_419 = 10'h18b == array_addr[14:5] ? valid_395 : _GEN_418; // @[DCache.scala 78:{33,33}]
  wire  _GEN_420 = 10'h18c == array_addr[14:5] ? valid_396 : _GEN_419; // @[DCache.scala 78:{33,33}]
  wire  _GEN_421 = 10'h18d == array_addr[14:5] ? valid_397 : _GEN_420; // @[DCache.scala 78:{33,33}]
  wire  _GEN_422 = 10'h18e == array_addr[14:5] ? valid_398 : _GEN_421; // @[DCache.scala 78:{33,33}]
  wire  _GEN_423 = 10'h18f == array_addr[14:5] ? valid_399 : _GEN_422; // @[DCache.scala 78:{33,33}]
  wire  _GEN_424 = 10'h190 == array_addr[14:5] ? valid_400 : _GEN_423; // @[DCache.scala 78:{33,33}]
  wire  _GEN_425 = 10'h191 == array_addr[14:5] ? valid_401 : _GEN_424; // @[DCache.scala 78:{33,33}]
  wire  _GEN_426 = 10'h192 == array_addr[14:5] ? valid_402 : _GEN_425; // @[DCache.scala 78:{33,33}]
  wire  _GEN_427 = 10'h193 == array_addr[14:5] ? valid_403 : _GEN_426; // @[DCache.scala 78:{33,33}]
  wire  _GEN_428 = 10'h194 == array_addr[14:5] ? valid_404 : _GEN_427; // @[DCache.scala 78:{33,33}]
  wire  _GEN_429 = 10'h195 == array_addr[14:5] ? valid_405 : _GEN_428; // @[DCache.scala 78:{33,33}]
  wire  _GEN_430 = 10'h196 == array_addr[14:5] ? valid_406 : _GEN_429; // @[DCache.scala 78:{33,33}]
  wire  _GEN_431 = 10'h197 == array_addr[14:5] ? valid_407 : _GEN_430; // @[DCache.scala 78:{33,33}]
  wire  _GEN_432 = 10'h198 == array_addr[14:5] ? valid_408 : _GEN_431; // @[DCache.scala 78:{33,33}]
  wire  _GEN_433 = 10'h199 == array_addr[14:5] ? valid_409 : _GEN_432; // @[DCache.scala 78:{33,33}]
  wire  _GEN_434 = 10'h19a == array_addr[14:5] ? valid_410 : _GEN_433; // @[DCache.scala 78:{33,33}]
  wire  _GEN_435 = 10'h19b == array_addr[14:5] ? valid_411 : _GEN_434; // @[DCache.scala 78:{33,33}]
  wire  _GEN_436 = 10'h19c == array_addr[14:5] ? valid_412 : _GEN_435; // @[DCache.scala 78:{33,33}]
  wire  _GEN_437 = 10'h19d == array_addr[14:5] ? valid_413 : _GEN_436; // @[DCache.scala 78:{33,33}]
  wire  _GEN_438 = 10'h19e == array_addr[14:5] ? valid_414 : _GEN_437; // @[DCache.scala 78:{33,33}]
  wire  _GEN_439 = 10'h19f == array_addr[14:5] ? valid_415 : _GEN_438; // @[DCache.scala 78:{33,33}]
  wire  _GEN_440 = 10'h1a0 == array_addr[14:5] ? valid_416 : _GEN_439; // @[DCache.scala 78:{33,33}]
  wire  _GEN_441 = 10'h1a1 == array_addr[14:5] ? valid_417 : _GEN_440; // @[DCache.scala 78:{33,33}]
  wire  _GEN_442 = 10'h1a2 == array_addr[14:5] ? valid_418 : _GEN_441; // @[DCache.scala 78:{33,33}]
  wire  _GEN_443 = 10'h1a3 == array_addr[14:5] ? valid_419 : _GEN_442; // @[DCache.scala 78:{33,33}]
  wire  _GEN_444 = 10'h1a4 == array_addr[14:5] ? valid_420 : _GEN_443; // @[DCache.scala 78:{33,33}]
  wire  _GEN_445 = 10'h1a5 == array_addr[14:5] ? valid_421 : _GEN_444; // @[DCache.scala 78:{33,33}]
  wire  _GEN_446 = 10'h1a6 == array_addr[14:5] ? valid_422 : _GEN_445; // @[DCache.scala 78:{33,33}]
  wire  _GEN_447 = 10'h1a7 == array_addr[14:5] ? valid_423 : _GEN_446; // @[DCache.scala 78:{33,33}]
  wire  _GEN_448 = 10'h1a8 == array_addr[14:5] ? valid_424 : _GEN_447; // @[DCache.scala 78:{33,33}]
  wire  _GEN_449 = 10'h1a9 == array_addr[14:5] ? valid_425 : _GEN_448; // @[DCache.scala 78:{33,33}]
  wire  _GEN_450 = 10'h1aa == array_addr[14:5] ? valid_426 : _GEN_449; // @[DCache.scala 78:{33,33}]
  wire  _GEN_451 = 10'h1ab == array_addr[14:5] ? valid_427 : _GEN_450; // @[DCache.scala 78:{33,33}]
  wire  _GEN_452 = 10'h1ac == array_addr[14:5] ? valid_428 : _GEN_451; // @[DCache.scala 78:{33,33}]
  wire  _GEN_453 = 10'h1ad == array_addr[14:5] ? valid_429 : _GEN_452; // @[DCache.scala 78:{33,33}]
  wire  _GEN_454 = 10'h1ae == array_addr[14:5] ? valid_430 : _GEN_453; // @[DCache.scala 78:{33,33}]
  wire  _GEN_455 = 10'h1af == array_addr[14:5] ? valid_431 : _GEN_454; // @[DCache.scala 78:{33,33}]
  wire  _GEN_456 = 10'h1b0 == array_addr[14:5] ? valid_432 : _GEN_455; // @[DCache.scala 78:{33,33}]
  wire  _GEN_457 = 10'h1b1 == array_addr[14:5] ? valid_433 : _GEN_456; // @[DCache.scala 78:{33,33}]
  wire  _GEN_458 = 10'h1b2 == array_addr[14:5] ? valid_434 : _GEN_457; // @[DCache.scala 78:{33,33}]
  wire  _GEN_459 = 10'h1b3 == array_addr[14:5] ? valid_435 : _GEN_458; // @[DCache.scala 78:{33,33}]
  wire  _GEN_460 = 10'h1b4 == array_addr[14:5] ? valid_436 : _GEN_459; // @[DCache.scala 78:{33,33}]
  wire  _GEN_461 = 10'h1b5 == array_addr[14:5] ? valid_437 : _GEN_460; // @[DCache.scala 78:{33,33}]
  wire  _GEN_462 = 10'h1b6 == array_addr[14:5] ? valid_438 : _GEN_461; // @[DCache.scala 78:{33,33}]
  wire  _GEN_463 = 10'h1b7 == array_addr[14:5] ? valid_439 : _GEN_462; // @[DCache.scala 78:{33,33}]
  wire  _GEN_464 = 10'h1b8 == array_addr[14:5] ? valid_440 : _GEN_463; // @[DCache.scala 78:{33,33}]
  wire  _GEN_465 = 10'h1b9 == array_addr[14:5] ? valid_441 : _GEN_464; // @[DCache.scala 78:{33,33}]
  wire  _GEN_466 = 10'h1ba == array_addr[14:5] ? valid_442 : _GEN_465; // @[DCache.scala 78:{33,33}]
  wire  _GEN_467 = 10'h1bb == array_addr[14:5] ? valid_443 : _GEN_466; // @[DCache.scala 78:{33,33}]
  wire  _GEN_468 = 10'h1bc == array_addr[14:5] ? valid_444 : _GEN_467; // @[DCache.scala 78:{33,33}]
  wire  _GEN_469 = 10'h1bd == array_addr[14:5] ? valid_445 : _GEN_468; // @[DCache.scala 78:{33,33}]
  wire  _GEN_470 = 10'h1be == array_addr[14:5] ? valid_446 : _GEN_469; // @[DCache.scala 78:{33,33}]
  wire  _GEN_471 = 10'h1bf == array_addr[14:5] ? valid_447 : _GEN_470; // @[DCache.scala 78:{33,33}]
  wire  _GEN_472 = 10'h1c0 == array_addr[14:5] ? valid_448 : _GEN_471; // @[DCache.scala 78:{33,33}]
  wire  _GEN_473 = 10'h1c1 == array_addr[14:5] ? valid_449 : _GEN_472; // @[DCache.scala 78:{33,33}]
  wire  _GEN_474 = 10'h1c2 == array_addr[14:5] ? valid_450 : _GEN_473; // @[DCache.scala 78:{33,33}]
  wire  _GEN_475 = 10'h1c3 == array_addr[14:5] ? valid_451 : _GEN_474; // @[DCache.scala 78:{33,33}]
  wire  _GEN_476 = 10'h1c4 == array_addr[14:5] ? valid_452 : _GEN_475; // @[DCache.scala 78:{33,33}]
  wire  _GEN_477 = 10'h1c5 == array_addr[14:5] ? valid_453 : _GEN_476; // @[DCache.scala 78:{33,33}]
  wire  _GEN_478 = 10'h1c6 == array_addr[14:5] ? valid_454 : _GEN_477; // @[DCache.scala 78:{33,33}]
  wire  _GEN_479 = 10'h1c7 == array_addr[14:5] ? valid_455 : _GEN_478; // @[DCache.scala 78:{33,33}]
  wire  _GEN_480 = 10'h1c8 == array_addr[14:5] ? valid_456 : _GEN_479; // @[DCache.scala 78:{33,33}]
  wire  _GEN_481 = 10'h1c9 == array_addr[14:5] ? valid_457 : _GEN_480; // @[DCache.scala 78:{33,33}]
  wire  _GEN_482 = 10'h1ca == array_addr[14:5] ? valid_458 : _GEN_481; // @[DCache.scala 78:{33,33}]
  wire  _GEN_483 = 10'h1cb == array_addr[14:5] ? valid_459 : _GEN_482; // @[DCache.scala 78:{33,33}]
  wire  _GEN_484 = 10'h1cc == array_addr[14:5] ? valid_460 : _GEN_483; // @[DCache.scala 78:{33,33}]
  wire  _GEN_485 = 10'h1cd == array_addr[14:5] ? valid_461 : _GEN_484; // @[DCache.scala 78:{33,33}]
  wire  _GEN_486 = 10'h1ce == array_addr[14:5] ? valid_462 : _GEN_485; // @[DCache.scala 78:{33,33}]
  wire  _GEN_487 = 10'h1cf == array_addr[14:5] ? valid_463 : _GEN_486; // @[DCache.scala 78:{33,33}]
  wire  _GEN_488 = 10'h1d0 == array_addr[14:5] ? valid_464 : _GEN_487; // @[DCache.scala 78:{33,33}]
  wire  _GEN_489 = 10'h1d1 == array_addr[14:5] ? valid_465 : _GEN_488; // @[DCache.scala 78:{33,33}]
  wire  _GEN_490 = 10'h1d2 == array_addr[14:5] ? valid_466 : _GEN_489; // @[DCache.scala 78:{33,33}]
  wire  _GEN_491 = 10'h1d3 == array_addr[14:5] ? valid_467 : _GEN_490; // @[DCache.scala 78:{33,33}]
  wire  _GEN_492 = 10'h1d4 == array_addr[14:5] ? valid_468 : _GEN_491; // @[DCache.scala 78:{33,33}]
  wire  _GEN_493 = 10'h1d5 == array_addr[14:5] ? valid_469 : _GEN_492; // @[DCache.scala 78:{33,33}]
  wire  _GEN_494 = 10'h1d6 == array_addr[14:5] ? valid_470 : _GEN_493; // @[DCache.scala 78:{33,33}]
  wire  _GEN_495 = 10'h1d7 == array_addr[14:5] ? valid_471 : _GEN_494; // @[DCache.scala 78:{33,33}]
  wire  _GEN_496 = 10'h1d8 == array_addr[14:5] ? valid_472 : _GEN_495; // @[DCache.scala 78:{33,33}]
  wire  _GEN_497 = 10'h1d9 == array_addr[14:5] ? valid_473 : _GEN_496; // @[DCache.scala 78:{33,33}]
  wire  _GEN_498 = 10'h1da == array_addr[14:5] ? valid_474 : _GEN_497; // @[DCache.scala 78:{33,33}]
  wire  _GEN_499 = 10'h1db == array_addr[14:5] ? valid_475 : _GEN_498; // @[DCache.scala 78:{33,33}]
  wire  _GEN_500 = 10'h1dc == array_addr[14:5] ? valid_476 : _GEN_499; // @[DCache.scala 78:{33,33}]
  wire  _GEN_501 = 10'h1dd == array_addr[14:5] ? valid_477 : _GEN_500; // @[DCache.scala 78:{33,33}]
  wire  _GEN_502 = 10'h1de == array_addr[14:5] ? valid_478 : _GEN_501; // @[DCache.scala 78:{33,33}]
  wire  _GEN_503 = 10'h1df == array_addr[14:5] ? valid_479 : _GEN_502; // @[DCache.scala 78:{33,33}]
  wire  _GEN_504 = 10'h1e0 == array_addr[14:5] ? valid_480 : _GEN_503; // @[DCache.scala 78:{33,33}]
  wire  _GEN_505 = 10'h1e1 == array_addr[14:5] ? valid_481 : _GEN_504; // @[DCache.scala 78:{33,33}]
  wire  _GEN_506 = 10'h1e2 == array_addr[14:5] ? valid_482 : _GEN_505; // @[DCache.scala 78:{33,33}]
  wire  _GEN_507 = 10'h1e3 == array_addr[14:5] ? valid_483 : _GEN_506; // @[DCache.scala 78:{33,33}]
  wire  _GEN_508 = 10'h1e4 == array_addr[14:5] ? valid_484 : _GEN_507; // @[DCache.scala 78:{33,33}]
  wire  _GEN_509 = 10'h1e5 == array_addr[14:5] ? valid_485 : _GEN_508; // @[DCache.scala 78:{33,33}]
  wire  _GEN_510 = 10'h1e6 == array_addr[14:5] ? valid_486 : _GEN_509; // @[DCache.scala 78:{33,33}]
  wire  _GEN_511 = 10'h1e7 == array_addr[14:5] ? valid_487 : _GEN_510; // @[DCache.scala 78:{33,33}]
  wire  _GEN_512 = 10'h1e8 == array_addr[14:5] ? valid_488 : _GEN_511; // @[DCache.scala 78:{33,33}]
  wire  _GEN_513 = 10'h1e9 == array_addr[14:5] ? valid_489 : _GEN_512; // @[DCache.scala 78:{33,33}]
  wire  _GEN_514 = 10'h1ea == array_addr[14:5] ? valid_490 : _GEN_513; // @[DCache.scala 78:{33,33}]
  wire  _GEN_515 = 10'h1eb == array_addr[14:5] ? valid_491 : _GEN_514; // @[DCache.scala 78:{33,33}]
  wire  _GEN_516 = 10'h1ec == array_addr[14:5] ? valid_492 : _GEN_515; // @[DCache.scala 78:{33,33}]
  wire  _GEN_517 = 10'h1ed == array_addr[14:5] ? valid_493 : _GEN_516; // @[DCache.scala 78:{33,33}]
  wire  _GEN_518 = 10'h1ee == array_addr[14:5] ? valid_494 : _GEN_517; // @[DCache.scala 78:{33,33}]
  wire  _GEN_519 = 10'h1ef == array_addr[14:5] ? valid_495 : _GEN_518; // @[DCache.scala 78:{33,33}]
  wire  _GEN_520 = 10'h1f0 == array_addr[14:5] ? valid_496 : _GEN_519; // @[DCache.scala 78:{33,33}]
  wire  _GEN_521 = 10'h1f1 == array_addr[14:5] ? valid_497 : _GEN_520; // @[DCache.scala 78:{33,33}]
  wire  _GEN_522 = 10'h1f2 == array_addr[14:5] ? valid_498 : _GEN_521; // @[DCache.scala 78:{33,33}]
  wire  _GEN_523 = 10'h1f3 == array_addr[14:5] ? valid_499 : _GEN_522; // @[DCache.scala 78:{33,33}]
  wire  _GEN_524 = 10'h1f4 == array_addr[14:5] ? valid_500 : _GEN_523; // @[DCache.scala 78:{33,33}]
  wire  _GEN_525 = 10'h1f5 == array_addr[14:5] ? valid_501 : _GEN_524; // @[DCache.scala 78:{33,33}]
  wire  _GEN_526 = 10'h1f6 == array_addr[14:5] ? valid_502 : _GEN_525; // @[DCache.scala 78:{33,33}]
  wire  _GEN_527 = 10'h1f7 == array_addr[14:5] ? valid_503 : _GEN_526; // @[DCache.scala 78:{33,33}]
  wire  _GEN_528 = 10'h1f8 == array_addr[14:5] ? valid_504 : _GEN_527; // @[DCache.scala 78:{33,33}]
  wire  _GEN_529 = 10'h1f9 == array_addr[14:5] ? valid_505 : _GEN_528; // @[DCache.scala 78:{33,33}]
  wire  _GEN_530 = 10'h1fa == array_addr[14:5] ? valid_506 : _GEN_529; // @[DCache.scala 78:{33,33}]
  wire  _GEN_531 = 10'h1fb == array_addr[14:5] ? valid_507 : _GEN_530; // @[DCache.scala 78:{33,33}]
  wire  _GEN_532 = 10'h1fc == array_addr[14:5] ? valid_508 : _GEN_531; // @[DCache.scala 78:{33,33}]
  wire  _GEN_533 = 10'h1fd == array_addr[14:5] ? valid_509 : _GEN_532; // @[DCache.scala 78:{33,33}]
  wire  _GEN_534 = 10'h1fe == array_addr[14:5] ? valid_510 : _GEN_533; // @[DCache.scala 78:{33,33}]
  wire  _GEN_535 = 10'h1ff == array_addr[14:5] ? valid_511 : _GEN_534; // @[DCache.scala 78:{33,33}]
  wire  _GEN_536 = 10'h200 == array_addr[14:5] ? valid_512 : _GEN_535; // @[DCache.scala 78:{33,33}]
  wire  _GEN_537 = 10'h201 == array_addr[14:5] ? valid_513 : _GEN_536; // @[DCache.scala 78:{33,33}]
  wire  _GEN_538 = 10'h202 == array_addr[14:5] ? valid_514 : _GEN_537; // @[DCache.scala 78:{33,33}]
  wire  _GEN_539 = 10'h203 == array_addr[14:5] ? valid_515 : _GEN_538; // @[DCache.scala 78:{33,33}]
  wire  _GEN_540 = 10'h204 == array_addr[14:5] ? valid_516 : _GEN_539; // @[DCache.scala 78:{33,33}]
  wire  _GEN_541 = 10'h205 == array_addr[14:5] ? valid_517 : _GEN_540; // @[DCache.scala 78:{33,33}]
  wire  _GEN_542 = 10'h206 == array_addr[14:5] ? valid_518 : _GEN_541; // @[DCache.scala 78:{33,33}]
  wire  _GEN_543 = 10'h207 == array_addr[14:5] ? valid_519 : _GEN_542; // @[DCache.scala 78:{33,33}]
  wire  _GEN_544 = 10'h208 == array_addr[14:5] ? valid_520 : _GEN_543; // @[DCache.scala 78:{33,33}]
  wire  _GEN_545 = 10'h209 == array_addr[14:5] ? valid_521 : _GEN_544; // @[DCache.scala 78:{33,33}]
  wire  _GEN_546 = 10'h20a == array_addr[14:5] ? valid_522 : _GEN_545; // @[DCache.scala 78:{33,33}]
  wire  _GEN_547 = 10'h20b == array_addr[14:5] ? valid_523 : _GEN_546; // @[DCache.scala 78:{33,33}]
  wire  _GEN_548 = 10'h20c == array_addr[14:5] ? valid_524 : _GEN_547; // @[DCache.scala 78:{33,33}]
  wire  _GEN_549 = 10'h20d == array_addr[14:5] ? valid_525 : _GEN_548; // @[DCache.scala 78:{33,33}]
  wire  _GEN_550 = 10'h20e == array_addr[14:5] ? valid_526 : _GEN_549; // @[DCache.scala 78:{33,33}]
  wire  _GEN_551 = 10'h20f == array_addr[14:5] ? valid_527 : _GEN_550; // @[DCache.scala 78:{33,33}]
  wire  _GEN_552 = 10'h210 == array_addr[14:5] ? valid_528 : _GEN_551; // @[DCache.scala 78:{33,33}]
  wire  _GEN_553 = 10'h211 == array_addr[14:5] ? valid_529 : _GEN_552; // @[DCache.scala 78:{33,33}]
  wire  _GEN_554 = 10'h212 == array_addr[14:5] ? valid_530 : _GEN_553; // @[DCache.scala 78:{33,33}]
  wire  _GEN_555 = 10'h213 == array_addr[14:5] ? valid_531 : _GEN_554; // @[DCache.scala 78:{33,33}]
  wire  _GEN_556 = 10'h214 == array_addr[14:5] ? valid_532 : _GEN_555; // @[DCache.scala 78:{33,33}]
  wire  _GEN_557 = 10'h215 == array_addr[14:5] ? valid_533 : _GEN_556; // @[DCache.scala 78:{33,33}]
  wire  _GEN_558 = 10'h216 == array_addr[14:5] ? valid_534 : _GEN_557; // @[DCache.scala 78:{33,33}]
  wire  _GEN_559 = 10'h217 == array_addr[14:5] ? valid_535 : _GEN_558; // @[DCache.scala 78:{33,33}]
  wire  _GEN_560 = 10'h218 == array_addr[14:5] ? valid_536 : _GEN_559; // @[DCache.scala 78:{33,33}]
  wire  _GEN_561 = 10'h219 == array_addr[14:5] ? valid_537 : _GEN_560; // @[DCache.scala 78:{33,33}]
  wire  _GEN_562 = 10'h21a == array_addr[14:5] ? valid_538 : _GEN_561; // @[DCache.scala 78:{33,33}]
  wire  _GEN_563 = 10'h21b == array_addr[14:5] ? valid_539 : _GEN_562; // @[DCache.scala 78:{33,33}]
  wire  _GEN_564 = 10'h21c == array_addr[14:5] ? valid_540 : _GEN_563; // @[DCache.scala 78:{33,33}]
  wire  _GEN_565 = 10'h21d == array_addr[14:5] ? valid_541 : _GEN_564; // @[DCache.scala 78:{33,33}]
  wire  _GEN_566 = 10'h21e == array_addr[14:5] ? valid_542 : _GEN_565; // @[DCache.scala 78:{33,33}]
  wire  _GEN_567 = 10'h21f == array_addr[14:5] ? valid_543 : _GEN_566; // @[DCache.scala 78:{33,33}]
  wire  _GEN_568 = 10'h220 == array_addr[14:5] ? valid_544 : _GEN_567; // @[DCache.scala 78:{33,33}]
  wire  _GEN_569 = 10'h221 == array_addr[14:5] ? valid_545 : _GEN_568; // @[DCache.scala 78:{33,33}]
  wire  _GEN_570 = 10'h222 == array_addr[14:5] ? valid_546 : _GEN_569; // @[DCache.scala 78:{33,33}]
  wire  _GEN_571 = 10'h223 == array_addr[14:5] ? valid_547 : _GEN_570; // @[DCache.scala 78:{33,33}]
  wire  _GEN_572 = 10'h224 == array_addr[14:5] ? valid_548 : _GEN_571; // @[DCache.scala 78:{33,33}]
  wire  _GEN_573 = 10'h225 == array_addr[14:5] ? valid_549 : _GEN_572; // @[DCache.scala 78:{33,33}]
  wire  _GEN_574 = 10'h226 == array_addr[14:5] ? valid_550 : _GEN_573; // @[DCache.scala 78:{33,33}]
  wire  _GEN_575 = 10'h227 == array_addr[14:5] ? valid_551 : _GEN_574; // @[DCache.scala 78:{33,33}]
  wire  _GEN_576 = 10'h228 == array_addr[14:5] ? valid_552 : _GEN_575; // @[DCache.scala 78:{33,33}]
  wire  _GEN_577 = 10'h229 == array_addr[14:5] ? valid_553 : _GEN_576; // @[DCache.scala 78:{33,33}]
  wire  _GEN_578 = 10'h22a == array_addr[14:5] ? valid_554 : _GEN_577; // @[DCache.scala 78:{33,33}]
  wire  _GEN_579 = 10'h22b == array_addr[14:5] ? valid_555 : _GEN_578; // @[DCache.scala 78:{33,33}]
  wire  _GEN_580 = 10'h22c == array_addr[14:5] ? valid_556 : _GEN_579; // @[DCache.scala 78:{33,33}]
  wire  _GEN_581 = 10'h22d == array_addr[14:5] ? valid_557 : _GEN_580; // @[DCache.scala 78:{33,33}]
  wire  _GEN_582 = 10'h22e == array_addr[14:5] ? valid_558 : _GEN_581; // @[DCache.scala 78:{33,33}]
  wire  _GEN_583 = 10'h22f == array_addr[14:5] ? valid_559 : _GEN_582; // @[DCache.scala 78:{33,33}]
  wire  _GEN_584 = 10'h230 == array_addr[14:5] ? valid_560 : _GEN_583; // @[DCache.scala 78:{33,33}]
  wire  _GEN_585 = 10'h231 == array_addr[14:5] ? valid_561 : _GEN_584; // @[DCache.scala 78:{33,33}]
  wire  _GEN_586 = 10'h232 == array_addr[14:5] ? valid_562 : _GEN_585; // @[DCache.scala 78:{33,33}]
  wire  _GEN_587 = 10'h233 == array_addr[14:5] ? valid_563 : _GEN_586; // @[DCache.scala 78:{33,33}]
  wire  _GEN_588 = 10'h234 == array_addr[14:5] ? valid_564 : _GEN_587; // @[DCache.scala 78:{33,33}]
  wire  _GEN_589 = 10'h235 == array_addr[14:5] ? valid_565 : _GEN_588; // @[DCache.scala 78:{33,33}]
  wire  _GEN_590 = 10'h236 == array_addr[14:5] ? valid_566 : _GEN_589; // @[DCache.scala 78:{33,33}]
  wire  _GEN_591 = 10'h237 == array_addr[14:5] ? valid_567 : _GEN_590; // @[DCache.scala 78:{33,33}]
  wire  _GEN_592 = 10'h238 == array_addr[14:5] ? valid_568 : _GEN_591; // @[DCache.scala 78:{33,33}]
  wire  _GEN_593 = 10'h239 == array_addr[14:5] ? valid_569 : _GEN_592; // @[DCache.scala 78:{33,33}]
  wire  _GEN_594 = 10'h23a == array_addr[14:5] ? valid_570 : _GEN_593; // @[DCache.scala 78:{33,33}]
  wire  _GEN_595 = 10'h23b == array_addr[14:5] ? valid_571 : _GEN_594; // @[DCache.scala 78:{33,33}]
  wire  _GEN_596 = 10'h23c == array_addr[14:5] ? valid_572 : _GEN_595; // @[DCache.scala 78:{33,33}]
  wire  _GEN_597 = 10'h23d == array_addr[14:5] ? valid_573 : _GEN_596; // @[DCache.scala 78:{33,33}]
  wire  _GEN_598 = 10'h23e == array_addr[14:5] ? valid_574 : _GEN_597; // @[DCache.scala 78:{33,33}]
  wire  _GEN_599 = 10'h23f == array_addr[14:5] ? valid_575 : _GEN_598; // @[DCache.scala 78:{33,33}]
  wire  _GEN_600 = 10'h240 == array_addr[14:5] ? valid_576 : _GEN_599; // @[DCache.scala 78:{33,33}]
  wire  _GEN_601 = 10'h241 == array_addr[14:5] ? valid_577 : _GEN_600; // @[DCache.scala 78:{33,33}]
  wire  _GEN_602 = 10'h242 == array_addr[14:5] ? valid_578 : _GEN_601; // @[DCache.scala 78:{33,33}]
  wire  _GEN_603 = 10'h243 == array_addr[14:5] ? valid_579 : _GEN_602; // @[DCache.scala 78:{33,33}]
  wire  _GEN_604 = 10'h244 == array_addr[14:5] ? valid_580 : _GEN_603; // @[DCache.scala 78:{33,33}]
  wire  _GEN_605 = 10'h245 == array_addr[14:5] ? valid_581 : _GEN_604; // @[DCache.scala 78:{33,33}]
  wire  _GEN_606 = 10'h246 == array_addr[14:5] ? valid_582 : _GEN_605; // @[DCache.scala 78:{33,33}]
  wire  _GEN_607 = 10'h247 == array_addr[14:5] ? valid_583 : _GEN_606; // @[DCache.scala 78:{33,33}]
  wire  _GEN_608 = 10'h248 == array_addr[14:5] ? valid_584 : _GEN_607; // @[DCache.scala 78:{33,33}]
  wire  _GEN_609 = 10'h249 == array_addr[14:5] ? valid_585 : _GEN_608; // @[DCache.scala 78:{33,33}]
  wire  _GEN_610 = 10'h24a == array_addr[14:5] ? valid_586 : _GEN_609; // @[DCache.scala 78:{33,33}]
  wire  _GEN_611 = 10'h24b == array_addr[14:5] ? valid_587 : _GEN_610; // @[DCache.scala 78:{33,33}]
  wire  _GEN_612 = 10'h24c == array_addr[14:5] ? valid_588 : _GEN_611; // @[DCache.scala 78:{33,33}]
  wire  _GEN_613 = 10'h24d == array_addr[14:5] ? valid_589 : _GEN_612; // @[DCache.scala 78:{33,33}]
  wire  _GEN_614 = 10'h24e == array_addr[14:5] ? valid_590 : _GEN_613; // @[DCache.scala 78:{33,33}]
  wire  _GEN_615 = 10'h24f == array_addr[14:5] ? valid_591 : _GEN_614; // @[DCache.scala 78:{33,33}]
  wire  _GEN_616 = 10'h250 == array_addr[14:5] ? valid_592 : _GEN_615; // @[DCache.scala 78:{33,33}]
  wire  _GEN_617 = 10'h251 == array_addr[14:5] ? valid_593 : _GEN_616; // @[DCache.scala 78:{33,33}]
  wire  _GEN_618 = 10'h252 == array_addr[14:5] ? valid_594 : _GEN_617; // @[DCache.scala 78:{33,33}]
  wire  _GEN_619 = 10'h253 == array_addr[14:5] ? valid_595 : _GEN_618; // @[DCache.scala 78:{33,33}]
  wire  _GEN_620 = 10'h254 == array_addr[14:5] ? valid_596 : _GEN_619; // @[DCache.scala 78:{33,33}]
  wire  _GEN_621 = 10'h255 == array_addr[14:5] ? valid_597 : _GEN_620; // @[DCache.scala 78:{33,33}]
  wire  _GEN_622 = 10'h256 == array_addr[14:5] ? valid_598 : _GEN_621; // @[DCache.scala 78:{33,33}]
  wire  _GEN_623 = 10'h257 == array_addr[14:5] ? valid_599 : _GEN_622; // @[DCache.scala 78:{33,33}]
  wire  _GEN_624 = 10'h258 == array_addr[14:5] ? valid_600 : _GEN_623; // @[DCache.scala 78:{33,33}]
  wire  _GEN_625 = 10'h259 == array_addr[14:5] ? valid_601 : _GEN_624; // @[DCache.scala 78:{33,33}]
  wire  _GEN_626 = 10'h25a == array_addr[14:5] ? valid_602 : _GEN_625; // @[DCache.scala 78:{33,33}]
  wire  _GEN_627 = 10'h25b == array_addr[14:5] ? valid_603 : _GEN_626; // @[DCache.scala 78:{33,33}]
  wire  _GEN_628 = 10'h25c == array_addr[14:5] ? valid_604 : _GEN_627; // @[DCache.scala 78:{33,33}]
  wire  _GEN_629 = 10'h25d == array_addr[14:5] ? valid_605 : _GEN_628; // @[DCache.scala 78:{33,33}]
  wire  _GEN_630 = 10'h25e == array_addr[14:5] ? valid_606 : _GEN_629; // @[DCache.scala 78:{33,33}]
  wire  _GEN_631 = 10'h25f == array_addr[14:5] ? valid_607 : _GEN_630; // @[DCache.scala 78:{33,33}]
  wire  _GEN_632 = 10'h260 == array_addr[14:5] ? valid_608 : _GEN_631; // @[DCache.scala 78:{33,33}]
  wire  _GEN_633 = 10'h261 == array_addr[14:5] ? valid_609 : _GEN_632; // @[DCache.scala 78:{33,33}]
  wire  _GEN_634 = 10'h262 == array_addr[14:5] ? valid_610 : _GEN_633; // @[DCache.scala 78:{33,33}]
  wire  _GEN_635 = 10'h263 == array_addr[14:5] ? valid_611 : _GEN_634; // @[DCache.scala 78:{33,33}]
  wire  _GEN_636 = 10'h264 == array_addr[14:5] ? valid_612 : _GEN_635; // @[DCache.scala 78:{33,33}]
  wire  _GEN_637 = 10'h265 == array_addr[14:5] ? valid_613 : _GEN_636; // @[DCache.scala 78:{33,33}]
  wire  _GEN_638 = 10'h266 == array_addr[14:5] ? valid_614 : _GEN_637; // @[DCache.scala 78:{33,33}]
  wire  _GEN_639 = 10'h267 == array_addr[14:5] ? valid_615 : _GEN_638; // @[DCache.scala 78:{33,33}]
  wire  _GEN_640 = 10'h268 == array_addr[14:5] ? valid_616 : _GEN_639; // @[DCache.scala 78:{33,33}]
  wire  _GEN_641 = 10'h269 == array_addr[14:5] ? valid_617 : _GEN_640; // @[DCache.scala 78:{33,33}]
  wire  _GEN_642 = 10'h26a == array_addr[14:5] ? valid_618 : _GEN_641; // @[DCache.scala 78:{33,33}]
  wire  _GEN_643 = 10'h26b == array_addr[14:5] ? valid_619 : _GEN_642; // @[DCache.scala 78:{33,33}]
  wire  _GEN_644 = 10'h26c == array_addr[14:5] ? valid_620 : _GEN_643; // @[DCache.scala 78:{33,33}]
  wire  _GEN_645 = 10'h26d == array_addr[14:5] ? valid_621 : _GEN_644; // @[DCache.scala 78:{33,33}]
  wire  _GEN_646 = 10'h26e == array_addr[14:5] ? valid_622 : _GEN_645; // @[DCache.scala 78:{33,33}]
  wire  _GEN_647 = 10'h26f == array_addr[14:5] ? valid_623 : _GEN_646; // @[DCache.scala 78:{33,33}]
  wire  _GEN_648 = 10'h270 == array_addr[14:5] ? valid_624 : _GEN_647; // @[DCache.scala 78:{33,33}]
  wire  _GEN_649 = 10'h271 == array_addr[14:5] ? valid_625 : _GEN_648; // @[DCache.scala 78:{33,33}]
  wire  _GEN_650 = 10'h272 == array_addr[14:5] ? valid_626 : _GEN_649; // @[DCache.scala 78:{33,33}]
  wire  _GEN_651 = 10'h273 == array_addr[14:5] ? valid_627 : _GEN_650; // @[DCache.scala 78:{33,33}]
  wire  _GEN_652 = 10'h274 == array_addr[14:5] ? valid_628 : _GEN_651; // @[DCache.scala 78:{33,33}]
  wire  _GEN_653 = 10'h275 == array_addr[14:5] ? valid_629 : _GEN_652; // @[DCache.scala 78:{33,33}]
  wire  _GEN_654 = 10'h276 == array_addr[14:5] ? valid_630 : _GEN_653; // @[DCache.scala 78:{33,33}]
  wire  _GEN_655 = 10'h277 == array_addr[14:5] ? valid_631 : _GEN_654; // @[DCache.scala 78:{33,33}]
  wire  _GEN_656 = 10'h278 == array_addr[14:5] ? valid_632 : _GEN_655; // @[DCache.scala 78:{33,33}]
  wire  _GEN_657 = 10'h279 == array_addr[14:5] ? valid_633 : _GEN_656; // @[DCache.scala 78:{33,33}]
  wire  _GEN_658 = 10'h27a == array_addr[14:5] ? valid_634 : _GEN_657; // @[DCache.scala 78:{33,33}]
  wire  _GEN_659 = 10'h27b == array_addr[14:5] ? valid_635 : _GEN_658; // @[DCache.scala 78:{33,33}]
  wire  _GEN_660 = 10'h27c == array_addr[14:5] ? valid_636 : _GEN_659; // @[DCache.scala 78:{33,33}]
  wire  _GEN_661 = 10'h27d == array_addr[14:5] ? valid_637 : _GEN_660; // @[DCache.scala 78:{33,33}]
  wire  _GEN_662 = 10'h27e == array_addr[14:5] ? valid_638 : _GEN_661; // @[DCache.scala 78:{33,33}]
  wire  _GEN_663 = 10'h27f == array_addr[14:5] ? valid_639 : _GEN_662; // @[DCache.scala 78:{33,33}]
  wire  _GEN_664 = 10'h280 == array_addr[14:5] ? valid_640 : _GEN_663; // @[DCache.scala 78:{33,33}]
  wire  _GEN_665 = 10'h281 == array_addr[14:5] ? valid_641 : _GEN_664; // @[DCache.scala 78:{33,33}]
  wire  _GEN_666 = 10'h282 == array_addr[14:5] ? valid_642 : _GEN_665; // @[DCache.scala 78:{33,33}]
  wire  _GEN_667 = 10'h283 == array_addr[14:5] ? valid_643 : _GEN_666; // @[DCache.scala 78:{33,33}]
  wire  _GEN_668 = 10'h284 == array_addr[14:5] ? valid_644 : _GEN_667; // @[DCache.scala 78:{33,33}]
  wire  _GEN_669 = 10'h285 == array_addr[14:5] ? valid_645 : _GEN_668; // @[DCache.scala 78:{33,33}]
  wire  _GEN_670 = 10'h286 == array_addr[14:5] ? valid_646 : _GEN_669; // @[DCache.scala 78:{33,33}]
  wire  _GEN_671 = 10'h287 == array_addr[14:5] ? valid_647 : _GEN_670; // @[DCache.scala 78:{33,33}]
  wire  _GEN_672 = 10'h288 == array_addr[14:5] ? valid_648 : _GEN_671; // @[DCache.scala 78:{33,33}]
  wire  _GEN_673 = 10'h289 == array_addr[14:5] ? valid_649 : _GEN_672; // @[DCache.scala 78:{33,33}]
  wire  _GEN_674 = 10'h28a == array_addr[14:5] ? valid_650 : _GEN_673; // @[DCache.scala 78:{33,33}]
  wire  _GEN_675 = 10'h28b == array_addr[14:5] ? valid_651 : _GEN_674; // @[DCache.scala 78:{33,33}]
  wire  _GEN_676 = 10'h28c == array_addr[14:5] ? valid_652 : _GEN_675; // @[DCache.scala 78:{33,33}]
  wire  _GEN_677 = 10'h28d == array_addr[14:5] ? valid_653 : _GEN_676; // @[DCache.scala 78:{33,33}]
  wire  _GEN_678 = 10'h28e == array_addr[14:5] ? valid_654 : _GEN_677; // @[DCache.scala 78:{33,33}]
  wire  _GEN_679 = 10'h28f == array_addr[14:5] ? valid_655 : _GEN_678; // @[DCache.scala 78:{33,33}]
  wire  _GEN_680 = 10'h290 == array_addr[14:5] ? valid_656 : _GEN_679; // @[DCache.scala 78:{33,33}]
  wire  _GEN_681 = 10'h291 == array_addr[14:5] ? valid_657 : _GEN_680; // @[DCache.scala 78:{33,33}]
  wire  _GEN_682 = 10'h292 == array_addr[14:5] ? valid_658 : _GEN_681; // @[DCache.scala 78:{33,33}]
  wire  _GEN_683 = 10'h293 == array_addr[14:5] ? valid_659 : _GEN_682; // @[DCache.scala 78:{33,33}]
  wire  _GEN_684 = 10'h294 == array_addr[14:5] ? valid_660 : _GEN_683; // @[DCache.scala 78:{33,33}]
  wire  _GEN_685 = 10'h295 == array_addr[14:5] ? valid_661 : _GEN_684; // @[DCache.scala 78:{33,33}]
  wire  _GEN_686 = 10'h296 == array_addr[14:5] ? valid_662 : _GEN_685; // @[DCache.scala 78:{33,33}]
  wire  _GEN_687 = 10'h297 == array_addr[14:5] ? valid_663 : _GEN_686; // @[DCache.scala 78:{33,33}]
  wire  _GEN_688 = 10'h298 == array_addr[14:5] ? valid_664 : _GEN_687; // @[DCache.scala 78:{33,33}]
  wire  _GEN_689 = 10'h299 == array_addr[14:5] ? valid_665 : _GEN_688; // @[DCache.scala 78:{33,33}]
  wire  _GEN_690 = 10'h29a == array_addr[14:5] ? valid_666 : _GEN_689; // @[DCache.scala 78:{33,33}]
  wire  _GEN_691 = 10'h29b == array_addr[14:5] ? valid_667 : _GEN_690; // @[DCache.scala 78:{33,33}]
  wire  _GEN_692 = 10'h29c == array_addr[14:5] ? valid_668 : _GEN_691; // @[DCache.scala 78:{33,33}]
  wire  _GEN_693 = 10'h29d == array_addr[14:5] ? valid_669 : _GEN_692; // @[DCache.scala 78:{33,33}]
  wire  _GEN_694 = 10'h29e == array_addr[14:5] ? valid_670 : _GEN_693; // @[DCache.scala 78:{33,33}]
  wire  _GEN_695 = 10'h29f == array_addr[14:5] ? valid_671 : _GEN_694; // @[DCache.scala 78:{33,33}]
  wire  _GEN_696 = 10'h2a0 == array_addr[14:5] ? valid_672 : _GEN_695; // @[DCache.scala 78:{33,33}]
  wire  _GEN_697 = 10'h2a1 == array_addr[14:5] ? valid_673 : _GEN_696; // @[DCache.scala 78:{33,33}]
  wire  _GEN_698 = 10'h2a2 == array_addr[14:5] ? valid_674 : _GEN_697; // @[DCache.scala 78:{33,33}]
  wire  _GEN_699 = 10'h2a3 == array_addr[14:5] ? valid_675 : _GEN_698; // @[DCache.scala 78:{33,33}]
  wire  _GEN_700 = 10'h2a4 == array_addr[14:5] ? valid_676 : _GEN_699; // @[DCache.scala 78:{33,33}]
  wire  _GEN_701 = 10'h2a5 == array_addr[14:5] ? valid_677 : _GEN_700; // @[DCache.scala 78:{33,33}]
  wire  _GEN_702 = 10'h2a6 == array_addr[14:5] ? valid_678 : _GEN_701; // @[DCache.scala 78:{33,33}]
  wire  _GEN_703 = 10'h2a7 == array_addr[14:5] ? valid_679 : _GEN_702; // @[DCache.scala 78:{33,33}]
  wire  _GEN_704 = 10'h2a8 == array_addr[14:5] ? valid_680 : _GEN_703; // @[DCache.scala 78:{33,33}]
  wire  _GEN_705 = 10'h2a9 == array_addr[14:5] ? valid_681 : _GEN_704; // @[DCache.scala 78:{33,33}]
  wire  _GEN_706 = 10'h2aa == array_addr[14:5] ? valid_682 : _GEN_705; // @[DCache.scala 78:{33,33}]
  wire  _GEN_707 = 10'h2ab == array_addr[14:5] ? valid_683 : _GEN_706; // @[DCache.scala 78:{33,33}]
  wire  _GEN_708 = 10'h2ac == array_addr[14:5] ? valid_684 : _GEN_707; // @[DCache.scala 78:{33,33}]
  wire  _GEN_709 = 10'h2ad == array_addr[14:5] ? valid_685 : _GEN_708; // @[DCache.scala 78:{33,33}]
  wire  _GEN_710 = 10'h2ae == array_addr[14:5] ? valid_686 : _GEN_709; // @[DCache.scala 78:{33,33}]
  wire  _GEN_711 = 10'h2af == array_addr[14:5] ? valid_687 : _GEN_710; // @[DCache.scala 78:{33,33}]
  wire  _GEN_712 = 10'h2b0 == array_addr[14:5] ? valid_688 : _GEN_711; // @[DCache.scala 78:{33,33}]
  wire  _GEN_713 = 10'h2b1 == array_addr[14:5] ? valid_689 : _GEN_712; // @[DCache.scala 78:{33,33}]
  wire  _GEN_714 = 10'h2b2 == array_addr[14:5] ? valid_690 : _GEN_713; // @[DCache.scala 78:{33,33}]
  wire  _GEN_715 = 10'h2b3 == array_addr[14:5] ? valid_691 : _GEN_714; // @[DCache.scala 78:{33,33}]
  wire  _GEN_716 = 10'h2b4 == array_addr[14:5] ? valid_692 : _GEN_715; // @[DCache.scala 78:{33,33}]
  wire  _GEN_717 = 10'h2b5 == array_addr[14:5] ? valid_693 : _GEN_716; // @[DCache.scala 78:{33,33}]
  wire  _GEN_718 = 10'h2b6 == array_addr[14:5] ? valid_694 : _GEN_717; // @[DCache.scala 78:{33,33}]
  wire  _GEN_719 = 10'h2b7 == array_addr[14:5] ? valid_695 : _GEN_718; // @[DCache.scala 78:{33,33}]
  wire  _GEN_720 = 10'h2b8 == array_addr[14:5] ? valid_696 : _GEN_719; // @[DCache.scala 78:{33,33}]
  wire  _GEN_721 = 10'h2b9 == array_addr[14:5] ? valid_697 : _GEN_720; // @[DCache.scala 78:{33,33}]
  wire  _GEN_722 = 10'h2ba == array_addr[14:5] ? valid_698 : _GEN_721; // @[DCache.scala 78:{33,33}]
  wire  _GEN_723 = 10'h2bb == array_addr[14:5] ? valid_699 : _GEN_722; // @[DCache.scala 78:{33,33}]
  wire  _GEN_724 = 10'h2bc == array_addr[14:5] ? valid_700 : _GEN_723; // @[DCache.scala 78:{33,33}]
  wire  _GEN_725 = 10'h2bd == array_addr[14:5] ? valid_701 : _GEN_724; // @[DCache.scala 78:{33,33}]
  wire  _GEN_726 = 10'h2be == array_addr[14:5] ? valid_702 : _GEN_725; // @[DCache.scala 78:{33,33}]
  wire  _GEN_727 = 10'h2bf == array_addr[14:5] ? valid_703 : _GEN_726; // @[DCache.scala 78:{33,33}]
  wire  _GEN_728 = 10'h2c0 == array_addr[14:5] ? valid_704 : _GEN_727; // @[DCache.scala 78:{33,33}]
  wire  _GEN_729 = 10'h2c1 == array_addr[14:5] ? valid_705 : _GEN_728; // @[DCache.scala 78:{33,33}]
  wire  _GEN_730 = 10'h2c2 == array_addr[14:5] ? valid_706 : _GEN_729; // @[DCache.scala 78:{33,33}]
  wire  _GEN_731 = 10'h2c3 == array_addr[14:5] ? valid_707 : _GEN_730; // @[DCache.scala 78:{33,33}]
  wire  _GEN_732 = 10'h2c4 == array_addr[14:5] ? valid_708 : _GEN_731; // @[DCache.scala 78:{33,33}]
  wire  _GEN_733 = 10'h2c5 == array_addr[14:5] ? valid_709 : _GEN_732; // @[DCache.scala 78:{33,33}]
  wire  _GEN_734 = 10'h2c6 == array_addr[14:5] ? valid_710 : _GEN_733; // @[DCache.scala 78:{33,33}]
  wire  _GEN_735 = 10'h2c7 == array_addr[14:5] ? valid_711 : _GEN_734; // @[DCache.scala 78:{33,33}]
  wire  _GEN_736 = 10'h2c8 == array_addr[14:5] ? valid_712 : _GEN_735; // @[DCache.scala 78:{33,33}]
  wire  _GEN_737 = 10'h2c9 == array_addr[14:5] ? valid_713 : _GEN_736; // @[DCache.scala 78:{33,33}]
  wire  _GEN_738 = 10'h2ca == array_addr[14:5] ? valid_714 : _GEN_737; // @[DCache.scala 78:{33,33}]
  wire  _GEN_739 = 10'h2cb == array_addr[14:5] ? valid_715 : _GEN_738; // @[DCache.scala 78:{33,33}]
  wire  _GEN_740 = 10'h2cc == array_addr[14:5] ? valid_716 : _GEN_739; // @[DCache.scala 78:{33,33}]
  wire  _GEN_741 = 10'h2cd == array_addr[14:5] ? valid_717 : _GEN_740; // @[DCache.scala 78:{33,33}]
  wire  _GEN_742 = 10'h2ce == array_addr[14:5] ? valid_718 : _GEN_741; // @[DCache.scala 78:{33,33}]
  wire  _GEN_743 = 10'h2cf == array_addr[14:5] ? valid_719 : _GEN_742; // @[DCache.scala 78:{33,33}]
  wire  _GEN_744 = 10'h2d0 == array_addr[14:5] ? valid_720 : _GEN_743; // @[DCache.scala 78:{33,33}]
  wire  _GEN_745 = 10'h2d1 == array_addr[14:5] ? valid_721 : _GEN_744; // @[DCache.scala 78:{33,33}]
  wire  _GEN_746 = 10'h2d2 == array_addr[14:5] ? valid_722 : _GEN_745; // @[DCache.scala 78:{33,33}]
  wire  _GEN_747 = 10'h2d3 == array_addr[14:5] ? valid_723 : _GEN_746; // @[DCache.scala 78:{33,33}]
  wire  _GEN_748 = 10'h2d4 == array_addr[14:5] ? valid_724 : _GEN_747; // @[DCache.scala 78:{33,33}]
  wire  _GEN_749 = 10'h2d5 == array_addr[14:5] ? valid_725 : _GEN_748; // @[DCache.scala 78:{33,33}]
  wire  _GEN_750 = 10'h2d6 == array_addr[14:5] ? valid_726 : _GEN_749; // @[DCache.scala 78:{33,33}]
  wire  _GEN_751 = 10'h2d7 == array_addr[14:5] ? valid_727 : _GEN_750; // @[DCache.scala 78:{33,33}]
  wire  _GEN_752 = 10'h2d8 == array_addr[14:5] ? valid_728 : _GEN_751; // @[DCache.scala 78:{33,33}]
  wire  _GEN_753 = 10'h2d9 == array_addr[14:5] ? valid_729 : _GEN_752; // @[DCache.scala 78:{33,33}]
  wire  _GEN_754 = 10'h2da == array_addr[14:5] ? valid_730 : _GEN_753; // @[DCache.scala 78:{33,33}]
  wire  _GEN_755 = 10'h2db == array_addr[14:5] ? valid_731 : _GEN_754; // @[DCache.scala 78:{33,33}]
  wire  _GEN_756 = 10'h2dc == array_addr[14:5] ? valid_732 : _GEN_755; // @[DCache.scala 78:{33,33}]
  wire  _GEN_757 = 10'h2dd == array_addr[14:5] ? valid_733 : _GEN_756; // @[DCache.scala 78:{33,33}]
  wire  _GEN_758 = 10'h2de == array_addr[14:5] ? valid_734 : _GEN_757; // @[DCache.scala 78:{33,33}]
  wire  _GEN_759 = 10'h2df == array_addr[14:5] ? valid_735 : _GEN_758; // @[DCache.scala 78:{33,33}]
  wire  _GEN_760 = 10'h2e0 == array_addr[14:5] ? valid_736 : _GEN_759; // @[DCache.scala 78:{33,33}]
  wire  _GEN_761 = 10'h2e1 == array_addr[14:5] ? valid_737 : _GEN_760; // @[DCache.scala 78:{33,33}]
  wire  _GEN_762 = 10'h2e2 == array_addr[14:5] ? valid_738 : _GEN_761; // @[DCache.scala 78:{33,33}]
  wire  _GEN_763 = 10'h2e3 == array_addr[14:5] ? valid_739 : _GEN_762; // @[DCache.scala 78:{33,33}]
  wire  _GEN_764 = 10'h2e4 == array_addr[14:5] ? valid_740 : _GEN_763; // @[DCache.scala 78:{33,33}]
  wire  _GEN_765 = 10'h2e5 == array_addr[14:5] ? valid_741 : _GEN_764; // @[DCache.scala 78:{33,33}]
  wire  _GEN_766 = 10'h2e6 == array_addr[14:5] ? valid_742 : _GEN_765; // @[DCache.scala 78:{33,33}]
  wire  _GEN_767 = 10'h2e7 == array_addr[14:5] ? valid_743 : _GEN_766; // @[DCache.scala 78:{33,33}]
  wire  _GEN_768 = 10'h2e8 == array_addr[14:5] ? valid_744 : _GEN_767; // @[DCache.scala 78:{33,33}]
  wire  _GEN_769 = 10'h2e9 == array_addr[14:5] ? valid_745 : _GEN_768; // @[DCache.scala 78:{33,33}]
  wire  _GEN_770 = 10'h2ea == array_addr[14:5] ? valid_746 : _GEN_769; // @[DCache.scala 78:{33,33}]
  wire  _GEN_771 = 10'h2eb == array_addr[14:5] ? valid_747 : _GEN_770; // @[DCache.scala 78:{33,33}]
  wire  _GEN_772 = 10'h2ec == array_addr[14:5] ? valid_748 : _GEN_771; // @[DCache.scala 78:{33,33}]
  wire  _GEN_773 = 10'h2ed == array_addr[14:5] ? valid_749 : _GEN_772; // @[DCache.scala 78:{33,33}]
  wire  _GEN_774 = 10'h2ee == array_addr[14:5] ? valid_750 : _GEN_773; // @[DCache.scala 78:{33,33}]
  wire  _GEN_775 = 10'h2ef == array_addr[14:5] ? valid_751 : _GEN_774; // @[DCache.scala 78:{33,33}]
  wire  _GEN_776 = 10'h2f0 == array_addr[14:5] ? valid_752 : _GEN_775; // @[DCache.scala 78:{33,33}]
  wire  _GEN_777 = 10'h2f1 == array_addr[14:5] ? valid_753 : _GEN_776; // @[DCache.scala 78:{33,33}]
  wire  _GEN_778 = 10'h2f2 == array_addr[14:5] ? valid_754 : _GEN_777; // @[DCache.scala 78:{33,33}]
  wire  _GEN_779 = 10'h2f3 == array_addr[14:5] ? valid_755 : _GEN_778; // @[DCache.scala 78:{33,33}]
  wire  _GEN_780 = 10'h2f4 == array_addr[14:5] ? valid_756 : _GEN_779; // @[DCache.scala 78:{33,33}]
  wire  _GEN_781 = 10'h2f5 == array_addr[14:5] ? valid_757 : _GEN_780; // @[DCache.scala 78:{33,33}]
  wire  _GEN_782 = 10'h2f6 == array_addr[14:5] ? valid_758 : _GEN_781; // @[DCache.scala 78:{33,33}]
  wire  _GEN_783 = 10'h2f7 == array_addr[14:5] ? valid_759 : _GEN_782; // @[DCache.scala 78:{33,33}]
  wire  _GEN_784 = 10'h2f8 == array_addr[14:5] ? valid_760 : _GEN_783; // @[DCache.scala 78:{33,33}]
  wire  _GEN_785 = 10'h2f9 == array_addr[14:5] ? valid_761 : _GEN_784; // @[DCache.scala 78:{33,33}]
  wire  _GEN_786 = 10'h2fa == array_addr[14:5] ? valid_762 : _GEN_785; // @[DCache.scala 78:{33,33}]
  wire  _GEN_787 = 10'h2fb == array_addr[14:5] ? valid_763 : _GEN_786; // @[DCache.scala 78:{33,33}]
  wire  _GEN_788 = 10'h2fc == array_addr[14:5] ? valid_764 : _GEN_787; // @[DCache.scala 78:{33,33}]
  wire  _GEN_789 = 10'h2fd == array_addr[14:5] ? valid_765 : _GEN_788; // @[DCache.scala 78:{33,33}]
  wire  _GEN_790 = 10'h2fe == array_addr[14:5] ? valid_766 : _GEN_789; // @[DCache.scala 78:{33,33}]
  wire  _GEN_791 = 10'h2ff == array_addr[14:5] ? valid_767 : _GEN_790; // @[DCache.scala 78:{33,33}]
  wire  _GEN_792 = 10'h300 == array_addr[14:5] ? valid_768 : _GEN_791; // @[DCache.scala 78:{33,33}]
  wire  _GEN_793 = 10'h301 == array_addr[14:5] ? valid_769 : _GEN_792; // @[DCache.scala 78:{33,33}]
  wire  _GEN_794 = 10'h302 == array_addr[14:5] ? valid_770 : _GEN_793; // @[DCache.scala 78:{33,33}]
  wire  _GEN_795 = 10'h303 == array_addr[14:5] ? valid_771 : _GEN_794; // @[DCache.scala 78:{33,33}]
  wire  _GEN_796 = 10'h304 == array_addr[14:5] ? valid_772 : _GEN_795; // @[DCache.scala 78:{33,33}]
  wire  _GEN_797 = 10'h305 == array_addr[14:5] ? valid_773 : _GEN_796; // @[DCache.scala 78:{33,33}]
  wire  _GEN_798 = 10'h306 == array_addr[14:5] ? valid_774 : _GEN_797; // @[DCache.scala 78:{33,33}]
  wire  _GEN_799 = 10'h307 == array_addr[14:5] ? valid_775 : _GEN_798; // @[DCache.scala 78:{33,33}]
  wire  _GEN_800 = 10'h308 == array_addr[14:5] ? valid_776 : _GEN_799; // @[DCache.scala 78:{33,33}]
  wire  _GEN_801 = 10'h309 == array_addr[14:5] ? valid_777 : _GEN_800; // @[DCache.scala 78:{33,33}]
  wire  _GEN_802 = 10'h30a == array_addr[14:5] ? valid_778 : _GEN_801; // @[DCache.scala 78:{33,33}]
  wire  _GEN_803 = 10'h30b == array_addr[14:5] ? valid_779 : _GEN_802; // @[DCache.scala 78:{33,33}]
  wire  _GEN_804 = 10'h30c == array_addr[14:5] ? valid_780 : _GEN_803; // @[DCache.scala 78:{33,33}]
  wire  _GEN_805 = 10'h30d == array_addr[14:5] ? valid_781 : _GEN_804; // @[DCache.scala 78:{33,33}]
  wire  _GEN_806 = 10'h30e == array_addr[14:5] ? valid_782 : _GEN_805; // @[DCache.scala 78:{33,33}]
  wire  _GEN_807 = 10'h30f == array_addr[14:5] ? valid_783 : _GEN_806; // @[DCache.scala 78:{33,33}]
  wire  _GEN_808 = 10'h310 == array_addr[14:5] ? valid_784 : _GEN_807; // @[DCache.scala 78:{33,33}]
  wire  _GEN_809 = 10'h311 == array_addr[14:5] ? valid_785 : _GEN_808; // @[DCache.scala 78:{33,33}]
  wire  _GEN_810 = 10'h312 == array_addr[14:5] ? valid_786 : _GEN_809; // @[DCache.scala 78:{33,33}]
  wire  _GEN_811 = 10'h313 == array_addr[14:5] ? valid_787 : _GEN_810; // @[DCache.scala 78:{33,33}]
  wire  _GEN_812 = 10'h314 == array_addr[14:5] ? valid_788 : _GEN_811; // @[DCache.scala 78:{33,33}]
  wire  _GEN_813 = 10'h315 == array_addr[14:5] ? valid_789 : _GEN_812; // @[DCache.scala 78:{33,33}]
  wire  _GEN_814 = 10'h316 == array_addr[14:5] ? valid_790 : _GEN_813; // @[DCache.scala 78:{33,33}]
  wire  _GEN_815 = 10'h317 == array_addr[14:5] ? valid_791 : _GEN_814; // @[DCache.scala 78:{33,33}]
  wire  _GEN_816 = 10'h318 == array_addr[14:5] ? valid_792 : _GEN_815; // @[DCache.scala 78:{33,33}]
  wire  _GEN_817 = 10'h319 == array_addr[14:5] ? valid_793 : _GEN_816; // @[DCache.scala 78:{33,33}]
  wire  _GEN_818 = 10'h31a == array_addr[14:5] ? valid_794 : _GEN_817; // @[DCache.scala 78:{33,33}]
  wire  _GEN_819 = 10'h31b == array_addr[14:5] ? valid_795 : _GEN_818; // @[DCache.scala 78:{33,33}]
  wire  _GEN_820 = 10'h31c == array_addr[14:5] ? valid_796 : _GEN_819; // @[DCache.scala 78:{33,33}]
  wire  _GEN_821 = 10'h31d == array_addr[14:5] ? valid_797 : _GEN_820; // @[DCache.scala 78:{33,33}]
  wire  _GEN_822 = 10'h31e == array_addr[14:5] ? valid_798 : _GEN_821; // @[DCache.scala 78:{33,33}]
  wire  _GEN_823 = 10'h31f == array_addr[14:5] ? valid_799 : _GEN_822; // @[DCache.scala 78:{33,33}]
  wire  _GEN_824 = 10'h320 == array_addr[14:5] ? valid_800 : _GEN_823; // @[DCache.scala 78:{33,33}]
  wire  _GEN_825 = 10'h321 == array_addr[14:5] ? valid_801 : _GEN_824; // @[DCache.scala 78:{33,33}]
  wire  _GEN_826 = 10'h322 == array_addr[14:5] ? valid_802 : _GEN_825; // @[DCache.scala 78:{33,33}]
  wire  _GEN_827 = 10'h323 == array_addr[14:5] ? valid_803 : _GEN_826; // @[DCache.scala 78:{33,33}]
  wire  _GEN_828 = 10'h324 == array_addr[14:5] ? valid_804 : _GEN_827; // @[DCache.scala 78:{33,33}]
  wire  _GEN_829 = 10'h325 == array_addr[14:5] ? valid_805 : _GEN_828; // @[DCache.scala 78:{33,33}]
  wire  _GEN_830 = 10'h326 == array_addr[14:5] ? valid_806 : _GEN_829; // @[DCache.scala 78:{33,33}]
  wire  _GEN_831 = 10'h327 == array_addr[14:5] ? valid_807 : _GEN_830; // @[DCache.scala 78:{33,33}]
  wire  _GEN_832 = 10'h328 == array_addr[14:5] ? valid_808 : _GEN_831; // @[DCache.scala 78:{33,33}]
  wire  _GEN_833 = 10'h329 == array_addr[14:5] ? valid_809 : _GEN_832; // @[DCache.scala 78:{33,33}]
  wire  _GEN_834 = 10'h32a == array_addr[14:5] ? valid_810 : _GEN_833; // @[DCache.scala 78:{33,33}]
  wire  _GEN_835 = 10'h32b == array_addr[14:5] ? valid_811 : _GEN_834; // @[DCache.scala 78:{33,33}]
  wire  _GEN_836 = 10'h32c == array_addr[14:5] ? valid_812 : _GEN_835; // @[DCache.scala 78:{33,33}]
  wire  _GEN_837 = 10'h32d == array_addr[14:5] ? valid_813 : _GEN_836; // @[DCache.scala 78:{33,33}]
  wire  _GEN_838 = 10'h32e == array_addr[14:5] ? valid_814 : _GEN_837; // @[DCache.scala 78:{33,33}]
  wire  _GEN_839 = 10'h32f == array_addr[14:5] ? valid_815 : _GEN_838; // @[DCache.scala 78:{33,33}]
  wire  _GEN_840 = 10'h330 == array_addr[14:5] ? valid_816 : _GEN_839; // @[DCache.scala 78:{33,33}]
  wire  _GEN_841 = 10'h331 == array_addr[14:5] ? valid_817 : _GEN_840; // @[DCache.scala 78:{33,33}]
  wire  _GEN_842 = 10'h332 == array_addr[14:5] ? valid_818 : _GEN_841; // @[DCache.scala 78:{33,33}]
  wire  _GEN_843 = 10'h333 == array_addr[14:5] ? valid_819 : _GEN_842; // @[DCache.scala 78:{33,33}]
  wire  _GEN_844 = 10'h334 == array_addr[14:5] ? valid_820 : _GEN_843; // @[DCache.scala 78:{33,33}]
  wire  _GEN_845 = 10'h335 == array_addr[14:5] ? valid_821 : _GEN_844; // @[DCache.scala 78:{33,33}]
  wire  _GEN_846 = 10'h336 == array_addr[14:5] ? valid_822 : _GEN_845; // @[DCache.scala 78:{33,33}]
  wire  _GEN_847 = 10'h337 == array_addr[14:5] ? valid_823 : _GEN_846; // @[DCache.scala 78:{33,33}]
  wire  _GEN_848 = 10'h338 == array_addr[14:5] ? valid_824 : _GEN_847; // @[DCache.scala 78:{33,33}]
  wire  _GEN_849 = 10'h339 == array_addr[14:5] ? valid_825 : _GEN_848; // @[DCache.scala 78:{33,33}]
  wire  _GEN_850 = 10'h33a == array_addr[14:5] ? valid_826 : _GEN_849; // @[DCache.scala 78:{33,33}]
  wire  _GEN_851 = 10'h33b == array_addr[14:5] ? valid_827 : _GEN_850; // @[DCache.scala 78:{33,33}]
  wire  _GEN_852 = 10'h33c == array_addr[14:5] ? valid_828 : _GEN_851; // @[DCache.scala 78:{33,33}]
  wire  _GEN_853 = 10'h33d == array_addr[14:5] ? valid_829 : _GEN_852; // @[DCache.scala 78:{33,33}]
  wire  _GEN_854 = 10'h33e == array_addr[14:5] ? valid_830 : _GEN_853; // @[DCache.scala 78:{33,33}]
  wire  _GEN_855 = 10'h33f == array_addr[14:5] ? valid_831 : _GEN_854; // @[DCache.scala 78:{33,33}]
  wire  _GEN_856 = 10'h340 == array_addr[14:5] ? valid_832 : _GEN_855; // @[DCache.scala 78:{33,33}]
  wire  _GEN_857 = 10'h341 == array_addr[14:5] ? valid_833 : _GEN_856; // @[DCache.scala 78:{33,33}]
  wire  _GEN_858 = 10'h342 == array_addr[14:5] ? valid_834 : _GEN_857; // @[DCache.scala 78:{33,33}]
  wire  _GEN_859 = 10'h343 == array_addr[14:5] ? valid_835 : _GEN_858; // @[DCache.scala 78:{33,33}]
  wire  _GEN_860 = 10'h344 == array_addr[14:5] ? valid_836 : _GEN_859; // @[DCache.scala 78:{33,33}]
  wire  _GEN_861 = 10'h345 == array_addr[14:5] ? valid_837 : _GEN_860; // @[DCache.scala 78:{33,33}]
  wire  _GEN_862 = 10'h346 == array_addr[14:5] ? valid_838 : _GEN_861; // @[DCache.scala 78:{33,33}]
  wire  _GEN_863 = 10'h347 == array_addr[14:5] ? valid_839 : _GEN_862; // @[DCache.scala 78:{33,33}]
  wire  _GEN_864 = 10'h348 == array_addr[14:5] ? valid_840 : _GEN_863; // @[DCache.scala 78:{33,33}]
  wire  _GEN_865 = 10'h349 == array_addr[14:5] ? valid_841 : _GEN_864; // @[DCache.scala 78:{33,33}]
  wire  _GEN_866 = 10'h34a == array_addr[14:5] ? valid_842 : _GEN_865; // @[DCache.scala 78:{33,33}]
  wire  _GEN_867 = 10'h34b == array_addr[14:5] ? valid_843 : _GEN_866; // @[DCache.scala 78:{33,33}]
  wire  _GEN_868 = 10'h34c == array_addr[14:5] ? valid_844 : _GEN_867; // @[DCache.scala 78:{33,33}]
  wire  _GEN_869 = 10'h34d == array_addr[14:5] ? valid_845 : _GEN_868; // @[DCache.scala 78:{33,33}]
  wire  _GEN_870 = 10'h34e == array_addr[14:5] ? valid_846 : _GEN_869; // @[DCache.scala 78:{33,33}]
  wire  _GEN_871 = 10'h34f == array_addr[14:5] ? valid_847 : _GEN_870; // @[DCache.scala 78:{33,33}]
  wire  _GEN_872 = 10'h350 == array_addr[14:5] ? valid_848 : _GEN_871; // @[DCache.scala 78:{33,33}]
  wire  _GEN_873 = 10'h351 == array_addr[14:5] ? valid_849 : _GEN_872; // @[DCache.scala 78:{33,33}]
  wire  _GEN_874 = 10'h352 == array_addr[14:5] ? valid_850 : _GEN_873; // @[DCache.scala 78:{33,33}]
  wire  _GEN_875 = 10'h353 == array_addr[14:5] ? valid_851 : _GEN_874; // @[DCache.scala 78:{33,33}]
  wire  _GEN_876 = 10'h354 == array_addr[14:5] ? valid_852 : _GEN_875; // @[DCache.scala 78:{33,33}]
  wire  _GEN_877 = 10'h355 == array_addr[14:5] ? valid_853 : _GEN_876; // @[DCache.scala 78:{33,33}]
  wire  _GEN_878 = 10'h356 == array_addr[14:5] ? valid_854 : _GEN_877; // @[DCache.scala 78:{33,33}]
  wire  _GEN_879 = 10'h357 == array_addr[14:5] ? valid_855 : _GEN_878; // @[DCache.scala 78:{33,33}]
  wire  _GEN_880 = 10'h358 == array_addr[14:5] ? valid_856 : _GEN_879; // @[DCache.scala 78:{33,33}]
  wire  _GEN_881 = 10'h359 == array_addr[14:5] ? valid_857 : _GEN_880; // @[DCache.scala 78:{33,33}]
  wire  _GEN_882 = 10'h35a == array_addr[14:5] ? valid_858 : _GEN_881; // @[DCache.scala 78:{33,33}]
  wire  _GEN_883 = 10'h35b == array_addr[14:5] ? valid_859 : _GEN_882; // @[DCache.scala 78:{33,33}]
  wire  _GEN_884 = 10'h35c == array_addr[14:5] ? valid_860 : _GEN_883; // @[DCache.scala 78:{33,33}]
  wire  _GEN_885 = 10'h35d == array_addr[14:5] ? valid_861 : _GEN_884; // @[DCache.scala 78:{33,33}]
  wire  _GEN_886 = 10'h35e == array_addr[14:5] ? valid_862 : _GEN_885; // @[DCache.scala 78:{33,33}]
  wire  _GEN_887 = 10'h35f == array_addr[14:5] ? valid_863 : _GEN_886; // @[DCache.scala 78:{33,33}]
  wire  _GEN_888 = 10'h360 == array_addr[14:5] ? valid_864 : _GEN_887; // @[DCache.scala 78:{33,33}]
  wire  _GEN_889 = 10'h361 == array_addr[14:5] ? valid_865 : _GEN_888; // @[DCache.scala 78:{33,33}]
  wire  _GEN_890 = 10'h362 == array_addr[14:5] ? valid_866 : _GEN_889; // @[DCache.scala 78:{33,33}]
  wire  _GEN_891 = 10'h363 == array_addr[14:5] ? valid_867 : _GEN_890; // @[DCache.scala 78:{33,33}]
  wire  _GEN_892 = 10'h364 == array_addr[14:5] ? valid_868 : _GEN_891; // @[DCache.scala 78:{33,33}]
  wire  _GEN_893 = 10'h365 == array_addr[14:5] ? valid_869 : _GEN_892; // @[DCache.scala 78:{33,33}]
  wire  _GEN_894 = 10'h366 == array_addr[14:5] ? valid_870 : _GEN_893; // @[DCache.scala 78:{33,33}]
  wire  _GEN_895 = 10'h367 == array_addr[14:5] ? valid_871 : _GEN_894; // @[DCache.scala 78:{33,33}]
  wire  _GEN_896 = 10'h368 == array_addr[14:5] ? valid_872 : _GEN_895; // @[DCache.scala 78:{33,33}]
  wire  _GEN_897 = 10'h369 == array_addr[14:5] ? valid_873 : _GEN_896; // @[DCache.scala 78:{33,33}]
  wire  _GEN_898 = 10'h36a == array_addr[14:5] ? valid_874 : _GEN_897; // @[DCache.scala 78:{33,33}]
  wire  _GEN_899 = 10'h36b == array_addr[14:5] ? valid_875 : _GEN_898; // @[DCache.scala 78:{33,33}]
  wire  _GEN_900 = 10'h36c == array_addr[14:5] ? valid_876 : _GEN_899; // @[DCache.scala 78:{33,33}]
  wire  _GEN_901 = 10'h36d == array_addr[14:5] ? valid_877 : _GEN_900; // @[DCache.scala 78:{33,33}]
  wire  _GEN_902 = 10'h36e == array_addr[14:5] ? valid_878 : _GEN_901; // @[DCache.scala 78:{33,33}]
  wire  _GEN_903 = 10'h36f == array_addr[14:5] ? valid_879 : _GEN_902; // @[DCache.scala 78:{33,33}]
  wire  _GEN_904 = 10'h370 == array_addr[14:5] ? valid_880 : _GEN_903; // @[DCache.scala 78:{33,33}]
  wire  _GEN_905 = 10'h371 == array_addr[14:5] ? valid_881 : _GEN_904; // @[DCache.scala 78:{33,33}]
  wire  _GEN_906 = 10'h372 == array_addr[14:5] ? valid_882 : _GEN_905; // @[DCache.scala 78:{33,33}]
  wire  _GEN_907 = 10'h373 == array_addr[14:5] ? valid_883 : _GEN_906; // @[DCache.scala 78:{33,33}]
  wire  _GEN_908 = 10'h374 == array_addr[14:5] ? valid_884 : _GEN_907; // @[DCache.scala 78:{33,33}]
  wire  _GEN_909 = 10'h375 == array_addr[14:5] ? valid_885 : _GEN_908; // @[DCache.scala 78:{33,33}]
  wire  _GEN_910 = 10'h376 == array_addr[14:5] ? valid_886 : _GEN_909; // @[DCache.scala 78:{33,33}]
  wire  _GEN_911 = 10'h377 == array_addr[14:5] ? valid_887 : _GEN_910; // @[DCache.scala 78:{33,33}]
  wire  _GEN_912 = 10'h378 == array_addr[14:5] ? valid_888 : _GEN_911; // @[DCache.scala 78:{33,33}]
  wire  _GEN_913 = 10'h379 == array_addr[14:5] ? valid_889 : _GEN_912; // @[DCache.scala 78:{33,33}]
  wire  _GEN_914 = 10'h37a == array_addr[14:5] ? valid_890 : _GEN_913; // @[DCache.scala 78:{33,33}]
  wire  _GEN_915 = 10'h37b == array_addr[14:5] ? valid_891 : _GEN_914; // @[DCache.scala 78:{33,33}]
  wire  _GEN_916 = 10'h37c == array_addr[14:5] ? valid_892 : _GEN_915; // @[DCache.scala 78:{33,33}]
  wire  _GEN_917 = 10'h37d == array_addr[14:5] ? valid_893 : _GEN_916; // @[DCache.scala 78:{33,33}]
  wire  _GEN_918 = 10'h37e == array_addr[14:5] ? valid_894 : _GEN_917; // @[DCache.scala 78:{33,33}]
  wire  _GEN_919 = 10'h37f == array_addr[14:5] ? valid_895 : _GEN_918; // @[DCache.scala 78:{33,33}]
  wire  _GEN_920 = 10'h380 == array_addr[14:5] ? valid_896 : _GEN_919; // @[DCache.scala 78:{33,33}]
  wire  _GEN_921 = 10'h381 == array_addr[14:5] ? valid_897 : _GEN_920; // @[DCache.scala 78:{33,33}]
  wire  _GEN_922 = 10'h382 == array_addr[14:5] ? valid_898 : _GEN_921; // @[DCache.scala 78:{33,33}]
  wire  _GEN_923 = 10'h383 == array_addr[14:5] ? valid_899 : _GEN_922; // @[DCache.scala 78:{33,33}]
  wire  _GEN_924 = 10'h384 == array_addr[14:5] ? valid_900 : _GEN_923; // @[DCache.scala 78:{33,33}]
  wire  _GEN_925 = 10'h385 == array_addr[14:5] ? valid_901 : _GEN_924; // @[DCache.scala 78:{33,33}]
  wire  _GEN_926 = 10'h386 == array_addr[14:5] ? valid_902 : _GEN_925; // @[DCache.scala 78:{33,33}]
  wire  _GEN_927 = 10'h387 == array_addr[14:5] ? valid_903 : _GEN_926; // @[DCache.scala 78:{33,33}]
  wire  _GEN_928 = 10'h388 == array_addr[14:5] ? valid_904 : _GEN_927; // @[DCache.scala 78:{33,33}]
  wire  _GEN_929 = 10'h389 == array_addr[14:5] ? valid_905 : _GEN_928; // @[DCache.scala 78:{33,33}]
  wire  _GEN_930 = 10'h38a == array_addr[14:5] ? valid_906 : _GEN_929; // @[DCache.scala 78:{33,33}]
  wire  _GEN_931 = 10'h38b == array_addr[14:5] ? valid_907 : _GEN_930; // @[DCache.scala 78:{33,33}]
  wire  _GEN_932 = 10'h38c == array_addr[14:5] ? valid_908 : _GEN_931; // @[DCache.scala 78:{33,33}]
  wire  _GEN_933 = 10'h38d == array_addr[14:5] ? valid_909 : _GEN_932; // @[DCache.scala 78:{33,33}]
  wire  _GEN_934 = 10'h38e == array_addr[14:5] ? valid_910 : _GEN_933; // @[DCache.scala 78:{33,33}]
  wire  _GEN_935 = 10'h38f == array_addr[14:5] ? valid_911 : _GEN_934; // @[DCache.scala 78:{33,33}]
  wire  _GEN_936 = 10'h390 == array_addr[14:5] ? valid_912 : _GEN_935; // @[DCache.scala 78:{33,33}]
  wire  _GEN_937 = 10'h391 == array_addr[14:5] ? valid_913 : _GEN_936; // @[DCache.scala 78:{33,33}]
  wire  _GEN_938 = 10'h392 == array_addr[14:5] ? valid_914 : _GEN_937; // @[DCache.scala 78:{33,33}]
  wire  _GEN_939 = 10'h393 == array_addr[14:5] ? valid_915 : _GEN_938; // @[DCache.scala 78:{33,33}]
  wire  _GEN_940 = 10'h394 == array_addr[14:5] ? valid_916 : _GEN_939; // @[DCache.scala 78:{33,33}]
  wire  _GEN_941 = 10'h395 == array_addr[14:5] ? valid_917 : _GEN_940; // @[DCache.scala 78:{33,33}]
  wire  _GEN_942 = 10'h396 == array_addr[14:5] ? valid_918 : _GEN_941; // @[DCache.scala 78:{33,33}]
  wire  _GEN_943 = 10'h397 == array_addr[14:5] ? valid_919 : _GEN_942; // @[DCache.scala 78:{33,33}]
  wire  _GEN_944 = 10'h398 == array_addr[14:5] ? valid_920 : _GEN_943; // @[DCache.scala 78:{33,33}]
  wire  _GEN_945 = 10'h399 == array_addr[14:5] ? valid_921 : _GEN_944; // @[DCache.scala 78:{33,33}]
  wire  _GEN_946 = 10'h39a == array_addr[14:5] ? valid_922 : _GEN_945; // @[DCache.scala 78:{33,33}]
  wire  _GEN_947 = 10'h39b == array_addr[14:5] ? valid_923 : _GEN_946; // @[DCache.scala 78:{33,33}]
  wire  _GEN_948 = 10'h39c == array_addr[14:5] ? valid_924 : _GEN_947; // @[DCache.scala 78:{33,33}]
  wire  _GEN_949 = 10'h39d == array_addr[14:5] ? valid_925 : _GEN_948; // @[DCache.scala 78:{33,33}]
  wire  _GEN_950 = 10'h39e == array_addr[14:5] ? valid_926 : _GEN_949; // @[DCache.scala 78:{33,33}]
  wire  _GEN_951 = 10'h39f == array_addr[14:5] ? valid_927 : _GEN_950; // @[DCache.scala 78:{33,33}]
  wire  _GEN_952 = 10'h3a0 == array_addr[14:5] ? valid_928 : _GEN_951; // @[DCache.scala 78:{33,33}]
  wire  _GEN_953 = 10'h3a1 == array_addr[14:5] ? valid_929 : _GEN_952; // @[DCache.scala 78:{33,33}]
  wire  _GEN_954 = 10'h3a2 == array_addr[14:5] ? valid_930 : _GEN_953; // @[DCache.scala 78:{33,33}]
  wire  _GEN_955 = 10'h3a3 == array_addr[14:5] ? valid_931 : _GEN_954; // @[DCache.scala 78:{33,33}]
  wire  _GEN_956 = 10'h3a4 == array_addr[14:5] ? valid_932 : _GEN_955; // @[DCache.scala 78:{33,33}]
  wire  _GEN_957 = 10'h3a5 == array_addr[14:5] ? valid_933 : _GEN_956; // @[DCache.scala 78:{33,33}]
  wire  _GEN_958 = 10'h3a6 == array_addr[14:5] ? valid_934 : _GEN_957; // @[DCache.scala 78:{33,33}]
  wire  _GEN_959 = 10'h3a7 == array_addr[14:5] ? valid_935 : _GEN_958; // @[DCache.scala 78:{33,33}]
  wire  _GEN_960 = 10'h3a8 == array_addr[14:5] ? valid_936 : _GEN_959; // @[DCache.scala 78:{33,33}]
  wire  _GEN_961 = 10'h3a9 == array_addr[14:5] ? valid_937 : _GEN_960; // @[DCache.scala 78:{33,33}]
  wire  _GEN_962 = 10'h3aa == array_addr[14:5] ? valid_938 : _GEN_961; // @[DCache.scala 78:{33,33}]
  wire  _GEN_963 = 10'h3ab == array_addr[14:5] ? valid_939 : _GEN_962; // @[DCache.scala 78:{33,33}]
  wire  _GEN_964 = 10'h3ac == array_addr[14:5] ? valid_940 : _GEN_963; // @[DCache.scala 78:{33,33}]
  wire  _GEN_965 = 10'h3ad == array_addr[14:5] ? valid_941 : _GEN_964; // @[DCache.scala 78:{33,33}]
  wire  _GEN_966 = 10'h3ae == array_addr[14:5] ? valid_942 : _GEN_965; // @[DCache.scala 78:{33,33}]
  wire  _GEN_967 = 10'h3af == array_addr[14:5] ? valid_943 : _GEN_966; // @[DCache.scala 78:{33,33}]
  wire  _GEN_968 = 10'h3b0 == array_addr[14:5] ? valid_944 : _GEN_967; // @[DCache.scala 78:{33,33}]
  wire  _GEN_969 = 10'h3b1 == array_addr[14:5] ? valid_945 : _GEN_968; // @[DCache.scala 78:{33,33}]
  wire  _GEN_970 = 10'h3b2 == array_addr[14:5] ? valid_946 : _GEN_969; // @[DCache.scala 78:{33,33}]
  wire  _GEN_971 = 10'h3b3 == array_addr[14:5] ? valid_947 : _GEN_970; // @[DCache.scala 78:{33,33}]
  wire  _GEN_972 = 10'h3b4 == array_addr[14:5] ? valid_948 : _GEN_971; // @[DCache.scala 78:{33,33}]
  wire  _GEN_973 = 10'h3b5 == array_addr[14:5] ? valid_949 : _GEN_972; // @[DCache.scala 78:{33,33}]
  wire  _GEN_974 = 10'h3b6 == array_addr[14:5] ? valid_950 : _GEN_973; // @[DCache.scala 78:{33,33}]
  wire  _GEN_975 = 10'h3b7 == array_addr[14:5] ? valid_951 : _GEN_974; // @[DCache.scala 78:{33,33}]
  wire  _GEN_976 = 10'h3b8 == array_addr[14:5] ? valid_952 : _GEN_975; // @[DCache.scala 78:{33,33}]
  wire  _GEN_977 = 10'h3b9 == array_addr[14:5] ? valid_953 : _GEN_976; // @[DCache.scala 78:{33,33}]
  wire  _GEN_978 = 10'h3ba == array_addr[14:5] ? valid_954 : _GEN_977; // @[DCache.scala 78:{33,33}]
  wire  _GEN_979 = 10'h3bb == array_addr[14:5] ? valid_955 : _GEN_978; // @[DCache.scala 78:{33,33}]
  wire  _GEN_980 = 10'h3bc == array_addr[14:5] ? valid_956 : _GEN_979; // @[DCache.scala 78:{33,33}]
  wire  _GEN_981 = 10'h3bd == array_addr[14:5] ? valid_957 : _GEN_980; // @[DCache.scala 78:{33,33}]
  wire  _GEN_982 = 10'h3be == array_addr[14:5] ? valid_958 : _GEN_981; // @[DCache.scala 78:{33,33}]
  wire  _GEN_983 = 10'h3bf == array_addr[14:5] ? valid_959 : _GEN_982; // @[DCache.scala 78:{33,33}]
  wire  _GEN_984 = 10'h3c0 == array_addr[14:5] ? valid_960 : _GEN_983; // @[DCache.scala 78:{33,33}]
  wire  _GEN_985 = 10'h3c1 == array_addr[14:5] ? valid_961 : _GEN_984; // @[DCache.scala 78:{33,33}]
  wire  _GEN_986 = 10'h3c2 == array_addr[14:5] ? valid_962 : _GEN_985; // @[DCache.scala 78:{33,33}]
  wire  _GEN_987 = 10'h3c3 == array_addr[14:5] ? valid_963 : _GEN_986; // @[DCache.scala 78:{33,33}]
  wire  _GEN_988 = 10'h3c4 == array_addr[14:5] ? valid_964 : _GEN_987; // @[DCache.scala 78:{33,33}]
  wire  _GEN_989 = 10'h3c5 == array_addr[14:5] ? valid_965 : _GEN_988; // @[DCache.scala 78:{33,33}]
  wire  _GEN_990 = 10'h3c6 == array_addr[14:5] ? valid_966 : _GEN_989; // @[DCache.scala 78:{33,33}]
  wire  _GEN_991 = 10'h3c7 == array_addr[14:5] ? valid_967 : _GEN_990; // @[DCache.scala 78:{33,33}]
  wire  _GEN_992 = 10'h3c8 == array_addr[14:5] ? valid_968 : _GEN_991; // @[DCache.scala 78:{33,33}]
  wire  _GEN_993 = 10'h3c9 == array_addr[14:5] ? valid_969 : _GEN_992; // @[DCache.scala 78:{33,33}]
  wire  _GEN_994 = 10'h3ca == array_addr[14:5] ? valid_970 : _GEN_993; // @[DCache.scala 78:{33,33}]
  wire  _GEN_995 = 10'h3cb == array_addr[14:5] ? valid_971 : _GEN_994; // @[DCache.scala 78:{33,33}]
  wire  _GEN_996 = 10'h3cc == array_addr[14:5] ? valid_972 : _GEN_995; // @[DCache.scala 78:{33,33}]
  wire  _GEN_997 = 10'h3cd == array_addr[14:5] ? valid_973 : _GEN_996; // @[DCache.scala 78:{33,33}]
  wire  _GEN_998 = 10'h3ce == array_addr[14:5] ? valid_974 : _GEN_997; // @[DCache.scala 78:{33,33}]
  wire  _GEN_999 = 10'h3cf == array_addr[14:5] ? valid_975 : _GEN_998; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1000 = 10'h3d0 == array_addr[14:5] ? valid_976 : _GEN_999; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1001 = 10'h3d1 == array_addr[14:5] ? valid_977 : _GEN_1000; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1002 = 10'h3d2 == array_addr[14:5] ? valid_978 : _GEN_1001; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1003 = 10'h3d3 == array_addr[14:5] ? valid_979 : _GEN_1002; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1004 = 10'h3d4 == array_addr[14:5] ? valid_980 : _GEN_1003; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1005 = 10'h3d5 == array_addr[14:5] ? valid_981 : _GEN_1004; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1006 = 10'h3d6 == array_addr[14:5] ? valid_982 : _GEN_1005; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1007 = 10'h3d7 == array_addr[14:5] ? valid_983 : _GEN_1006; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1008 = 10'h3d8 == array_addr[14:5] ? valid_984 : _GEN_1007; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1009 = 10'h3d9 == array_addr[14:5] ? valid_985 : _GEN_1008; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1010 = 10'h3da == array_addr[14:5] ? valid_986 : _GEN_1009; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1011 = 10'h3db == array_addr[14:5] ? valid_987 : _GEN_1010; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1012 = 10'h3dc == array_addr[14:5] ? valid_988 : _GEN_1011; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1013 = 10'h3dd == array_addr[14:5] ? valid_989 : _GEN_1012; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1014 = 10'h3de == array_addr[14:5] ? valid_990 : _GEN_1013; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1015 = 10'h3df == array_addr[14:5] ? valid_991 : _GEN_1014; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1016 = 10'h3e0 == array_addr[14:5] ? valid_992 : _GEN_1015; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1017 = 10'h3e1 == array_addr[14:5] ? valid_993 : _GEN_1016; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1018 = 10'h3e2 == array_addr[14:5] ? valid_994 : _GEN_1017; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1019 = 10'h3e3 == array_addr[14:5] ? valid_995 : _GEN_1018; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1020 = 10'h3e4 == array_addr[14:5] ? valid_996 : _GEN_1019; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1021 = 10'h3e5 == array_addr[14:5] ? valid_997 : _GEN_1020; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1022 = 10'h3e6 == array_addr[14:5] ? valid_998 : _GEN_1021; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1023 = 10'h3e7 == array_addr[14:5] ? valid_999 : _GEN_1022; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1024 = 10'h3e8 == array_addr[14:5] ? valid_1000 : _GEN_1023; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1025 = 10'h3e9 == array_addr[14:5] ? valid_1001 : _GEN_1024; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1026 = 10'h3ea == array_addr[14:5] ? valid_1002 : _GEN_1025; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1027 = 10'h3eb == array_addr[14:5] ? valid_1003 : _GEN_1026; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1028 = 10'h3ec == array_addr[14:5] ? valid_1004 : _GEN_1027; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1029 = 10'h3ed == array_addr[14:5] ? valid_1005 : _GEN_1028; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1030 = 10'h3ee == array_addr[14:5] ? valid_1006 : _GEN_1029; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1031 = 10'h3ef == array_addr[14:5] ? valid_1007 : _GEN_1030; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1032 = 10'h3f0 == array_addr[14:5] ? valid_1008 : _GEN_1031; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1033 = 10'h3f1 == array_addr[14:5] ? valid_1009 : _GEN_1032; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1034 = 10'h3f2 == array_addr[14:5] ? valid_1010 : _GEN_1033; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1035 = 10'h3f3 == array_addr[14:5] ? valid_1011 : _GEN_1034; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1036 = 10'h3f4 == array_addr[14:5] ? valid_1012 : _GEN_1035; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1037 = 10'h3f5 == array_addr[14:5] ? valid_1013 : _GEN_1036; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1038 = 10'h3f6 == array_addr[14:5] ? valid_1014 : _GEN_1037; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1039 = 10'h3f7 == array_addr[14:5] ? valid_1015 : _GEN_1038; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1040 = 10'h3f8 == array_addr[14:5] ? valid_1016 : _GEN_1039; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1041 = 10'h3f9 == array_addr[14:5] ? valid_1017 : _GEN_1040; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1042 = 10'h3fa == array_addr[14:5] ? valid_1018 : _GEN_1041; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1043 = 10'h3fb == array_addr[14:5] ? valid_1019 : _GEN_1042; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1044 = 10'h3fc == array_addr[14:5] ? valid_1020 : _GEN_1043; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1045 = 10'h3fd == array_addr[14:5] ? valid_1021 : _GEN_1044; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1046 = 10'h3fe == array_addr[14:5] ? valid_1022 : _GEN_1045; // @[DCache.scala 78:{33,33}]
  wire  _GEN_1047 = 10'h3ff == array_addr[14:5] ? valid_1023 : _GEN_1046; // @[DCache.scala 78:{33,33}]
  wire  array_hit = _GEN_1047 & array_wdata_tag == array_out_tag; // @[DCache.scala 78:33]
  reg [26:0] lrsc_addr; // @[DCache.scala 128:30]
  wire  is_lr_r = req_r_lrsc & ~req_r_wen; // @[DCache.scala 131:34]
  wire  _GEN_1048 = _array_io_en_T_1 & is_lr_r | lrsc_reserved; // @[DCache.scala 132:30 133:19 127:30]
  wire [4:0] _lrsc_counter_T_1 = lrsc_counter + 5'h1; // @[DCache.scala 137:34]
  wire  is_sc = io_cache_req_bits_lrsc & io_cache_req_bits_wen; // @[DCache.scala 143:33]
  wire  sc_fail = is_sc & (_x1_b_ready_T_1 | io_cache_req_bits_addr[31:5] != lrsc_addr); // @[DCache.scala 144:25]
  wire  is_sc_r = req_r_lrsc & req_r_wen; // @[DCache.scala 145:30]
  reg  sc_fail_r; // @[Reg.scala 35:20]
  wire [5:0] _sc_rdata_64_T_1 = {req_r_addr[2], 5'h0}; // @[DCache.scala 153:42]
  wire [63:0] _sc_rdata_64_T_2 = 64'h1 << _sc_rdata_64_T_1; // @[DCache.scala 153:24]
  wire [63:0] sc_rdata_64 = sc_fail_r ? _sc_rdata_64_T_2 : 64'h0; // @[DCache.scala 152:19 153:17 151:32]
  wire  _T_12 = ~sc_fail_r; // @[DCache.scala 171:12]
  wire  _GEN_1057 = 10'h0 == array_addr[14:5] | valid_0; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1058 = 10'h1 == array_addr[14:5] | valid_1; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1059 = 10'h2 == array_addr[14:5] | valid_2; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1060 = 10'h3 == array_addr[14:5] | valid_3; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1061 = 10'h4 == array_addr[14:5] | valid_4; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1062 = 10'h5 == array_addr[14:5] | valid_5; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1063 = 10'h6 == array_addr[14:5] | valid_6; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1064 = 10'h7 == array_addr[14:5] | valid_7; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1065 = 10'h8 == array_addr[14:5] | valid_8; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1066 = 10'h9 == array_addr[14:5] | valid_9; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1067 = 10'ha == array_addr[14:5] | valid_10; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1068 = 10'hb == array_addr[14:5] | valid_11; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1069 = 10'hc == array_addr[14:5] | valid_12; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1070 = 10'hd == array_addr[14:5] | valid_13; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1071 = 10'he == array_addr[14:5] | valid_14; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1072 = 10'hf == array_addr[14:5] | valid_15; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1073 = 10'h10 == array_addr[14:5] | valid_16; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1074 = 10'h11 == array_addr[14:5] | valid_17; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1075 = 10'h12 == array_addr[14:5] | valid_18; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1076 = 10'h13 == array_addr[14:5] | valid_19; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1077 = 10'h14 == array_addr[14:5] | valid_20; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1078 = 10'h15 == array_addr[14:5] | valid_21; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1079 = 10'h16 == array_addr[14:5] | valid_22; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1080 = 10'h17 == array_addr[14:5] | valid_23; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1081 = 10'h18 == array_addr[14:5] | valid_24; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1082 = 10'h19 == array_addr[14:5] | valid_25; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1083 = 10'h1a == array_addr[14:5] | valid_26; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1084 = 10'h1b == array_addr[14:5] | valid_27; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1085 = 10'h1c == array_addr[14:5] | valid_28; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1086 = 10'h1d == array_addr[14:5] | valid_29; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1087 = 10'h1e == array_addr[14:5] | valid_30; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1088 = 10'h1f == array_addr[14:5] | valid_31; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1089 = 10'h20 == array_addr[14:5] | valid_32; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1090 = 10'h21 == array_addr[14:5] | valid_33; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1091 = 10'h22 == array_addr[14:5] | valid_34; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1092 = 10'h23 == array_addr[14:5] | valid_35; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1093 = 10'h24 == array_addr[14:5] | valid_36; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1094 = 10'h25 == array_addr[14:5] | valid_37; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1095 = 10'h26 == array_addr[14:5] | valid_38; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1096 = 10'h27 == array_addr[14:5] | valid_39; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1097 = 10'h28 == array_addr[14:5] | valid_40; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1098 = 10'h29 == array_addr[14:5] | valid_41; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1099 = 10'h2a == array_addr[14:5] | valid_42; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1100 = 10'h2b == array_addr[14:5] | valid_43; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1101 = 10'h2c == array_addr[14:5] | valid_44; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1102 = 10'h2d == array_addr[14:5] | valid_45; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1103 = 10'h2e == array_addr[14:5] | valid_46; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1104 = 10'h2f == array_addr[14:5] | valid_47; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1105 = 10'h30 == array_addr[14:5] | valid_48; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1106 = 10'h31 == array_addr[14:5] | valid_49; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1107 = 10'h32 == array_addr[14:5] | valid_50; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1108 = 10'h33 == array_addr[14:5] | valid_51; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1109 = 10'h34 == array_addr[14:5] | valid_52; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1110 = 10'h35 == array_addr[14:5] | valid_53; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1111 = 10'h36 == array_addr[14:5] | valid_54; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1112 = 10'h37 == array_addr[14:5] | valid_55; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1113 = 10'h38 == array_addr[14:5] | valid_56; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1114 = 10'h39 == array_addr[14:5] | valid_57; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1115 = 10'h3a == array_addr[14:5] | valid_58; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1116 = 10'h3b == array_addr[14:5] | valid_59; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1117 = 10'h3c == array_addr[14:5] | valid_60; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1118 = 10'h3d == array_addr[14:5] | valid_61; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1119 = 10'h3e == array_addr[14:5] | valid_62; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1120 = 10'h3f == array_addr[14:5] | valid_63; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1121 = 10'h40 == array_addr[14:5] | valid_64; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1122 = 10'h41 == array_addr[14:5] | valid_65; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1123 = 10'h42 == array_addr[14:5] | valid_66; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1124 = 10'h43 == array_addr[14:5] | valid_67; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1125 = 10'h44 == array_addr[14:5] | valid_68; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1126 = 10'h45 == array_addr[14:5] | valid_69; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1127 = 10'h46 == array_addr[14:5] | valid_70; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1128 = 10'h47 == array_addr[14:5] | valid_71; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1129 = 10'h48 == array_addr[14:5] | valid_72; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1130 = 10'h49 == array_addr[14:5] | valid_73; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1131 = 10'h4a == array_addr[14:5] | valid_74; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1132 = 10'h4b == array_addr[14:5] | valid_75; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1133 = 10'h4c == array_addr[14:5] | valid_76; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1134 = 10'h4d == array_addr[14:5] | valid_77; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1135 = 10'h4e == array_addr[14:5] | valid_78; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1136 = 10'h4f == array_addr[14:5] | valid_79; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1137 = 10'h50 == array_addr[14:5] | valid_80; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1138 = 10'h51 == array_addr[14:5] | valid_81; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1139 = 10'h52 == array_addr[14:5] | valid_82; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1140 = 10'h53 == array_addr[14:5] | valid_83; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1141 = 10'h54 == array_addr[14:5] | valid_84; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1142 = 10'h55 == array_addr[14:5] | valid_85; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1143 = 10'h56 == array_addr[14:5] | valid_86; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1144 = 10'h57 == array_addr[14:5] | valid_87; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1145 = 10'h58 == array_addr[14:5] | valid_88; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1146 = 10'h59 == array_addr[14:5] | valid_89; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1147 = 10'h5a == array_addr[14:5] | valid_90; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1148 = 10'h5b == array_addr[14:5] | valid_91; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1149 = 10'h5c == array_addr[14:5] | valid_92; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1150 = 10'h5d == array_addr[14:5] | valid_93; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1151 = 10'h5e == array_addr[14:5] | valid_94; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1152 = 10'h5f == array_addr[14:5] | valid_95; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1153 = 10'h60 == array_addr[14:5] | valid_96; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1154 = 10'h61 == array_addr[14:5] | valid_97; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1155 = 10'h62 == array_addr[14:5] | valid_98; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1156 = 10'h63 == array_addr[14:5] | valid_99; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1157 = 10'h64 == array_addr[14:5] | valid_100; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1158 = 10'h65 == array_addr[14:5] | valid_101; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1159 = 10'h66 == array_addr[14:5] | valid_102; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1160 = 10'h67 == array_addr[14:5] | valid_103; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1161 = 10'h68 == array_addr[14:5] | valid_104; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1162 = 10'h69 == array_addr[14:5] | valid_105; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1163 = 10'h6a == array_addr[14:5] | valid_106; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1164 = 10'h6b == array_addr[14:5] | valid_107; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1165 = 10'h6c == array_addr[14:5] | valid_108; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1166 = 10'h6d == array_addr[14:5] | valid_109; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1167 = 10'h6e == array_addr[14:5] | valid_110; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1168 = 10'h6f == array_addr[14:5] | valid_111; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1169 = 10'h70 == array_addr[14:5] | valid_112; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1170 = 10'h71 == array_addr[14:5] | valid_113; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1171 = 10'h72 == array_addr[14:5] | valid_114; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1172 = 10'h73 == array_addr[14:5] | valid_115; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1173 = 10'h74 == array_addr[14:5] | valid_116; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1174 = 10'h75 == array_addr[14:5] | valid_117; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1175 = 10'h76 == array_addr[14:5] | valid_118; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1176 = 10'h77 == array_addr[14:5] | valid_119; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1177 = 10'h78 == array_addr[14:5] | valid_120; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1178 = 10'h79 == array_addr[14:5] | valid_121; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1179 = 10'h7a == array_addr[14:5] | valid_122; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1180 = 10'h7b == array_addr[14:5] | valid_123; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1181 = 10'h7c == array_addr[14:5] | valid_124; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1182 = 10'h7d == array_addr[14:5] | valid_125; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1183 = 10'h7e == array_addr[14:5] | valid_126; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1184 = 10'h7f == array_addr[14:5] | valid_127; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1185 = 10'h80 == array_addr[14:5] | valid_128; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1186 = 10'h81 == array_addr[14:5] | valid_129; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1187 = 10'h82 == array_addr[14:5] | valid_130; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1188 = 10'h83 == array_addr[14:5] | valid_131; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1189 = 10'h84 == array_addr[14:5] | valid_132; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1190 = 10'h85 == array_addr[14:5] | valid_133; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1191 = 10'h86 == array_addr[14:5] | valid_134; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1192 = 10'h87 == array_addr[14:5] | valid_135; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1193 = 10'h88 == array_addr[14:5] | valid_136; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1194 = 10'h89 == array_addr[14:5] | valid_137; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1195 = 10'h8a == array_addr[14:5] | valid_138; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1196 = 10'h8b == array_addr[14:5] | valid_139; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1197 = 10'h8c == array_addr[14:5] | valid_140; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1198 = 10'h8d == array_addr[14:5] | valid_141; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1199 = 10'h8e == array_addr[14:5] | valid_142; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1200 = 10'h8f == array_addr[14:5] | valid_143; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1201 = 10'h90 == array_addr[14:5] | valid_144; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1202 = 10'h91 == array_addr[14:5] | valid_145; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1203 = 10'h92 == array_addr[14:5] | valid_146; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1204 = 10'h93 == array_addr[14:5] | valid_147; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1205 = 10'h94 == array_addr[14:5] | valid_148; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1206 = 10'h95 == array_addr[14:5] | valid_149; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1207 = 10'h96 == array_addr[14:5] | valid_150; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1208 = 10'h97 == array_addr[14:5] | valid_151; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1209 = 10'h98 == array_addr[14:5] | valid_152; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1210 = 10'h99 == array_addr[14:5] | valid_153; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1211 = 10'h9a == array_addr[14:5] | valid_154; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1212 = 10'h9b == array_addr[14:5] | valid_155; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1213 = 10'h9c == array_addr[14:5] | valid_156; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1214 = 10'h9d == array_addr[14:5] | valid_157; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1215 = 10'h9e == array_addr[14:5] | valid_158; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1216 = 10'h9f == array_addr[14:5] | valid_159; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1217 = 10'ha0 == array_addr[14:5] | valid_160; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1218 = 10'ha1 == array_addr[14:5] | valid_161; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1219 = 10'ha2 == array_addr[14:5] | valid_162; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1220 = 10'ha3 == array_addr[14:5] | valid_163; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1221 = 10'ha4 == array_addr[14:5] | valid_164; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1222 = 10'ha5 == array_addr[14:5] | valid_165; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1223 = 10'ha6 == array_addr[14:5] | valid_166; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1224 = 10'ha7 == array_addr[14:5] | valid_167; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1225 = 10'ha8 == array_addr[14:5] | valid_168; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1226 = 10'ha9 == array_addr[14:5] | valid_169; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1227 = 10'haa == array_addr[14:5] | valid_170; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1228 = 10'hab == array_addr[14:5] | valid_171; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1229 = 10'hac == array_addr[14:5] | valid_172; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1230 = 10'had == array_addr[14:5] | valid_173; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1231 = 10'hae == array_addr[14:5] | valid_174; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1232 = 10'haf == array_addr[14:5] | valid_175; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1233 = 10'hb0 == array_addr[14:5] | valid_176; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1234 = 10'hb1 == array_addr[14:5] | valid_177; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1235 = 10'hb2 == array_addr[14:5] | valid_178; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1236 = 10'hb3 == array_addr[14:5] | valid_179; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1237 = 10'hb4 == array_addr[14:5] | valid_180; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1238 = 10'hb5 == array_addr[14:5] | valid_181; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1239 = 10'hb6 == array_addr[14:5] | valid_182; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1240 = 10'hb7 == array_addr[14:5] | valid_183; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1241 = 10'hb8 == array_addr[14:5] | valid_184; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1242 = 10'hb9 == array_addr[14:5] | valid_185; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1243 = 10'hba == array_addr[14:5] | valid_186; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1244 = 10'hbb == array_addr[14:5] | valid_187; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1245 = 10'hbc == array_addr[14:5] | valid_188; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1246 = 10'hbd == array_addr[14:5] | valid_189; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1247 = 10'hbe == array_addr[14:5] | valid_190; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1248 = 10'hbf == array_addr[14:5] | valid_191; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1249 = 10'hc0 == array_addr[14:5] | valid_192; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1250 = 10'hc1 == array_addr[14:5] | valid_193; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1251 = 10'hc2 == array_addr[14:5] | valid_194; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1252 = 10'hc3 == array_addr[14:5] | valid_195; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1253 = 10'hc4 == array_addr[14:5] | valid_196; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1254 = 10'hc5 == array_addr[14:5] | valid_197; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1255 = 10'hc6 == array_addr[14:5] | valid_198; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1256 = 10'hc7 == array_addr[14:5] | valid_199; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1257 = 10'hc8 == array_addr[14:5] | valid_200; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1258 = 10'hc9 == array_addr[14:5] | valid_201; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1259 = 10'hca == array_addr[14:5] | valid_202; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1260 = 10'hcb == array_addr[14:5] | valid_203; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1261 = 10'hcc == array_addr[14:5] | valid_204; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1262 = 10'hcd == array_addr[14:5] | valid_205; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1263 = 10'hce == array_addr[14:5] | valid_206; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1264 = 10'hcf == array_addr[14:5] | valid_207; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1265 = 10'hd0 == array_addr[14:5] | valid_208; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1266 = 10'hd1 == array_addr[14:5] | valid_209; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1267 = 10'hd2 == array_addr[14:5] | valid_210; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1268 = 10'hd3 == array_addr[14:5] | valid_211; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1269 = 10'hd4 == array_addr[14:5] | valid_212; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1270 = 10'hd5 == array_addr[14:5] | valid_213; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1271 = 10'hd6 == array_addr[14:5] | valid_214; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1272 = 10'hd7 == array_addr[14:5] | valid_215; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1273 = 10'hd8 == array_addr[14:5] | valid_216; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1274 = 10'hd9 == array_addr[14:5] | valid_217; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1275 = 10'hda == array_addr[14:5] | valid_218; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1276 = 10'hdb == array_addr[14:5] | valid_219; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1277 = 10'hdc == array_addr[14:5] | valid_220; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1278 = 10'hdd == array_addr[14:5] | valid_221; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1279 = 10'hde == array_addr[14:5] | valid_222; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1280 = 10'hdf == array_addr[14:5] | valid_223; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1281 = 10'he0 == array_addr[14:5] | valid_224; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1282 = 10'he1 == array_addr[14:5] | valid_225; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1283 = 10'he2 == array_addr[14:5] | valid_226; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1284 = 10'he3 == array_addr[14:5] | valid_227; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1285 = 10'he4 == array_addr[14:5] | valid_228; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1286 = 10'he5 == array_addr[14:5] | valid_229; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1287 = 10'he6 == array_addr[14:5] | valid_230; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1288 = 10'he7 == array_addr[14:5] | valid_231; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1289 = 10'he8 == array_addr[14:5] | valid_232; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1290 = 10'he9 == array_addr[14:5] | valid_233; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1291 = 10'hea == array_addr[14:5] | valid_234; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1292 = 10'heb == array_addr[14:5] | valid_235; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1293 = 10'hec == array_addr[14:5] | valid_236; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1294 = 10'hed == array_addr[14:5] | valid_237; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1295 = 10'hee == array_addr[14:5] | valid_238; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1296 = 10'hef == array_addr[14:5] | valid_239; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1297 = 10'hf0 == array_addr[14:5] | valid_240; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1298 = 10'hf1 == array_addr[14:5] | valid_241; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1299 = 10'hf2 == array_addr[14:5] | valid_242; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1300 = 10'hf3 == array_addr[14:5] | valid_243; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1301 = 10'hf4 == array_addr[14:5] | valid_244; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1302 = 10'hf5 == array_addr[14:5] | valid_245; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1303 = 10'hf6 == array_addr[14:5] | valid_246; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1304 = 10'hf7 == array_addr[14:5] | valid_247; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1305 = 10'hf8 == array_addr[14:5] | valid_248; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1306 = 10'hf9 == array_addr[14:5] | valid_249; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1307 = 10'hfa == array_addr[14:5] | valid_250; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1308 = 10'hfb == array_addr[14:5] | valid_251; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1309 = 10'hfc == array_addr[14:5] | valid_252; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1310 = 10'hfd == array_addr[14:5] | valid_253; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1311 = 10'hfe == array_addr[14:5] | valid_254; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1312 = 10'hff == array_addr[14:5] | valid_255; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1313 = 10'h100 == array_addr[14:5] | valid_256; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1314 = 10'h101 == array_addr[14:5] | valid_257; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1315 = 10'h102 == array_addr[14:5] | valid_258; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1316 = 10'h103 == array_addr[14:5] | valid_259; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1317 = 10'h104 == array_addr[14:5] | valid_260; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1318 = 10'h105 == array_addr[14:5] | valid_261; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1319 = 10'h106 == array_addr[14:5] | valid_262; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1320 = 10'h107 == array_addr[14:5] | valid_263; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1321 = 10'h108 == array_addr[14:5] | valid_264; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1322 = 10'h109 == array_addr[14:5] | valid_265; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1323 = 10'h10a == array_addr[14:5] | valid_266; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1324 = 10'h10b == array_addr[14:5] | valid_267; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1325 = 10'h10c == array_addr[14:5] | valid_268; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1326 = 10'h10d == array_addr[14:5] | valid_269; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1327 = 10'h10e == array_addr[14:5] | valid_270; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1328 = 10'h10f == array_addr[14:5] | valid_271; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1329 = 10'h110 == array_addr[14:5] | valid_272; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1330 = 10'h111 == array_addr[14:5] | valid_273; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1331 = 10'h112 == array_addr[14:5] | valid_274; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1332 = 10'h113 == array_addr[14:5] | valid_275; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1333 = 10'h114 == array_addr[14:5] | valid_276; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1334 = 10'h115 == array_addr[14:5] | valid_277; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1335 = 10'h116 == array_addr[14:5] | valid_278; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1336 = 10'h117 == array_addr[14:5] | valid_279; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1337 = 10'h118 == array_addr[14:5] | valid_280; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1338 = 10'h119 == array_addr[14:5] | valid_281; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1339 = 10'h11a == array_addr[14:5] | valid_282; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1340 = 10'h11b == array_addr[14:5] | valid_283; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1341 = 10'h11c == array_addr[14:5] | valid_284; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1342 = 10'h11d == array_addr[14:5] | valid_285; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1343 = 10'h11e == array_addr[14:5] | valid_286; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1344 = 10'h11f == array_addr[14:5] | valid_287; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1345 = 10'h120 == array_addr[14:5] | valid_288; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1346 = 10'h121 == array_addr[14:5] | valid_289; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1347 = 10'h122 == array_addr[14:5] | valid_290; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1348 = 10'h123 == array_addr[14:5] | valid_291; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1349 = 10'h124 == array_addr[14:5] | valid_292; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1350 = 10'h125 == array_addr[14:5] | valid_293; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1351 = 10'h126 == array_addr[14:5] | valid_294; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1352 = 10'h127 == array_addr[14:5] | valid_295; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1353 = 10'h128 == array_addr[14:5] | valid_296; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1354 = 10'h129 == array_addr[14:5] | valid_297; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1355 = 10'h12a == array_addr[14:5] | valid_298; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1356 = 10'h12b == array_addr[14:5] | valid_299; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1357 = 10'h12c == array_addr[14:5] | valid_300; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1358 = 10'h12d == array_addr[14:5] | valid_301; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1359 = 10'h12e == array_addr[14:5] | valid_302; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1360 = 10'h12f == array_addr[14:5] | valid_303; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1361 = 10'h130 == array_addr[14:5] | valid_304; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1362 = 10'h131 == array_addr[14:5] | valid_305; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1363 = 10'h132 == array_addr[14:5] | valid_306; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1364 = 10'h133 == array_addr[14:5] | valid_307; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1365 = 10'h134 == array_addr[14:5] | valid_308; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1366 = 10'h135 == array_addr[14:5] | valid_309; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1367 = 10'h136 == array_addr[14:5] | valid_310; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1368 = 10'h137 == array_addr[14:5] | valid_311; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1369 = 10'h138 == array_addr[14:5] | valid_312; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1370 = 10'h139 == array_addr[14:5] | valid_313; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1371 = 10'h13a == array_addr[14:5] | valid_314; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1372 = 10'h13b == array_addr[14:5] | valid_315; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1373 = 10'h13c == array_addr[14:5] | valid_316; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1374 = 10'h13d == array_addr[14:5] | valid_317; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1375 = 10'h13e == array_addr[14:5] | valid_318; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1376 = 10'h13f == array_addr[14:5] | valid_319; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1377 = 10'h140 == array_addr[14:5] | valid_320; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1378 = 10'h141 == array_addr[14:5] | valid_321; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1379 = 10'h142 == array_addr[14:5] | valid_322; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1380 = 10'h143 == array_addr[14:5] | valid_323; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1381 = 10'h144 == array_addr[14:5] | valid_324; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1382 = 10'h145 == array_addr[14:5] | valid_325; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1383 = 10'h146 == array_addr[14:5] | valid_326; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1384 = 10'h147 == array_addr[14:5] | valid_327; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1385 = 10'h148 == array_addr[14:5] | valid_328; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1386 = 10'h149 == array_addr[14:5] | valid_329; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1387 = 10'h14a == array_addr[14:5] | valid_330; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1388 = 10'h14b == array_addr[14:5] | valid_331; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1389 = 10'h14c == array_addr[14:5] | valid_332; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1390 = 10'h14d == array_addr[14:5] | valid_333; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1391 = 10'h14e == array_addr[14:5] | valid_334; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1392 = 10'h14f == array_addr[14:5] | valid_335; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1393 = 10'h150 == array_addr[14:5] | valid_336; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1394 = 10'h151 == array_addr[14:5] | valid_337; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1395 = 10'h152 == array_addr[14:5] | valid_338; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1396 = 10'h153 == array_addr[14:5] | valid_339; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1397 = 10'h154 == array_addr[14:5] | valid_340; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1398 = 10'h155 == array_addr[14:5] | valid_341; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1399 = 10'h156 == array_addr[14:5] | valid_342; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1400 = 10'h157 == array_addr[14:5] | valid_343; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1401 = 10'h158 == array_addr[14:5] | valid_344; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1402 = 10'h159 == array_addr[14:5] | valid_345; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1403 = 10'h15a == array_addr[14:5] | valid_346; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1404 = 10'h15b == array_addr[14:5] | valid_347; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1405 = 10'h15c == array_addr[14:5] | valid_348; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1406 = 10'h15d == array_addr[14:5] | valid_349; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1407 = 10'h15e == array_addr[14:5] | valid_350; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1408 = 10'h15f == array_addr[14:5] | valid_351; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1409 = 10'h160 == array_addr[14:5] | valid_352; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1410 = 10'h161 == array_addr[14:5] | valid_353; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1411 = 10'h162 == array_addr[14:5] | valid_354; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1412 = 10'h163 == array_addr[14:5] | valid_355; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1413 = 10'h164 == array_addr[14:5] | valid_356; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1414 = 10'h165 == array_addr[14:5] | valid_357; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1415 = 10'h166 == array_addr[14:5] | valid_358; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1416 = 10'h167 == array_addr[14:5] | valid_359; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1417 = 10'h168 == array_addr[14:5] | valid_360; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1418 = 10'h169 == array_addr[14:5] | valid_361; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1419 = 10'h16a == array_addr[14:5] | valid_362; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1420 = 10'h16b == array_addr[14:5] | valid_363; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1421 = 10'h16c == array_addr[14:5] | valid_364; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1422 = 10'h16d == array_addr[14:5] | valid_365; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1423 = 10'h16e == array_addr[14:5] | valid_366; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1424 = 10'h16f == array_addr[14:5] | valid_367; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1425 = 10'h170 == array_addr[14:5] | valid_368; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1426 = 10'h171 == array_addr[14:5] | valid_369; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1427 = 10'h172 == array_addr[14:5] | valid_370; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1428 = 10'h173 == array_addr[14:5] | valid_371; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1429 = 10'h174 == array_addr[14:5] | valid_372; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1430 = 10'h175 == array_addr[14:5] | valid_373; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1431 = 10'h176 == array_addr[14:5] | valid_374; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1432 = 10'h177 == array_addr[14:5] | valid_375; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1433 = 10'h178 == array_addr[14:5] | valid_376; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1434 = 10'h179 == array_addr[14:5] | valid_377; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1435 = 10'h17a == array_addr[14:5] | valid_378; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1436 = 10'h17b == array_addr[14:5] | valid_379; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1437 = 10'h17c == array_addr[14:5] | valid_380; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1438 = 10'h17d == array_addr[14:5] | valid_381; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1439 = 10'h17e == array_addr[14:5] | valid_382; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1440 = 10'h17f == array_addr[14:5] | valid_383; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1441 = 10'h180 == array_addr[14:5] | valid_384; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1442 = 10'h181 == array_addr[14:5] | valid_385; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1443 = 10'h182 == array_addr[14:5] | valid_386; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1444 = 10'h183 == array_addr[14:5] | valid_387; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1445 = 10'h184 == array_addr[14:5] | valid_388; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1446 = 10'h185 == array_addr[14:5] | valid_389; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1447 = 10'h186 == array_addr[14:5] | valid_390; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1448 = 10'h187 == array_addr[14:5] | valid_391; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1449 = 10'h188 == array_addr[14:5] | valid_392; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1450 = 10'h189 == array_addr[14:5] | valid_393; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1451 = 10'h18a == array_addr[14:5] | valid_394; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1452 = 10'h18b == array_addr[14:5] | valid_395; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1453 = 10'h18c == array_addr[14:5] | valid_396; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1454 = 10'h18d == array_addr[14:5] | valid_397; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1455 = 10'h18e == array_addr[14:5] | valid_398; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1456 = 10'h18f == array_addr[14:5] | valid_399; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1457 = 10'h190 == array_addr[14:5] | valid_400; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1458 = 10'h191 == array_addr[14:5] | valid_401; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1459 = 10'h192 == array_addr[14:5] | valid_402; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1460 = 10'h193 == array_addr[14:5] | valid_403; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1461 = 10'h194 == array_addr[14:5] | valid_404; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1462 = 10'h195 == array_addr[14:5] | valid_405; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1463 = 10'h196 == array_addr[14:5] | valid_406; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1464 = 10'h197 == array_addr[14:5] | valid_407; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1465 = 10'h198 == array_addr[14:5] | valid_408; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1466 = 10'h199 == array_addr[14:5] | valid_409; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1467 = 10'h19a == array_addr[14:5] | valid_410; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1468 = 10'h19b == array_addr[14:5] | valid_411; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1469 = 10'h19c == array_addr[14:5] | valid_412; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1470 = 10'h19d == array_addr[14:5] | valid_413; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1471 = 10'h19e == array_addr[14:5] | valid_414; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1472 = 10'h19f == array_addr[14:5] | valid_415; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1473 = 10'h1a0 == array_addr[14:5] | valid_416; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1474 = 10'h1a1 == array_addr[14:5] | valid_417; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1475 = 10'h1a2 == array_addr[14:5] | valid_418; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1476 = 10'h1a3 == array_addr[14:5] | valid_419; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1477 = 10'h1a4 == array_addr[14:5] | valid_420; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1478 = 10'h1a5 == array_addr[14:5] | valid_421; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1479 = 10'h1a6 == array_addr[14:5] | valid_422; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1480 = 10'h1a7 == array_addr[14:5] | valid_423; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1481 = 10'h1a8 == array_addr[14:5] | valid_424; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1482 = 10'h1a9 == array_addr[14:5] | valid_425; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1483 = 10'h1aa == array_addr[14:5] | valid_426; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1484 = 10'h1ab == array_addr[14:5] | valid_427; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1485 = 10'h1ac == array_addr[14:5] | valid_428; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1486 = 10'h1ad == array_addr[14:5] | valid_429; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1487 = 10'h1ae == array_addr[14:5] | valid_430; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1488 = 10'h1af == array_addr[14:5] | valid_431; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1489 = 10'h1b0 == array_addr[14:5] | valid_432; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1490 = 10'h1b1 == array_addr[14:5] | valid_433; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1491 = 10'h1b2 == array_addr[14:5] | valid_434; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1492 = 10'h1b3 == array_addr[14:5] | valid_435; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1493 = 10'h1b4 == array_addr[14:5] | valid_436; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1494 = 10'h1b5 == array_addr[14:5] | valid_437; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1495 = 10'h1b6 == array_addr[14:5] | valid_438; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1496 = 10'h1b7 == array_addr[14:5] | valid_439; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1497 = 10'h1b8 == array_addr[14:5] | valid_440; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1498 = 10'h1b9 == array_addr[14:5] | valid_441; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1499 = 10'h1ba == array_addr[14:5] | valid_442; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1500 = 10'h1bb == array_addr[14:5] | valid_443; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1501 = 10'h1bc == array_addr[14:5] | valid_444; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1502 = 10'h1bd == array_addr[14:5] | valid_445; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1503 = 10'h1be == array_addr[14:5] | valid_446; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1504 = 10'h1bf == array_addr[14:5] | valid_447; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1505 = 10'h1c0 == array_addr[14:5] | valid_448; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1506 = 10'h1c1 == array_addr[14:5] | valid_449; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1507 = 10'h1c2 == array_addr[14:5] | valid_450; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1508 = 10'h1c3 == array_addr[14:5] | valid_451; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1509 = 10'h1c4 == array_addr[14:5] | valid_452; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1510 = 10'h1c5 == array_addr[14:5] | valid_453; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1511 = 10'h1c6 == array_addr[14:5] | valid_454; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1512 = 10'h1c7 == array_addr[14:5] | valid_455; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1513 = 10'h1c8 == array_addr[14:5] | valid_456; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1514 = 10'h1c9 == array_addr[14:5] | valid_457; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1515 = 10'h1ca == array_addr[14:5] | valid_458; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1516 = 10'h1cb == array_addr[14:5] | valid_459; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1517 = 10'h1cc == array_addr[14:5] | valid_460; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1518 = 10'h1cd == array_addr[14:5] | valid_461; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1519 = 10'h1ce == array_addr[14:5] | valid_462; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1520 = 10'h1cf == array_addr[14:5] | valid_463; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1521 = 10'h1d0 == array_addr[14:5] | valid_464; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1522 = 10'h1d1 == array_addr[14:5] | valid_465; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1523 = 10'h1d2 == array_addr[14:5] | valid_466; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1524 = 10'h1d3 == array_addr[14:5] | valid_467; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1525 = 10'h1d4 == array_addr[14:5] | valid_468; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1526 = 10'h1d5 == array_addr[14:5] | valid_469; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1527 = 10'h1d6 == array_addr[14:5] | valid_470; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1528 = 10'h1d7 == array_addr[14:5] | valid_471; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1529 = 10'h1d8 == array_addr[14:5] | valid_472; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1530 = 10'h1d9 == array_addr[14:5] | valid_473; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1531 = 10'h1da == array_addr[14:5] | valid_474; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1532 = 10'h1db == array_addr[14:5] | valid_475; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1533 = 10'h1dc == array_addr[14:5] | valid_476; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1534 = 10'h1dd == array_addr[14:5] | valid_477; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1535 = 10'h1de == array_addr[14:5] | valid_478; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1536 = 10'h1df == array_addr[14:5] | valid_479; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1537 = 10'h1e0 == array_addr[14:5] | valid_480; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1538 = 10'h1e1 == array_addr[14:5] | valid_481; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1539 = 10'h1e2 == array_addr[14:5] | valid_482; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1540 = 10'h1e3 == array_addr[14:5] | valid_483; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1541 = 10'h1e4 == array_addr[14:5] | valid_484; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1542 = 10'h1e5 == array_addr[14:5] | valid_485; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1543 = 10'h1e6 == array_addr[14:5] | valid_486; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1544 = 10'h1e7 == array_addr[14:5] | valid_487; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1545 = 10'h1e8 == array_addr[14:5] | valid_488; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1546 = 10'h1e9 == array_addr[14:5] | valid_489; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1547 = 10'h1ea == array_addr[14:5] | valid_490; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1548 = 10'h1eb == array_addr[14:5] | valid_491; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1549 = 10'h1ec == array_addr[14:5] | valid_492; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1550 = 10'h1ed == array_addr[14:5] | valid_493; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1551 = 10'h1ee == array_addr[14:5] | valid_494; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1552 = 10'h1ef == array_addr[14:5] | valid_495; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1553 = 10'h1f0 == array_addr[14:5] | valid_496; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1554 = 10'h1f1 == array_addr[14:5] | valid_497; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1555 = 10'h1f2 == array_addr[14:5] | valid_498; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1556 = 10'h1f3 == array_addr[14:5] | valid_499; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1557 = 10'h1f4 == array_addr[14:5] | valid_500; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1558 = 10'h1f5 == array_addr[14:5] | valid_501; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1559 = 10'h1f6 == array_addr[14:5] | valid_502; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1560 = 10'h1f7 == array_addr[14:5] | valid_503; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1561 = 10'h1f8 == array_addr[14:5] | valid_504; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1562 = 10'h1f9 == array_addr[14:5] | valid_505; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1563 = 10'h1fa == array_addr[14:5] | valid_506; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1564 = 10'h1fb == array_addr[14:5] | valid_507; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1565 = 10'h1fc == array_addr[14:5] | valid_508; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1566 = 10'h1fd == array_addr[14:5] | valid_509; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1567 = 10'h1fe == array_addr[14:5] | valid_510; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1568 = 10'h1ff == array_addr[14:5] | valid_511; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1569 = 10'h200 == array_addr[14:5] | valid_512; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1570 = 10'h201 == array_addr[14:5] | valid_513; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1571 = 10'h202 == array_addr[14:5] | valid_514; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1572 = 10'h203 == array_addr[14:5] | valid_515; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1573 = 10'h204 == array_addr[14:5] | valid_516; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1574 = 10'h205 == array_addr[14:5] | valid_517; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1575 = 10'h206 == array_addr[14:5] | valid_518; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1576 = 10'h207 == array_addr[14:5] | valid_519; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1577 = 10'h208 == array_addr[14:5] | valid_520; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1578 = 10'h209 == array_addr[14:5] | valid_521; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1579 = 10'h20a == array_addr[14:5] | valid_522; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1580 = 10'h20b == array_addr[14:5] | valid_523; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1581 = 10'h20c == array_addr[14:5] | valid_524; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1582 = 10'h20d == array_addr[14:5] | valid_525; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1583 = 10'h20e == array_addr[14:5] | valid_526; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1584 = 10'h20f == array_addr[14:5] | valid_527; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1585 = 10'h210 == array_addr[14:5] | valid_528; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1586 = 10'h211 == array_addr[14:5] | valid_529; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1587 = 10'h212 == array_addr[14:5] | valid_530; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1588 = 10'h213 == array_addr[14:5] | valid_531; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1589 = 10'h214 == array_addr[14:5] | valid_532; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1590 = 10'h215 == array_addr[14:5] | valid_533; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1591 = 10'h216 == array_addr[14:5] | valid_534; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1592 = 10'h217 == array_addr[14:5] | valid_535; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1593 = 10'h218 == array_addr[14:5] | valid_536; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1594 = 10'h219 == array_addr[14:5] | valid_537; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1595 = 10'h21a == array_addr[14:5] | valid_538; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1596 = 10'h21b == array_addr[14:5] | valid_539; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1597 = 10'h21c == array_addr[14:5] | valid_540; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1598 = 10'h21d == array_addr[14:5] | valid_541; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1599 = 10'h21e == array_addr[14:5] | valid_542; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1600 = 10'h21f == array_addr[14:5] | valid_543; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1601 = 10'h220 == array_addr[14:5] | valid_544; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1602 = 10'h221 == array_addr[14:5] | valid_545; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1603 = 10'h222 == array_addr[14:5] | valid_546; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1604 = 10'h223 == array_addr[14:5] | valid_547; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1605 = 10'h224 == array_addr[14:5] | valid_548; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1606 = 10'h225 == array_addr[14:5] | valid_549; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1607 = 10'h226 == array_addr[14:5] | valid_550; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1608 = 10'h227 == array_addr[14:5] | valid_551; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1609 = 10'h228 == array_addr[14:5] | valid_552; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1610 = 10'h229 == array_addr[14:5] | valid_553; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1611 = 10'h22a == array_addr[14:5] | valid_554; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1612 = 10'h22b == array_addr[14:5] | valid_555; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1613 = 10'h22c == array_addr[14:5] | valid_556; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1614 = 10'h22d == array_addr[14:5] | valid_557; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1615 = 10'h22e == array_addr[14:5] | valid_558; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1616 = 10'h22f == array_addr[14:5] | valid_559; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1617 = 10'h230 == array_addr[14:5] | valid_560; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1618 = 10'h231 == array_addr[14:5] | valid_561; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1619 = 10'h232 == array_addr[14:5] | valid_562; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1620 = 10'h233 == array_addr[14:5] | valid_563; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1621 = 10'h234 == array_addr[14:5] | valid_564; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1622 = 10'h235 == array_addr[14:5] | valid_565; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1623 = 10'h236 == array_addr[14:5] | valid_566; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1624 = 10'h237 == array_addr[14:5] | valid_567; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1625 = 10'h238 == array_addr[14:5] | valid_568; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1626 = 10'h239 == array_addr[14:5] | valid_569; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1627 = 10'h23a == array_addr[14:5] | valid_570; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1628 = 10'h23b == array_addr[14:5] | valid_571; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1629 = 10'h23c == array_addr[14:5] | valid_572; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1630 = 10'h23d == array_addr[14:5] | valid_573; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1631 = 10'h23e == array_addr[14:5] | valid_574; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1632 = 10'h23f == array_addr[14:5] | valid_575; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1633 = 10'h240 == array_addr[14:5] | valid_576; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1634 = 10'h241 == array_addr[14:5] | valid_577; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1635 = 10'h242 == array_addr[14:5] | valid_578; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1636 = 10'h243 == array_addr[14:5] | valid_579; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1637 = 10'h244 == array_addr[14:5] | valid_580; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1638 = 10'h245 == array_addr[14:5] | valid_581; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1639 = 10'h246 == array_addr[14:5] | valid_582; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1640 = 10'h247 == array_addr[14:5] | valid_583; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1641 = 10'h248 == array_addr[14:5] | valid_584; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1642 = 10'h249 == array_addr[14:5] | valid_585; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1643 = 10'h24a == array_addr[14:5] | valid_586; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1644 = 10'h24b == array_addr[14:5] | valid_587; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1645 = 10'h24c == array_addr[14:5] | valid_588; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1646 = 10'h24d == array_addr[14:5] | valid_589; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1647 = 10'h24e == array_addr[14:5] | valid_590; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1648 = 10'h24f == array_addr[14:5] | valid_591; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1649 = 10'h250 == array_addr[14:5] | valid_592; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1650 = 10'h251 == array_addr[14:5] | valid_593; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1651 = 10'h252 == array_addr[14:5] | valid_594; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1652 = 10'h253 == array_addr[14:5] | valid_595; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1653 = 10'h254 == array_addr[14:5] | valid_596; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1654 = 10'h255 == array_addr[14:5] | valid_597; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1655 = 10'h256 == array_addr[14:5] | valid_598; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1656 = 10'h257 == array_addr[14:5] | valid_599; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1657 = 10'h258 == array_addr[14:5] | valid_600; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1658 = 10'h259 == array_addr[14:5] | valid_601; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1659 = 10'h25a == array_addr[14:5] | valid_602; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1660 = 10'h25b == array_addr[14:5] | valid_603; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1661 = 10'h25c == array_addr[14:5] | valid_604; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1662 = 10'h25d == array_addr[14:5] | valid_605; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1663 = 10'h25e == array_addr[14:5] | valid_606; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1664 = 10'h25f == array_addr[14:5] | valid_607; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1665 = 10'h260 == array_addr[14:5] | valid_608; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1666 = 10'h261 == array_addr[14:5] | valid_609; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1667 = 10'h262 == array_addr[14:5] | valid_610; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1668 = 10'h263 == array_addr[14:5] | valid_611; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1669 = 10'h264 == array_addr[14:5] | valid_612; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1670 = 10'h265 == array_addr[14:5] | valid_613; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1671 = 10'h266 == array_addr[14:5] | valid_614; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1672 = 10'h267 == array_addr[14:5] | valid_615; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1673 = 10'h268 == array_addr[14:5] | valid_616; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1674 = 10'h269 == array_addr[14:5] | valid_617; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1675 = 10'h26a == array_addr[14:5] | valid_618; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1676 = 10'h26b == array_addr[14:5] | valid_619; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1677 = 10'h26c == array_addr[14:5] | valid_620; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1678 = 10'h26d == array_addr[14:5] | valid_621; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1679 = 10'h26e == array_addr[14:5] | valid_622; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1680 = 10'h26f == array_addr[14:5] | valid_623; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1681 = 10'h270 == array_addr[14:5] | valid_624; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1682 = 10'h271 == array_addr[14:5] | valid_625; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1683 = 10'h272 == array_addr[14:5] | valid_626; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1684 = 10'h273 == array_addr[14:5] | valid_627; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1685 = 10'h274 == array_addr[14:5] | valid_628; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1686 = 10'h275 == array_addr[14:5] | valid_629; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1687 = 10'h276 == array_addr[14:5] | valid_630; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1688 = 10'h277 == array_addr[14:5] | valid_631; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1689 = 10'h278 == array_addr[14:5] | valid_632; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1690 = 10'h279 == array_addr[14:5] | valid_633; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1691 = 10'h27a == array_addr[14:5] | valid_634; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1692 = 10'h27b == array_addr[14:5] | valid_635; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1693 = 10'h27c == array_addr[14:5] | valid_636; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1694 = 10'h27d == array_addr[14:5] | valid_637; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1695 = 10'h27e == array_addr[14:5] | valid_638; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1696 = 10'h27f == array_addr[14:5] | valid_639; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1697 = 10'h280 == array_addr[14:5] | valid_640; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1698 = 10'h281 == array_addr[14:5] | valid_641; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1699 = 10'h282 == array_addr[14:5] | valid_642; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1700 = 10'h283 == array_addr[14:5] | valid_643; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1701 = 10'h284 == array_addr[14:5] | valid_644; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1702 = 10'h285 == array_addr[14:5] | valid_645; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1703 = 10'h286 == array_addr[14:5] | valid_646; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1704 = 10'h287 == array_addr[14:5] | valid_647; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1705 = 10'h288 == array_addr[14:5] | valid_648; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1706 = 10'h289 == array_addr[14:5] | valid_649; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1707 = 10'h28a == array_addr[14:5] | valid_650; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1708 = 10'h28b == array_addr[14:5] | valid_651; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1709 = 10'h28c == array_addr[14:5] | valid_652; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1710 = 10'h28d == array_addr[14:5] | valid_653; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1711 = 10'h28e == array_addr[14:5] | valid_654; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1712 = 10'h28f == array_addr[14:5] | valid_655; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1713 = 10'h290 == array_addr[14:5] | valid_656; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1714 = 10'h291 == array_addr[14:5] | valid_657; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1715 = 10'h292 == array_addr[14:5] | valid_658; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1716 = 10'h293 == array_addr[14:5] | valid_659; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1717 = 10'h294 == array_addr[14:5] | valid_660; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1718 = 10'h295 == array_addr[14:5] | valid_661; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1719 = 10'h296 == array_addr[14:5] | valid_662; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1720 = 10'h297 == array_addr[14:5] | valid_663; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1721 = 10'h298 == array_addr[14:5] | valid_664; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1722 = 10'h299 == array_addr[14:5] | valid_665; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1723 = 10'h29a == array_addr[14:5] | valid_666; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1724 = 10'h29b == array_addr[14:5] | valid_667; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1725 = 10'h29c == array_addr[14:5] | valid_668; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1726 = 10'h29d == array_addr[14:5] | valid_669; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1727 = 10'h29e == array_addr[14:5] | valid_670; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1728 = 10'h29f == array_addr[14:5] | valid_671; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1729 = 10'h2a0 == array_addr[14:5] | valid_672; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1730 = 10'h2a1 == array_addr[14:5] | valid_673; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1731 = 10'h2a2 == array_addr[14:5] | valid_674; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1732 = 10'h2a3 == array_addr[14:5] | valid_675; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1733 = 10'h2a4 == array_addr[14:5] | valid_676; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1734 = 10'h2a5 == array_addr[14:5] | valid_677; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1735 = 10'h2a6 == array_addr[14:5] | valid_678; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1736 = 10'h2a7 == array_addr[14:5] | valid_679; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1737 = 10'h2a8 == array_addr[14:5] | valid_680; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1738 = 10'h2a9 == array_addr[14:5] | valid_681; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1739 = 10'h2aa == array_addr[14:5] | valid_682; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1740 = 10'h2ab == array_addr[14:5] | valid_683; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1741 = 10'h2ac == array_addr[14:5] | valid_684; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1742 = 10'h2ad == array_addr[14:5] | valid_685; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1743 = 10'h2ae == array_addr[14:5] | valid_686; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1744 = 10'h2af == array_addr[14:5] | valid_687; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1745 = 10'h2b0 == array_addr[14:5] | valid_688; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1746 = 10'h2b1 == array_addr[14:5] | valid_689; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1747 = 10'h2b2 == array_addr[14:5] | valid_690; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1748 = 10'h2b3 == array_addr[14:5] | valid_691; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1749 = 10'h2b4 == array_addr[14:5] | valid_692; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1750 = 10'h2b5 == array_addr[14:5] | valid_693; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1751 = 10'h2b6 == array_addr[14:5] | valid_694; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1752 = 10'h2b7 == array_addr[14:5] | valid_695; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1753 = 10'h2b8 == array_addr[14:5] | valid_696; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1754 = 10'h2b9 == array_addr[14:5] | valid_697; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1755 = 10'h2ba == array_addr[14:5] | valid_698; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1756 = 10'h2bb == array_addr[14:5] | valid_699; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1757 = 10'h2bc == array_addr[14:5] | valid_700; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1758 = 10'h2bd == array_addr[14:5] | valid_701; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1759 = 10'h2be == array_addr[14:5] | valid_702; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1760 = 10'h2bf == array_addr[14:5] | valid_703; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1761 = 10'h2c0 == array_addr[14:5] | valid_704; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1762 = 10'h2c1 == array_addr[14:5] | valid_705; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1763 = 10'h2c2 == array_addr[14:5] | valid_706; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1764 = 10'h2c3 == array_addr[14:5] | valid_707; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1765 = 10'h2c4 == array_addr[14:5] | valid_708; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1766 = 10'h2c5 == array_addr[14:5] | valid_709; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1767 = 10'h2c6 == array_addr[14:5] | valid_710; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1768 = 10'h2c7 == array_addr[14:5] | valid_711; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1769 = 10'h2c8 == array_addr[14:5] | valid_712; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1770 = 10'h2c9 == array_addr[14:5] | valid_713; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1771 = 10'h2ca == array_addr[14:5] | valid_714; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1772 = 10'h2cb == array_addr[14:5] | valid_715; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1773 = 10'h2cc == array_addr[14:5] | valid_716; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1774 = 10'h2cd == array_addr[14:5] | valid_717; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1775 = 10'h2ce == array_addr[14:5] | valid_718; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1776 = 10'h2cf == array_addr[14:5] | valid_719; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1777 = 10'h2d0 == array_addr[14:5] | valid_720; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1778 = 10'h2d1 == array_addr[14:5] | valid_721; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1779 = 10'h2d2 == array_addr[14:5] | valid_722; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1780 = 10'h2d3 == array_addr[14:5] | valid_723; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1781 = 10'h2d4 == array_addr[14:5] | valid_724; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1782 = 10'h2d5 == array_addr[14:5] | valid_725; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1783 = 10'h2d6 == array_addr[14:5] | valid_726; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1784 = 10'h2d7 == array_addr[14:5] | valid_727; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1785 = 10'h2d8 == array_addr[14:5] | valid_728; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1786 = 10'h2d9 == array_addr[14:5] | valid_729; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1787 = 10'h2da == array_addr[14:5] | valid_730; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1788 = 10'h2db == array_addr[14:5] | valid_731; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1789 = 10'h2dc == array_addr[14:5] | valid_732; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1790 = 10'h2dd == array_addr[14:5] | valid_733; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1791 = 10'h2de == array_addr[14:5] | valid_734; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1792 = 10'h2df == array_addr[14:5] | valid_735; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1793 = 10'h2e0 == array_addr[14:5] | valid_736; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1794 = 10'h2e1 == array_addr[14:5] | valid_737; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1795 = 10'h2e2 == array_addr[14:5] | valid_738; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1796 = 10'h2e3 == array_addr[14:5] | valid_739; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1797 = 10'h2e4 == array_addr[14:5] | valid_740; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1798 = 10'h2e5 == array_addr[14:5] | valid_741; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1799 = 10'h2e6 == array_addr[14:5] | valid_742; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1800 = 10'h2e7 == array_addr[14:5] | valid_743; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1801 = 10'h2e8 == array_addr[14:5] | valid_744; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1802 = 10'h2e9 == array_addr[14:5] | valid_745; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1803 = 10'h2ea == array_addr[14:5] | valid_746; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1804 = 10'h2eb == array_addr[14:5] | valid_747; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1805 = 10'h2ec == array_addr[14:5] | valid_748; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1806 = 10'h2ed == array_addr[14:5] | valid_749; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1807 = 10'h2ee == array_addr[14:5] | valid_750; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1808 = 10'h2ef == array_addr[14:5] | valid_751; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1809 = 10'h2f0 == array_addr[14:5] | valid_752; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1810 = 10'h2f1 == array_addr[14:5] | valid_753; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1811 = 10'h2f2 == array_addr[14:5] | valid_754; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1812 = 10'h2f3 == array_addr[14:5] | valid_755; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1813 = 10'h2f4 == array_addr[14:5] | valid_756; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1814 = 10'h2f5 == array_addr[14:5] | valid_757; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1815 = 10'h2f6 == array_addr[14:5] | valid_758; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1816 = 10'h2f7 == array_addr[14:5] | valid_759; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1817 = 10'h2f8 == array_addr[14:5] | valid_760; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1818 = 10'h2f9 == array_addr[14:5] | valid_761; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1819 = 10'h2fa == array_addr[14:5] | valid_762; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1820 = 10'h2fb == array_addr[14:5] | valid_763; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1821 = 10'h2fc == array_addr[14:5] | valid_764; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1822 = 10'h2fd == array_addr[14:5] | valid_765; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1823 = 10'h2fe == array_addr[14:5] | valid_766; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1824 = 10'h2ff == array_addr[14:5] | valid_767; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1825 = 10'h300 == array_addr[14:5] | valid_768; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1826 = 10'h301 == array_addr[14:5] | valid_769; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1827 = 10'h302 == array_addr[14:5] | valid_770; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1828 = 10'h303 == array_addr[14:5] | valid_771; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1829 = 10'h304 == array_addr[14:5] | valid_772; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1830 = 10'h305 == array_addr[14:5] | valid_773; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1831 = 10'h306 == array_addr[14:5] | valid_774; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1832 = 10'h307 == array_addr[14:5] | valid_775; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1833 = 10'h308 == array_addr[14:5] | valid_776; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1834 = 10'h309 == array_addr[14:5] | valid_777; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1835 = 10'h30a == array_addr[14:5] | valid_778; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1836 = 10'h30b == array_addr[14:5] | valid_779; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1837 = 10'h30c == array_addr[14:5] | valid_780; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1838 = 10'h30d == array_addr[14:5] | valid_781; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1839 = 10'h30e == array_addr[14:5] | valid_782; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1840 = 10'h30f == array_addr[14:5] | valid_783; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1841 = 10'h310 == array_addr[14:5] | valid_784; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1842 = 10'h311 == array_addr[14:5] | valid_785; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1843 = 10'h312 == array_addr[14:5] | valid_786; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1844 = 10'h313 == array_addr[14:5] | valid_787; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1845 = 10'h314 == array_addr[14:5] | valid_788; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1846 = 10'h315 == array_addr[14:5] | valid_789; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1847 = 10'h316 == array_addr[14:5] | valid_790; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1848 = 10'h317 == array_addr[14:5] | valid_791; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1849 = 10'h318 == array_addr[14:5] | valid_792; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1850 = 10'h319 == array_addr[14:5] | valid_793; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1851 = 10'h31a == array_addr[14:5] | valid_794; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1852 = 10'h31b == array_addr[14:5] | valid_795; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1853 = 10'h31c == array_addr[14:5] | valid_796; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1854 = 10'h31d == array_addr[14:5] | valid_797; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1855 = 10'h31e == array_addr[14:5] | valid_798; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1856 = 10'h31f == array_addr[14:5] | valid_799; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1857 = 10'h320 == array_addr[14:5] | valid_800; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1858 = 10'h321 == array_addr[14:5] | valid_801; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1859 = 10'h322 == array_addr[14:5] | valid_802; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1860 = 10'h323 == array_addr[14:5] | valid_803; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1861 = 10'h324 == array_addr[14:5] | valid_804; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1862 = 10'h325 == array_addr[14:5] | valid_805; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1863 = 10'h326 == array_addr[14:5] | valid_806; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1864 = 10'h327 == array_addr[14:5] | valid_807; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1865 = 10'h328 == array_addr[14:5] | valid_808; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1866 = 10'h329 == array_addr[14:5] | valid_809; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1867 = 10'h32a == array_addr[14:5] | valid_810; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1868 = 10'h32b == array_addr[14:5] | valid_811; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1869 = 10'h32c == array_addr[14:5] | valid_812; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1870 = 10'h32d == array_addr[14:5] | valid_813; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1871 = 10'h32e == array_addr[14:5] | valid_814; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1872 = 10'h32f == array_addr[14:5] | valid_815; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1873 = 10'h330 == array_addr[14:5] | valid_816; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1874 = 10'h331 == array_addr[14:5] | valid_817; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1875 = 10'h332 == array_addr[14:5] | valid_818; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1876 = 10'h333 == array_addr[14:5] | valid_819; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1877 = 10'h334 == array_addr[14:5] | valid_820; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1878 = 10'h335 == array_addr[14:5] | valid_821; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1879 = 10'h336 == array_addr[14:5] | valid_822; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1880 = 10'h337 == array_addr[14:5] | valid_823; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1881 = 10'h338 == array_addr[14:5] | valid_824; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1882 = 10'h339 == array_addr[14:5] | valid_825; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1883 = 10'h33a == array_addr[14:5] | valid_826; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1884 = 10'h33b == array_addr[14:5] | valid_827; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1885 = 10'h33c == array_addr[14:5] | valid_828; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1886 = 10'h33d == array_addr[14:5] | valid_829; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1887 = 10'h33e == array_addr[14:5] | valid_830; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1888 = 10'h33f == array_addr[14:5] | valid_831; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1889 = 10'h340 == array_addr[14:5] | valid_832; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1890 = 10'h341 == array_addr[14:5] | valid_833; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1891 = 10'h342 == array_addr[14:5] | valid_834; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1892 = 10'h343 == array_addr[14:5] | valid_835; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1893 = 10'h344 == array_addr[14:5] | valid_836; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1894 = 10'h345 == array_addr[14:5] | valid_837; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1895 = 10'h346 == array_addr[14:5] | valid_838; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1896 = 10'h347 == array_addr[14:5] | valid_839; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1897 = 10'h348 == array_addr[14:5] | valid_840; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1898 = 10'h349 == array_addr[14:5] | valid_841; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1899 = 10'h34a == array_addr[14:5] | valid_842; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1900 = 10'h34b == array_addr[14:5] | valid_843; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1901 = 10'h34c == array_addr[14:5] | valid_844; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1902 = 10'h34d == array_addr[14:5] | valid_845; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1903 = 10'h34e == array_addr[14:5] | valid_846; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1904 = 10'h34f == array_addr[14:5] | valid_847; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1905 = 10'h350 == array_addr[14:5] | valid_848; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1906 = 10'h351 == array_addr[14:5] | valid_849; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1907 = 10'h352 == array_addr[14:5] | valid_850; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1908 = 10'h353 == array_addr[14:5] | valid_851; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1909 = 10'h354 == array_addr[14:5] | valid_852; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1910 = 10'h355 == array_addr[14:5] | valid_853; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1911 = 10'h356 == array_addr[14:5] | valid_854; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1912 = 10'h357 == array_addr[14:5] | valid_855; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1913 = 10'h358 == array_addr[14:5] | valid_856; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1914 = 10'h359 == array_addr[14:5] | valid_857; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1915 = 10'h35a == array_addr[14:5] | valid_858; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1916 = 10'h35b == array_addr[14:5] | valid_859; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1917 = 10'h35c == array_addr[14:5] | valid_860; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1918 = 10'h35d == array_addr[14:5] | valid_861; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1919 = 10'h35e == array_addr[14:5] | valid_862; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1920 = 10'h35f == array_addr[14:5] | valid_863; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1921 = 10'h360 == array_addr[14:5] | valid_864; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1922 = 10'h361 == array_addr[14:5] | valid_865; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1923 = 10'h362 == array_addr[14:5] | valid_866; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1924 = 10'h363 == array_addr[14:5] | valid_867; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1925 = 10'h364 == array_addr[14:5] | valid_868; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1926 = 10'h365 == array_addr[14:5] | valid_869; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1927 = 10'h366 == array_addr[14:5] | valid_870; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1928 = 10'h367 == array_addr[14:5] | valid_871; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1929 = 10'h368 == array_addr[14:5] | valid_872; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1930 = 10'h369 == array_addr[14:5] | valid_873; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1931 = 10'h36a == array_addr[14:5] | valid_874; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1932 = 10'h36b == array_addr[14:5] | valid_875; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1933 = 10'h36c == array_addr[14:5] | valid_876; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1934 = 10'h36d == array_addr[14:5] | valid_877; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1935 = 10'h36e == array_addr[14:5] | valid_878; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1936 = 10'h36f == array_addr[14:5] | valid_879; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1937 = 10'h370 == array_addr[14:5] | valid_880; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1938 = 10'h371 == array_addr[14:5] | valid_881; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1939 = 10'h372 == array_addr[14:5] | valid_882; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1940 = 10'h373 == array_addr[14:5] | valid_883; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1941 = 10'h374 == array_addr[14:5] | valid_884; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1942 = 10'h375 == array_addr[14:5] | valid_885; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1943 = 10'h376 == array_addr[14:5] | valid_886; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1944 = 10'h377 == array_addr[14:5] | valid_887; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1945 = 10'h378 == array_addr[14:5] | valid_888; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1946 = 10'h379 == array_addr[14:5] | valid_889; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1947 = 10'h37a == array_addr[14:5] | valid_890; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1948 = 10'h37b == array_addr[14:5] | valid_891; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1949 = 10'h37c == array_addr[14:5] | valid_892; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1950 = 10'h37d == array_addr[14:5] | valid_893; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1951 = 10'h37e == array_addr[14:5] | valid_894; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1952 = 10'h37f == array_addr[14:5] | valid_895; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1953 = 10'h380 == array_addr[14:5] | valid_896; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1954 = 10'h381 == array_addr[14:5] | valid_897; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1955 = 10'h382 == array_addr[14:5] | valid_898; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1956 = 10'h383 == array_addr[14:5] | valid_899; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1957 = 10'h384 == array_addr[14:5] | valid_900; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1958 = 10'h385 == array_addr[14:5] | valid_901; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1959 = 10'h386 == array_addr[14:5] | valid_902; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1960 = 10'h387 == array_addr[14:5] | valid_903; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1961 = 10'h388 == array_addr[14:5] | valid_904; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1962 = 10'h389 == array_addr[14:5] | valid_905; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1963 = 10'h38a == array_addr[14:5] | valid_906; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1964 = 10'h38b == array_addr[14:5] | valid_907; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1965 = 10'h38c == array_addr[14:5] | valid_908; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1966 = 10'h38d == array_addr[14:5] | valid_909; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1967 = 10'h38e == array_addr[14:5] | valid_910; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1968 = 10'h38f == array_addr[14:5] | valid_911; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1969 = 10'h390 == array_addr[14:5] | valid_912; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1970 = 10'h391 == array_addr[14:5] | valid_913; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1971 = 10'h392 == array_addr[14:5] | valid_914; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1972 = 10'h393 == array_addr[14:5] | valid_915; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1973 = 10'h394 == array_addr[14:5] | valid_916; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1974 = 10'h395 == array_addr[14:5] | valid_917; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1975 = 10'h396 == array_addr[14:5] | valid_918; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1976 = 10'h397 == array_addr[14:5] | valid_919; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1977 = 10'h398 == array_addr[14:5] | valid_920; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1978 = 10'h399 == array_addr[14:5] | valid_921; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1979 = 10'h39a == array_addr[14:5] | valid_922; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1980 = 10'h39b == array_addr[14:5] | valid_923; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1981 = 10'h39c == array_addr[14:5] | valid_924; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1982 = 10'h39d == array_addr[14:5] | valid_925; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1983 = 10'h39e == array_addr[14:5] | valid_926; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1984 = 10'h39f == array_addr[14:5] | valid_927; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1985 = 10'h3a0 == array_addr[14:5] | valid_928; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1986 = 10'h3a1 == array_addr[14:5] | valid_929; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1987 = 10'h3a2 == array_addr[14:5] | valid_930; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1988 = 10'h3a3 == array_addr[14:5] | valid_931; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1989 = 10'h3a4 == array_addr[14:5] | valid_932; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1990 = 10'h3a5 == array_addr[14:5] | valid_933; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1991 = 10'h3a6 == array_addr[14:5] | valid_934; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1992 = 10'h3a7 == array_addr[14:5] | valid_935; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1993 = 10'h3a8 == array_addr[14:5] | valid_936; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1994 = 10'h3a9 == array_addr[14:5] | valid_937; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1995 = 10'h3aa == array_addr[14:5] | valid_938; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1996 = 10'h3ab == array_addr[14:5] | valid_939; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1997 = 10'h3ac == array_addr[14:5] | valid_940; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1998 = 10'h3ad == array_addr[14:5] | valid_941; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_1999 = 10'h3ae == array_addr[14:5] | valid_942; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2000 = 10'h3af == array_addr[14:5] | valid_943; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2001 = 10'h3b0 == array_addr[14:5] | valid_944; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2002 = 10'h3b1 == array_addr[14:5] | valid_945; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2003 = 10'h3b2 == array_addr[14:5] | valid_946; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2004 = 10'h3b3 == array_addr[14:5] | valid_947; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2005 = 10'h3b4 == array_addr[14:5] | valid_948; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2006 = 10'h3b5 == array_addr[14:5] | valid_949; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2007 = 10'h3b6 == array_addr[14:5] | valid_950; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2008 = 10'h3b7 == array_addr[14:5] | valid_951; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2009 = 10'h3b8 == array_addr[14:5] | valid_952; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2010 = 10'h3b9 == array_addr[14:5] | valid_953; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2011 = 10'h3ba == array_addr[14:5] | valid_954; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2012 = 10'h3bb == array_addr[14:5] | valid_955; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2013 = 10'h3bc == array_addr[14:5] | valid_956; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2014 = 10'h3bd == array_addr[14:5] | valid_957; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2015 = 10'h3be == array_addr[14:5] | valid_958; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2016 = 10'h3bf == array_addr[14:5] | valid_959; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2017 = 10'h3c0 == array_addr[14:5] | valid_960; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2018 = 10'h3c1 == array_addr[14:5] | valid_961; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2019 = 10'h3c2 == array_addr[14:5] | valid_962; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2020 = 10'h3c3 == array_addr[14:5] | valid_963; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2021 = 10'h3c4 == array_addr[14:5] | valid_964; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2022 = 10'h3c5 == array_addr[14:5] | valid_965; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2023 = 10'h3c6 == array_addr[14:5] | valid_966; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2024 = 10'h3c7 == array_addr[14:5] | valid_967; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2025 = 10'h3c8 == array_addr[14:5] | valid_968; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2026 = 10'h3c9 == array_addr[14:5] | valid_969; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2027 = 10'h3ca == array_addr[14:5] | valid_970; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2028 = 10'h3cb == array_addr[14:5] | valid_971; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2029 = 10'h3cc == array_addr[14:5] | valid_972; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2030 = 10'h3cd == array_addr[14:5] | valid_973; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2031 = 10'h3ce == array_addr[14:5] | valid_974; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2032 = 10'h3cf == array_addr[14:5] | valid_975; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2033 = 10'h3d0 == array_addr[14:5] | valid_976; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2034 = 10'h3d1 == array_addr[14:5] | valid_977; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2035 = 10'h3d2 == array_addr[14:5] | valid_978; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2036 = 10'h3d3 == array_addr[14:5] | valid_979; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2037 = 10'h3d4 == array_addr[14:5] | valid_980; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2038 = 10'h3d5 == array_addr[14:5] | valid_981; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2039 = 10'h3d6 == array_addr[14:5] | valid_982; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2040 = 10'h3d7 == array_addr[14:5] | valid_983; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2041 = 10'h3d8 == array_addr[14:5] | valid_984; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2042 = 10'h3d9 == array_addr[14:5] | valid_985; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2043 = 10'h3da == array_addr[14:5] | valid_986; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2044 = 10'h3db == array_addr[14:5] | valid_987; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2045 = 10'h3dc == array_addr[14:5] | valid_988; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2046 = 10'h3dd == array_addr[14:5] | valid_989; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2047 = 10'h3de == array_addr[14:5] | valid_990; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2048 = 10'h3df == array_addr[14:5] | valid_991; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2049 = 10'h3e0 == array_addr[14:5] | valid_992; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2050 = 10'h3e1 == array_addr[14:5] | valid_993; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2051 = 10'h3e2 == array_addr[14:5] | valid_994; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2052 = 10'h3e3 == array_addr[14:5] | valid_995; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2053 = 10'h3e4 == array_addr[14:5] | valid_996; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2054 = 10'h3e5 == array_addr[14:5] | valid_997; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2055 = 10'h3e6 == array_addr[14:5] | valid_998; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2056 = 10'h3e7 == array_addr[14:5] | valid_999; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2057 = 10'h3e8 == array_addr[14:5] | valid_1000; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2058 = 10'h3e9 == array_addr[14:5] | valid_1001; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2059 = 10'h3ea == array_addr[14:5] | valid_1002; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2060 = 10'h3eb == array_addr[14:5] | valid_1003; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2061 = 10'h3ec == array_addr[14:5] | valid_1004; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2062 = 10'h3ed == array_addr[14:5] | valid_1005; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2063 = 10'h3ee == array_addr[14:5] | valid_1006; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2064 = 10'h3ef == array_addr[14:5] | valid_1007; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2065 = 10'h3f0 == array_addr[14:5] | valid_1008; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2066 = 10'h3f1 == array_addr[14:5] | valid_1009; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2067 = 10'h3f2 == array_addr[14:5] | valid_1010; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2068 = 10'h3f3 == array_addr[14:5] | valid_1011; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2069 = 10'h3f4 == array_addr[14:5] | valid_1012; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2070 = 10'h3f5 == array_addr[14:5] | valid_1013; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2071 = 10'h3f6 == array_addr[14:5] | valid_1014; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2072 = 10'h3f7 == array_addr[14:5] | valid_1015; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2073 = 10'h3f8 == array_addr[14:5] | valid_1016; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2074 = 10'h3f9 == array_addr[14:5] | valid_1017; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2075 = 10'h3fa == array_addr[14:5] | valid_1018; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2076 = 10'h3fb == array_addr[14:5] | valid_1019; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2077 = 10'h3fc == array_addr[14:5] | valid_1020; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2078 = 10'h3fd == array_addr[14:5] | valid_1021; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2079 = 10'h3fe == array_addr[14:5] | valid_1022; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2080 = 10'h3ff == array_addr[14:5] | valid_1023; // @[DCache.scala 173:{37,37} 56:22]
  wire  _GEN_2082 = ~sc_fail_r ? _GEN_1057 : valid_0; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2083 = ~sc_fail_r ? _GEN_1058 : valid_1; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2084 = ~sc_fail_r ? _GEN_1059 : valid_2; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2085 = ~sc_fail_r ? _GEN_1060 : valid_3; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2086 = ~sc_fail_r ? _GEN_1061 : valid_4; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2087 = ~sc_fail_r ? _GEN_1062 : valid_5; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2088 = ~sc_fail_r ? _GEN_1063 : valid_6; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2089 = ~sc_fail_r ? _GEN_1064 : valid_7; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2090 = ~sc_fail_r ? _GEN_1065 : valid_8; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2091 = ~sc_fail_r ? _GEN_1066 : valid_9; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2092 = ~sc_fail_r ? _GEN_1067 : valid_10; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2093 = ~sc_fail_r ? _GEN_1068 : valid_11; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2094 = ~sc_fail_r ? _GEN_1069 : valid_12; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2095 = ~sc_fail_r ? _GEN_1070 : valid_13; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2096 = ~sc_fail_r ? _GEN_1071 : valid_14; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2097 = ~sc_fail_r ? _GEN_1072 : valid_15; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2098 = ~sc_fail_r ? _GEN_1073 : valid_16; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2099 = ~sc_fail_r ? _GEN_1074 : valid_17; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2100 = ~sc_fail_r ? _GEN_1075 : valid_18; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2101 = ~sc_fail_r ? _GEN_1076 : valid_19; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2102 = ~sc_fail_r ? _GEN_1077 : valid_20; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2103 = ~sc_fail_r ? _GEN_1078 : valid_21; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2104 = ~sc_fail_r ? _GEN_1079 : valid_22; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2105 = ~sc_fail_r ? _GEN_1080 : valid_23; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2106 = ~sc_fail_r ? _GEN_1081 : valid_24; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2107 = ~sc_fail_r ? _GEN_1082 : valid_25; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2108 = ~sc_fail_r ? _GEN_1083 : valid_26; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2109 = ~sc_fail_r ? _GEN_1084 : valid_27; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2110 = ~sc_fail_r ? _GEN_1085 : valid_28; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2111 = ~sc_fail_r ? _GEN_1086 : valid_29; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2112 = ~sc_fail_r ? _GEN_1087 : valid_30; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2113 = ~sc_fail_r ? _GEN_1088 : valid_31; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2114 = ~sc_fail_r ? _GEN_1089 : valid_32; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2115 = ~sc_fail_r ? _GEN_1090 : valid_33; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2116 = ~sc_fail_r ? _GEN_1091 : valid_34; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2117 = ~sc_fail_r ? _GEN_1092 : valid_35; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2118 = ~sc_fail_r ? _GEN_1093 : valid_36; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2119 = ~sc_fail_r ? _GEN_1094 : valid_37; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2120 = ~sc_fail_r ? _GEN_1095 : valid_38; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2121 = ~sc_fail_r ? _GEN_1096 : valid_39; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2122 = ~sc_fail_r ? _GEN_1097 : valid_40; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2123 = ~sc_fail_r ? _GEN_1098 : valid_41; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2124 = ~sc_fail_r ? _GEN_1099 : valid_42; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2125 = ~sc_fail_r ? _GEN_1100 : valid_43; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2126 = ~sc_fail_r ? _GEN_1101 : valid_44; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2127 = ~sc_fail_r ? _GEN_1102 : valid_45; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2128 = ~sc_fail_r ? _GEN_1103 : valid_46; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2129 = ~sc_fail_r ? _GEN_1104 : valid_47; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2130 = ~sc_fail_r ? _GEN_1105 : valid_48; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2131 = ~sc_fail_r ? _GEN_1106 : valid_49; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2132 = ~sc_fail_r ? _GEN_1107 : valid_50; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2133 = ~sc_fail_r ? _GEN_1108 : valid_51; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2134 = ~sc_fail_r ? _GEN_1109 : valid_52; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2135 = ~sc_fail_r ? _GEN_1110 : valid_53; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2136 = ~sc_fail_r ? _GEN_1111 : valid_54; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2137 = ~sc_fail_r ? _GEN_1112 : valid_55; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2138 = ~sc_fail_r ? _GEN_1113 : valid_56; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2139 = ~sc_fail_r ? _GEN_1114 : valid_57; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2140 = ~sc_fail_r ? _GEN_1115 : valid_58; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2141 = ~sc_fail_r ? _GEN_1116 : valid_59; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2142 = ~sc_fail_r ? _GEN_1117 : valid_60; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2143 = ~sc_fail_r ? _GEN_1118 : valid_61; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2144 = ~sc_fail_r ? _GEN_1119 : valid_62; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2145 = ~sc_fail_r ? _GEN_1120 : valid_63; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2146 = ~sc_fail_r ? _GEN_1121 : valid_64; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2147 = ~sc_fail_r ? _GEN_1122 : valid_65; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2148 = ~sc_fail_r ? _GEN_1123 : valid_66; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2149 = ~sc_fail_r ? _GEN_1124 : valid_67; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2150 = ~sc_fail_r ? _GEN_1125 : valid_68; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2151 = ~sc_fail_r ? _GEN_1126 : valid_69; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2152 = ~sc_fail_r ? _GEN_1127 : valid_70; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2153 = ~sc_fail_r ? _GEN_1128 : valid_71; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2154 = ~sc_fail_r ? _GEN_1129 : valid_72; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2155 = ~sc_fail_r ? _GEN_1130 : valid_73; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2156 = ~sc_fail_r ? _GEN_1131 : valid_74; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2157 = ~sc_fail_r ? _GEN_1132 : valid_75; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2158 = ~sc_fail_r ? _GEN_1133 : valid_76; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2159 = ~sc_fail_r ? _GEN_1134 : valid_77; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2160 = ~sc_fail_r ? _GEN_1135 : valid_78; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2161 = ~sc_fail_r ? _GEN_1136 : valid_79; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2162 = ~sc_fail_r ? _GEN_1137 : valid_80; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2163 = ~sc_fail_r ? _GEN_1138 : valid_81; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2164 = ~sc_fail_r ? _GEN_1139 : valid_82; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2165 = ~sc_fail_r ? _GEN_1140 : valid_83; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2166 = ~sc_fail_r ? _GEN_1141 : valid_84; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2167 = ~sc_fail_r ? _GEN_1142 : valid_85; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2168 = ~sc_fail_r ? _GEN_1143 : valid_86; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2169 = ~sc_fail_r ? _GEN_1144 : valid_87; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2170 = ~sc_fail_r ? _GEN_1145 : valid_88; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2171 = ~sc_fail_r ? _GEN_1146 : valid_89; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2172 = ~sc_fail_r ? _GEN_1147 : valid_90; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2173 = ~sc_fail_r ? _GEN_1148 : valid_91; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2174 = ~sc_fail_r ? _GEN_1149 : valid_92; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2175 = ~sc_fail_r ? _GEN_1150 : valid_93; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2176 = ~sc_fail_r ? _GEN_1151 : valid_94; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2177 = ~sc_fail_r ? _GEN_1152 : valid_95; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2178 = ~sc_fail_r ? _GEN_1153 : valid_96; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2179 = ~sc_fail_r ? _GEN_1154 : valid_97; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2180 = ~sc_fail_r ? _GEN_1155 : valid_98; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2181 = ~sc_fail_r ? _GEN_1156 : valid_99; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2182 = ~sc_fail_r ? _GEN_1157 : valid_100; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2183 = ~sc_fail_r ? _GEN_1158 : valid_101; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2184 = ~sc_fail_r ? _GEN_1159 : valid_102; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2185 = ~sc_fail_r ? _GEN_1160 : valid_103; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2186 = ~sc_fail_r ? _GEN_1161 : valid_104; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2187 = ~sc_fail_r ? _GEN_1162 : valid_105; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2188 = ~sc_fail_r ? _GEN_1163 : valid_106; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2189 = ~sc_fail_r ? _GEN_1164 : valid_107; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2190 = ~sc_fail_r ? _GEN_1165 : valid_108; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2191 = ~sc_fail_r ? _GEN_1166 : valid_109; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2192 = ~sc_fail_r ? _GEN_1167 : valid_110; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2193 = ~sc_fail_r ? _GEN_1168 : valid_111; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2194 = ~sc_fail_r ? _GEN_1169 : valid_112; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2195 = ~sc_fail_r ? _GEN_1170 : valid_113; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2196 = ~sc_fail_r ? _GEN_1171 : valid_114; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2197 = ~sc_fail_r ? _GEN_1172 : valid_115; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2198 = ~sc_fail_r ? _GEN_1173 : valid_116; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2199 = ~sc_fail_r ? _GEN_1174 : valid_117; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2200 = ~sc_fail_r ? _GEN_1175 : valid_118; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2201 = ~sc_fail_r ? _GEN_1176 : valid_119; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2202 = ~sc_fail_r ? _GEN_1177 : valid_120; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2203 = ~sc_fail_r ? _GEN_1178 : valid_121; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2204 = ~sc_fail_r ? _GEN_1179 : valid_122; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2205 = ~sc_fail_r ? _GEN_1180 : valid_123; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2206 = ~sc_fail_r ? _GEN_1181 : valid_124; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2207 = ~sc_fail_r ? _GEN_1182 : valid_125; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2208 = ~sc_fail_r ? _GEN_1183 : valid_126; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2209 = ~sc_fail_r ? _GEN_1184 : valid_127; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2210 = ~sc_fail_r ? _GEN_1185 : valid_128; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2211 = ~sc_fail_r ? _GEN_1186 : valid_129; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2212 = ~sc_fail_r ? _GEN_1187 : valid_130; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2213 = ~sc_fail_r ? _GEN_1188 : valid_131; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2214 = ~sc_fail_r ? _GEN_1189 : valid_132; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2215 = ~sc_fail_r ? _GEN_1190 : valid_133; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2216 = ~sc_fail_r ? _GEN_1191 : valid_134; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2217 = ~sc_fail_r ? _GEN_1192 : valid_135; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2218 = ~sc_fail_r ? _GEN_1193 : valid_136; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2219 = ~sc_fail_r ? _GEN_1194 : valid_137; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2220 = ~sc_fail_r ? _GEN_1195 : valid_138; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2221 = ~sc_fail_r ? _GEN_1196 : valid_139; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2222 = ~sc_fail_r ? _GEN_1197 : valid_140; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2223 = ~sc_fail_r ? _GEN_1198 : valid_141; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2224 = ~sc_fail_r ? _GEN_1199 : valid_142; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2225 = ~sc_fail_r ? _GEN_1200 : valid_143; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2226 = ~sc_fail_r ? _GEN_1201 : valid_144; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2227 = ~sc_fail_r ? _GEN_1202 : valid_145; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2228 = ~sc_fail_r ? _GEN_1203 : valid_146; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2229 = ~sc_fail_r ? _GEN_1204 : valid_147; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2230 = ~sc_fail_r ? _GEN_1205 : valid_148; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2231 = ~sc_fail_r ? _GEN_1206 : valid_149; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2232 = ~sc_fail_r ? _GEN_1207 : valid_150; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2233 = ~sc_fail_r ? _GEN_1208 : valid_151; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2234 = ~sc_fail_r ? _GEN_1209 : valid_152; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2235 = ~sc_fail_r ? _GEN_1210 : valid_153; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2236 = ~sc_fail_r ? _GEN_1211 : valid_154; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2237 = ~sc_fail_r ? _GEN_1212 : valid_155; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2238 = ~sc_fail_r ? _GEN_1213 : valid_156; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2239 = ~sc_fail_r ? _GEN_1214 : valid_157; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2240 = ~sc_fail_r ? _GEN_1215 : valid_158; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2241 = ~sc_fail_r ? _GEN_1216 : valid_159; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2242 = ~sc_fail_r ? _GEN_1217 : valid_160; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2243 = ~sc_fail_r ? _GEN_1218 : valid_161; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2244 = ~sc_fail_r ? _GEN_1219 : valid_162; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2245 = ~sc_fail_r ? _GEN_1220 : valid_163; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2246 = ~sc_fail_r ? _GEN_1221 : valid_164; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2247 = ~sc_fail_r ? _GEN_1222 : valid_165; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2248 = ~sc_fail_r ? _GEN_1223 : valid_166; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2249 = ~sc_fail_r ? _GEN_1224 : valid_167; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2250 = ~sc_fail_r ? _GEN_1225 : valid_168; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2251 = ~sc_fail_r ? _GEN_1226 : valid_169; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2252 = ~sc_fail_r ? _GEN_1227 : valid_170; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2253 = ~sc_fail_r ? _GEN_1228 : valid_171; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2254 = ~sc_fail_r ? _GEN_1229 : valid_172; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2255 = ~sc_fail_r ? _GEN_1230 : valid_173; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2256 = ~sc_fail_r ? _GEN_1231 : valid_174; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2257 = ~sc_fail_r ? _GEN_1232 : valid_175; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2258 = ~sc_fail_r ? _GEN_1233 : valid_176; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2259 = ~sc_fail_r ? _GEN_1234 : valid_177; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2260 = ~sc_fail_r ? _GEN_1235 : valid_178; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2261 = ~sc_fail_r ? _GEN_1236 : valid_179; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2262 = ~sc_fail_r ? _GEN_1237 : valid_180; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2263 = ~sc_fail_r ? _GEN_1238 : valid_181; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2264 = ~sc_fail_r ? _GEN_1239 : valid_182; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2265 = ~sc_fail_r ? _GEN_1240 : valid_183; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2266 = ~sc_fail_r ? _GEN_1241 : valid_184; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2267 = ~sc_fail_r ? _GEN_1242 : valid_185; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2268 = ~sc_fail_r ? _GEN_1243 : valid_186; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2269 = ~sc_fail_r ? _GEN_1244 : valid_187; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2270 = ~sc_fail_r ? _GEN_1245 : valid_188; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2271 = ~sc_fail_r ? _GEN_1246 : valid_189; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2272 = ~sc_fail_r ? _GEN_1247 : valid_190; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2273 = ~sc_fail_r ? _GEN_1248 : valid_191; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2274 = ~sc_fail_r ? _GEN_1249 : valid_192; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2275 = ~sc_fail_r ? _GEN_1250 : valid_193; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2276 = ~sc_fail_r ? _GEN_1251 : valid_194; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2277 = ~sc_fail_r ? _GEN_1252 : valid_195; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2278 = ~sc_fail_r ? _GEN_1253 : valid_196; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2279 = ~sc_fail_r ? _GEN_1254 : valid_197; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2280 = ~sc_fail_r ? _GEN_1255 : valid_198; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2281 = ~sc_fail_r ? _GEN_1256 : valid_199; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2282 = ~sc_fail_r ? _GEN_1257 : valid_200; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2283 = ~sc_fail_r ? _GEN_1258 : valid_201; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2284 = ~sc_fail_r ? _GEN_1259 : valid_202; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2285 = ~sc_fail_r ? _GEN_1260 : valid_203; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2286 = ~sc_fail_r ? _GEN_1261 : valid_204; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2287 = ~sc_fail_r ? _GEN_1262 : valid_205; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2288 = ~sc_fail_r ? _GEN_1263 : valid_206; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2289 = ~sc_fail_r ? _GEN_1264 : valid_207; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2290 = ~sc_fail_r ? _GEN_1265 : valid_208; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2291 = ~sc_fail_r ? _GEN_1266 : valid_209; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2292 = ~sc_fail_r ? _GEN_1267 : valid_210; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2293 = ~sc_fail_r ? _GEN_1268 : valid_211; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2294 = ~sc_fail_r ? _GEN_1269 : valid_212; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2295 = ~sc_fail_r ? _GEN_1270 : valid_213; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2296 = ~sc_fail_r ? _GEN_1271 : valid_214; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2297 = ~sc_fail_r ? _GEN_1272 : valid_215; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2298 = ~sc_fail_r ? _GEN_1273 : valid_216; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2299 = ~sc_fail_r ? _GEN_1274 : valid_217; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2300 = ~sc_fail_r ? _GEN_1275 : valid_218; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2301 = ~sc_fail_r ? _GEN_1276 : valid_219; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2302 = ~sc_fail_r ? _GEN_1277 : valid_220; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2303 = ~sc_fail_r ? _GEN_1278 : valid_221; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2304 = ~sc_fail_r ? _GEN_1279 : valid_222; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2305 = ~sc_fail_r ? _GEN_1280 : valid_223; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2306 = ~sc_fail_r ? _GEN_1281 : valid_224; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2307 = ~sc_fail_r ? _GEN_1282 : valid_225; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2308 = ~sc_fail_r ? _GEN_1283 : valid_226; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2309 = ~sc_fail_r ? _GEN_1284 : valid_227; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2310 = ~sc_fail_r ? _GEN_1285 : valid_228; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2311 = ~sc_fail_r ? _GEN_1286 : valid_229; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2312 = ~sc_fail_r ? _GEN_1287 : valid_230; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2313 = ~sc_fail_r ? _GEN_1288 : valid_231; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2314 = ~sc_fail_r ? _GEN_1289 : valid_232; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2315 = ~sc_fail_r ? _GEN_1290 : valid_233; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2316 = ~sc_fail_r ? _GEN_1291 : valid_234; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2317 = ~sc_fail_r ? _GEN_1292 : valid_235; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2318 = ~sc_fail_r ? _GEN_1293 : valid_236; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2319 = ~sc_fail_r ? _GEN_1294 : valid_237; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2320 = ~sc_fail_r ? _GEN_1295 : valid_238; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2321 = ~sc_fail_r ? _GEN_1296 : valid_239; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2322 = ~sc_fail_r ? _GEN_1297 : valid_240; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2323 = ~sc_fail_r ? _GEN_1298 : valid_241; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2324 = ~sc_fail_r ? _GEN_1299 : valid_242; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2325 = ~sc_fail_r ? _GEN_1300 : valid_243; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2326 = ~sc_fail_r ? _GEN_1301 : valid_244; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2327 = ~sc_fail_r ? _GEN_1302 : valid_245; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2328 = ~sc_fail_r ? _GEN_1303 : valid_246; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2329 = ~sc_fail_r ? _GEN_1304 : valid_247; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2330 = ~sc_fail_r ? _GEN_1305 : valid_248; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2331 = ~sc_fail_r ? _GEN_1306 : valid_249; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2332 = ~sc_fail_r ? _GEN_1307 : valid_250; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2333 = ~sc_fail_r ? _GEN_1308 : valid_251; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2334 = ~sc_fail_r ? _GEN_1309 : valid_252; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2335 = ~sc_fail_r ? _GEN_1310 : valid_253; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2336 = ~sc_fail_r ? _GEN_1311 : valid_254; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2337 = ~sc_fail_r ? _GEN_1312 : valid_255; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2338 = ~sc_fail_r ? _GEN_1313 : valid_256; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2339 = ~sc_fail_r ? _GEN_1314 : valid_257; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2340 = ~sc_fail_r ? _GEN_1315 : valid_258; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2341 = ~sc_fail_r ? _GEN_1316 : valid_259; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2342 = ~sc_fail_r ? _GEN_1317 : valid_260; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2343 = ~sc_fail_r ? _GEN_1318 : valid_261; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2344 = ~sc_fail_r ? _GEN_1319 : valid_262; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2345 = ~sc_fail_r ? _GEN_1320 : valid_263; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2346 = ~sc_fail_r ? _GEN_1321 : valid_264; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2347 = ~sc_fail_r ? _GEN_1322 : valid_265; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2348 = ~sc_fail_r ? _GEN_1323 : valid_266; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2349 = ~sc_fail_r ? _GEN_1324 : valid_267; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2350 = ~sc_fail_r ? _GEN_1325 : valid_268; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2351 = ~sc_fail_r ? _GEN_1326 : valid_269; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2352 = ~sc_fail_r ? _GEN_1327 : valid_270; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2353 = ~sc_fail_r ? _GEN_1328 : valid_271; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2354 = ~sc_fail_r ? _GEN_1329 : valid_272; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2355 = ~sc_fail_r ? _GEN_1330 : valid_273; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2356 = ~sc_fail_r ? _GEN_1331 : valid_274; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2357 = ~sc_fail_r ? _GEN_1332 : valid_275; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2358 = ~sc_fail_r ? _GEN_1333 : valid_276; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2359 = ~sc_fail_r ? _GEN_1334 : valid_277; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2360 = ~sc_fail_r ? _GEN_1335 : valid_278; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2361 = ~sc_fail_r ? _GEN_1336 : valid_279; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2362 = ~sc_fail_r ? _GEN_1337 : valid_280; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2363 = ~sc_fail_r ? _GEN_1338 : valid_281; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2364 = ~sc_fail_r ? _GEN_1339 : valid_282; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2365 = ~sc_fail_r ? _GEN_1340 : valid_283; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2366 = ~sc_fail_r ? _GEN_1341 : valid_284; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2367 = ~sc_fail_r ? _GEN_1342 : valid_285; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2368 = ~sc_fail_r ? _GEN_1343 : valid_286; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2369 = ~sc_fail_r ? _GEN_1344 : valid_287; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2370 = ~sc_fail_r ? _GEN_1345 : valid_288; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2371 = ~sc_fail_r ? _GEN_1346 : valid_289; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2372 = ~sc_fail_r ? _GEN_1347 : valid_290; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2373 = ~sc_fail_r ? _GEN_1348 : valid_291; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2374 = ~sc_fail_r ? _GEN_1349 : valid_292; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2375 = ~sc_fail_r ? _GEN_1350 : valid_293; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2376 = ~sc_fail_r ? _GEN_1351 : valid_294; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2377 = ~sc_fail_r ? _GEN_1352 : valid_295; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2378 = ~sc_fail_r ? _GEN_1353 : valid_296; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2379 = ~sc_fail_r ? _GEN_1354 : valid_297; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2380 = ~sc_fail_r ? _GEN_1355 : valid_298; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2381 = ~sc_fail_r ? _GEN_1356 : valid_299; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2382 = ~sc_fail_r ? _GEN_1357 : valid_300; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2383 = ~sc_fail_r ? _GEN_1358 : valid_301; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2384 = ~sc_fail_r ? _GEN_1359 : valid_302; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2385 = ~sc_fail_r ? _GEN_1360 : valid_303; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2386 = ~sc_fail_r ? _GEN_1361 : valid_304; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2387 = ~sc_fail_r ? _GEN_1362 : valid_305; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2388 = ~sc_fail_r ? _GEN_1363 : valid_306; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2389 = ~sc_fail_r ? _GEN_1364 : valid_307; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2390 = ~sc_fail_r ? _GEN_1365 : valid_308; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2391 = ~sc_fail_r ? _GEN_1366 : valid_309; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2392 = ~sc_fail_r ? _GEN_1367 : valid_310; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2393 = ~sc_fail_r ? _GEN_1368 : valid_311; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2394 = ~sc_fail_r ? _GEN_1369 : valid_312; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2395 = ~sc_fail_r ? _GEN_1370 : valid_313; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2396 = ~sc_fail_r ? _GEN_1371 : valid_314; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2397 = ~sc_fail_r ? _GEN_1372 : valid_315; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2398 = ~sc_fail_r ? _GEN_1373 : valid_316; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2399 = ~sc_fail_r ? _GEN_1374 : valid_317; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2400 = ~sc_fail_r ? _GEN_1375 : valid_318; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2401 = ~sc_fail_r ? _GEN_1376 : valid_319; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2402 = ~sc_fail_r ? _GEN_1377 : valid_320; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2403 = ~sc_fail_r ? _GEN_1378 : valid_321; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2404 = ~sc_fail_r ? _GEN_1379 : valid_322; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2405 = ~sc_fail_r ? _GEN_1380 : valid_323; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2406 = ~sc_fail_r ? _GEN_1381 : valid_324; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2407 = ~sc_fail_r ? _GEN_1382 : valid_325; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2408 = ~sc_fail_r ? _GEN_1383 : valid_326; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2409 = ~sc_fail_r ? _GEN_1384 : valid_327; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2410 = ~sc_fail_r ? _GEN_1385 : valid_328; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2411 = ~sc_fail_r ? _GEN_1386 : valid_329; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2412 = ~sc_fail_r ? _GEN_1387 : valid_330; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2413 = ~sc_fail_r ? _GEN_1388 : valid_331; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2414 = ~sc_fail_r ? _GEN_1389 : valid_332; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2415 = ~sc_fail_r ? _GEN_1390 : valid_333; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2416 = ~sc_fail_r ? _GEN_1391 : valid_334; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2417 = ~sc_fail_r ? _GEN_1392 : valid_335; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2418 = ~sc_fail_r ? _GEN_1393 : valid_336; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2419 = ~sc_fail_r ? _GEN_1394 : valid_337; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2420 = ~sc_fail_r ? _GEN_1395 : valid_338; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2421 = ~sc_fail_r ? _GEN_1396 : valid_339; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2422 = ~sc_fail_r ? _GEN_1397 : valid_340; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2423 = ~sc_fail_r ? _GEN_1398 : valid_341; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2424 = ~sc_fail_r ? _GEN_1399 : valid_342; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2425 = ~sc_fail_r ? _GEN_1400 : valid_343; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2426 = ~sc_fail_r ? _GEN_1401 : valid_344; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2427 = ~sc_fail_r ? _GEN_1402 : valid_345; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2428 = ~sc_fail_r ? _GEN_1403 : valid_346; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2429 = ~sc_fail_r ? _GEN_1404 : valid_347; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2430 = ~sc_fail_r ? _GEN_1405 : valid_348; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2431 = ~sc_fail_r ? _GEN_1406 : valid_349; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2432 = ~sc_fail_r ? _GEN_1407 : valid_350; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2433 = ~sc_fail_r ? _GEN_1408 : valid_351; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2434 = ~sc_fail_r ? _GEN_1409 : valid_352; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2435 = ~sc_fail_r ? _GEN_1410 : valid_353; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2436 = ~sc_fail_r ? _GEN_1411 : valid_354; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2437 = ~sc_fail_r ? _GEN_1412 : valid_355; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2438 = ~sc_fail_r ? _GEN_1413 : valid_356; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2439 = ~sc_fail_r ? _GEN_1414 : valid_357; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2440 = ~sc_fail_r ? _GEN_1415 : valid_358; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2441 = ~sc_fail_r ? _GEN_1416 : valid_359; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2442 = ~sc_fail_r ? _GEN_1417 : valid_360; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2443 = ~sc_fail_r ? _GEN_1418 : valid_361; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2444 = ~sc_fail_r ? _GEN_1419 : valid_362; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2445 = ~sc_fail_r ? _GEN_1420 : valid_363; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2446 = ~sc_fail_r ? _GEN_1421 : valid_364; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2447 = ~sc_fail_r ? _GEN_1422 : valid_365; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2448 = ~sc_fail_r ? _GEN_1423 : valid_366; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2449 = ~sc_fail_r ? _GEN_1424 : valid_367; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2450 = ~sc_fail_r ? _GEN_1425 : valid_368; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2451 = ~sc_fail_r ? _GEN_1426 : valid_369; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2452 = ~sc_fail_r ? _GEN_1427 : valid_370; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2453 = ~sc_fail_r ? _GEN_1428 : valid_371; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2454 = ~sc_fail_r ? _GEN_1429 : valid_372; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2455 = ~sc_fail_r ? _GEN_1430 : valid_373; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2456 = ~sc_fail_r ? _GEN_1431 : valid_374; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2457 = ~sc_fail_r ? _GEN_1432 : valid_375; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2458 = ~sc_fail_r ? _GEN_1433 : valid_376; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2459 = ~sc_fail_r ? _GEN_1434 : valid_377; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2460 = ~sc_fail_r ? _GEN_1435 : valid_378; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2461 = ~sc_fail_r ? _GEN_1436 : valid_379; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2462 = ~sc_fail_r ? _GEN_1437 : valid_380; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2463 = ~sc_fail_r ? _GEN_1438 : valid_381; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2464 = ~sc_fail_r ? _GEN_1439 : valid_382; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2465 = ~sc_fail_r ? _GEN_1440 : valid_383; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2466 = ~sc_fail_r ? _GEN_1441 : valid_384; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2467 = ~sc_fail_r ? _GEN_1442 : valid_385; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2468 = ~sc_fail_r ? _GEN_1443 : valid_386; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2469 = ~sc_fail_r ? _GEN_1444 : valid_387; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2470 = ~sc_fail_r ? _GEN_1445 : valid_388; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2471 = ~sc_fail_r ? _GEN_1446 : valid_389; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2472 = ~sc_fail_r ? _GEN_1447 : valid_390; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2473 = ~sc_fail_r ? _GEN_1448 : valid_391; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2474 = ~sc_fail_r ? _GEN_1449 : valid_392; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2475 = ~sc_fail_r ? _GEN_1450 : valid_393; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2476 = ~sc_fail_r ? _GEN_1451 : valid_394; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2477 = ~sc_fail_r ? _GEN_1452 : valid_395; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2478 = ~sc_fail_r ? _GEN_1453 : valid_396; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2479 = ~sc_fail_r ? _GEN_1454 : valid_397; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2480 = ~sc_fail_r ? _GEN_1455 : valid_398; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2481 = ~sc_fail_r ? _GEN_1456 : valid_399; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2482 = ~sc_fail_r ? _GEN_1457 : valid_400; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2483 = ~sc_fail_r ? _GEN_1458 : valid_401; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2484 = ~sc_fail_r ? _GEN_1459 : valid_402; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2485 = ~sc_fail_r ? _GEN_1460 : valid_403; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2486 = ~sc_fail_r ? _GEN_1461 : valid_404; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2487 = ~sc_fail_r ? _GEN_1462 : valid_405; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2488 = ~sc_fail_r ? _GEN_1463 : valid_406; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2489 = ~sc_fail_r ? _GEN_1464 : valid_407; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2490 = ~sc_fail_r ? _GEN_1465 : valid_408; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2491 = ~sc_fail_r ? _GEN_1466 : valid_409; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2492 = ~sc_fail_r ? _GEN_1467 : valid_410; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2493 = ~sc_fail_r ? _GEN_1468 : valid_411; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2494 = ~sc_fail_r ? _GEN_1469 : valid_412; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2495 = ~sc_fail_r ? _GEN_1470 : valid_413; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2496 = ~sc_fail_r ? _GEN_1471 : valid_414; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2497 = ~sc_fail_r ? _GEN_1472 : valid_415; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2498 = ~sc_fail_r ? _GEN_1473 : valid_416; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2499 = ~sc_fail_r ? _GEN_1474 : valid_417; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2500 = ~sc_fail_r ? _GEN_1475 : valid_418; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2501 = ~sc_fail_r ? _GEN_1476 : valid_419; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2502 = ~sc_fail_r ? _GEN_1477 : valid_420; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2503 = ~sc_fail_r ? _GEN_1478 : valid_421; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2504 = ~sc_fail_r ? _GEN_1479 : valid_422; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2505 = ~sc_fail_r ? _GEN_1480 : valid_423; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2506 = ~sc_fail_r ? _GEN_1481 : valid_424; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2507 = ~sc_fail_r ? _GEN_1482 : valid_425; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2508 = ~sc_fail_r ? _GEN_1483 : valid_426; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2509 = ~sc_fail_r ? _GEN_1484 : valid_427; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2510 = ~sc_fail_r ? _GEN_1485 : valid_428; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2511 = ~sc_fail_r ? _GEN_1486 : valid_429; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2512 = ~sc_fail_r ? _GEN_1487 : valid_430; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2513 = ~sc_fail_r ? _GEN_1488 : valid_431; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2514 = ~sc_fail_r ? _GEN_1489 : valid_432; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2515 = ~sc_fail_r ? _GEN_1490 : valid_433; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2516 = ~sc_fail_r ? _GEN_1491 : valid_434; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2517 = ~sc_fail_r ? _GEN_1492 : valid_435; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2518 = ~sc_fail_r ? _GEN_1493 : valid_436; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2519 = ~sc_fail_r ? _GEN_1494 : valid_437; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2520 = ~sc_fail_r ? _GEN_1495 : valid_438; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2521 = ~sc_fail_r ? _GEN_1496 : valid_439; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2522 = ~sc_fail_r ? _GEN_1497 : valid_440; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2523 = ~sc_fail_r ? _GEN_1498 : valid_441; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2524 = ~sc_fail_r ? _GEN_1499 : valid_442; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2525 = ~sc_fail_r ? _GEN_1500 : valid_443; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2526 = ~sc_fail_r ? _GEN_1501 : valid_444; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2527 = ~sc_fail_r ? _GEN_1502 : valid_445; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2528 = ~sc_fail_r ? _GEN_1503 : valid_446; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2529 = ~sc_fail_r ? _GEN_1504 : valid_447; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2530 = ~sc_fail_r ? _GEN_1505 : valid_448; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2531 = ~sc_fail_r ? _GEN_1506 : valid_449; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2532 = ~sc_fail_r ? _GEN_1507 : valid_450; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2533 = ~sc_fail_r ? _GEN_1508 : valid_451; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2534 = ~sc_fail_r ? _GEN_1509 : valid_452; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2535 = ~sc_fail_r ? _GEN_1510 : valid_453; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2536 = ~sc_fail_r ? _GEN_1511 : valid_454; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2537 = ~sc_fail_r ? _GEN_1512 : valid_455; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2538 = ~sc_fail_r ? _GEN_1513 : valid_456; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2539 = ~sc_fail_r ? _GEN_1514 : valid_457; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2540 = ~sc_fail_r ? _GEN_1515 : valid_458; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2541 = ~sc_fail_r ? _GEN_1516 : valid_459; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2542 = ~sc_fail_r ? _GEN_1517 : valid_460; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2543 = ~sc_fail_r ? _GEN_1518 : valid_461; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2544 = ~sc_fail_r ? _GEN_1519 : valid_462; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2545 = ~sc_fail_r ? _GEN_1520 : valid_463; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2546 = ~sc_fail_r ? _GEN_1521 : valid_464; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2547 = ~sc_fail_r ? _GEN_1522 : valid_465; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2548 = ~sc_fail_r ? _GEN_1523 : valid_466; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2549 = ~sc_fail_r ? _GEN_1524 : valid_467; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2550 = ~sc_fail_r ? _GEN_1525 : valid_468; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2551 = ~sc_fail_r ? _GEN_1526 : valid_469; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2552 = ~sc_fail_r ? _GEN_1527 : valid_470; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2553 = ~sc_fail_r ? _GEN_1528 : valid_471; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2554 = ~sc_fail_r ? _GEN_1529 : valid_472; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2555 = ~sc_fail_r ? _GEN_1530 : valid_473; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2556 = ~sc_fail_r ? _GEN_1531 : valid_474; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2557 = ~sc_fail_r ? _GEN_1532 : valid_475; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2558 = ~sc_fail_r ? _GEN_1533 : valid_476; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2559 = ~sc_fail_r ? _GEN_1534 : valid_477; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2560 = ~sc_fail_r ? _GEN_1535 : valid_478; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2561 = ~sc_fail_r ? _GEN_1536 : valid_479; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2562 = ~sc_fail_r ? _GEN_1537 : valid_480; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2563 = ~sc_fail_r ? _GEN_1538 : valid_481; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2564 = ~sc_fail_r ? _GEN_1539 : valid_482; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2565 = ~sc_fail_r ? _GEN_1540 : valid_483; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2566 = ~sc_fail_r ? _GEN_1541 : valid_484; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2567 = ~sc_fail_r ? _GEN_1542 : valid_485; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2568 = ~sc_fail_r ? _GEN_1543 : valid_486; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2569 = ~sc_fail_r ? _GEN_1544 : valid_487; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2570 = ~sc_fail_r ? _GEN_1545 : valid_488; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2571 = ~sc_fail_r ? _GEN_1546 : valid_489; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2572 = ~sc_fail_r ? _GEN_1547 : valid_490; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2573 = ~sc_fail_r ? _GEN_1548 : valid_491; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2574 = ~sc_fail_r ? _GEN_1549 : valid_492; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2575 = ~sc_fail_r ? _GEN_1550 : valid_493; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2576 = ~sc_fail_r ? _GEN_1551 : valid_494; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2577 = ~sc_fail_r ? _GEN_1552 : valid_495; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2578 = ~sc_fail_r ? _GEN_1553 : valid_496; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2579 = ~sc_fail_r ? _GEN_1554 : valid_497; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2580 = ~sc_fail_r ? _GEN_1555 : valid_498; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2581 = ~sc_fail_r ? _GEN_1556 : valid_499; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2582 = ~sc_fail_r ? _GEN_1557 : valid_500; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2583 = ~sc_fail_r ? _GEN_1558 : valid_501; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2584 = ~sc_fail_r ? _GEN_1559 : valid_502; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2585 = ~sc_fail_r ? _GEN_1560 : valid_503; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2586 = ~sc_fail_r ? _GEN_1561 : valid_504; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2587 = ~sc_fail_r ? _GEN_1562 : valid_505; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2588 = ~sc_fail_r ? _GEN_1563 : valid_506; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2589 = ~sc_fail_r ? _GEN_1564 : valid_507; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2590 = ~sc_fail_r ? _GEN_1565 : valid_508; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2591 = ~sc_fail_r ? _GEN_1566 : valid_509; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2592 = ~sc_fail_r ? _GEN_1567 : valid_510; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2593 = ~sc_fail_r ? _GEN_1568 : valid_511; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2594 = ~sc_fail_r ? _GEN_1569 : valid_512; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2595 = ~sc_fail_r ? _GEN_1570 : valid_513; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2596 = ~sc_fail_r ? _GEN_1571 : valid_514; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2597 = ~sc_fail_r ? _GEN_1572 : valid_515; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2598 = ~sc_fail_r ? _GEN_1573 : valid_516; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2599 = ~sc_fail_r ? _GEN_1574 : valid_517; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2600 = ~sc_fail_r ? _GEN_1575 : valid_518; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2601 = ~sc_fail_r ? _GEN_1576 : valid_519; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2602 = ~sc_fail_r ? _GEN_1577 : valid_520; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2603 = ~sc_fail_r ? _GEN_1578 : valid_521; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2604 = ~sc_fail_r ? _GEN_1579 : valid_522; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2605 = ~sc_fail_r ? _GEN_1580 : valid_523; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2606 = ~sc_fail_r ? _GEN_1581 : valid_524; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2607 = ~sc_fail_r ? _GEN_1582 : valid_525; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2608 = ~sc_fail_r ? _GEN_1583 : valid_526; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2609 = ~sc_fail_r ? _GEN_1584 : valid_527; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2610 = ~sc_fail_r ? _GEN_1585 : valid_528; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2611 = ~sc_fail_r ? _GEN_1586 : valid_529; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2612 = ~sc_fail_r ? _GEN_1587 : valid_530; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2613 = ~sc_fail_r ? _GEN_1588 : valid_531; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2614 = ~sc_fail_r ? _GEN_1589 : valid_532; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2615 = ~sc_fail_r ? _GEN_1590 : valid_533; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2616 = ~sc_fail_r ? _GEN_1591 : valid_534; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2617 = ~sc_fail_r ? _GEN_1592 : valid_535; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2618 = ~sc_fail_r ? _GEN_1593 : valid_536; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2619 = ~sc_fail_r ? _GEN_1594 : valid_537; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2620 = ~sc_fail_r ? _GEN_1595 : valid_538; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2621 = ~sc_fail_r ? _GEN_1596 : valid_539; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2622 = ~sc_fail_r ? _GEN_1597 : valid_540; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2623 = ~sc_fail_r ? _GEN_1598 : valid_541; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2624 = ~sc_fail_r ? _GEN_1599 : valid_542; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2625 = ~sc_fail_r ? _GEN_1600 : valid_543; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2626 = ~sc_fail_r ? _GEN_1601 : valid_544; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2627 = ~sc_fail_r ? _GEN_1602 : valid_545; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2628 = ~sc_fail_r ? _GEN_1603 : valid_546; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2629 = ~sc_fail_r ? _GEN_1604 : valid_547; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2630 = ~sc_fail_r ? _GEN_1605 : valid_548; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2631 = ~sc_fail_r ? _GEN_1606 : valid_549; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2632 = ~sc_fail_r ? _GEN_1607 : valid_550; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2633 = ~sc_fail_r ? _GEN_1608 : valid_551; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2634 = ~sc_fail_r ? _GEN_1609 : valid_552; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2635 = ~sc_fail_r ? _GEN_1610 : valid_553; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2636 = ~sc_fail_r ? _GEN_1611 : valid_554; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2637 = ~sc_fail_r ? _GEN_1612 : valid_555; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2638 = ~sc_fail_r ? _GEN_1613 : valid_556; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2639 = ~sc_fail_r ? _GEN_1614 : valid_557; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2640 = ~sc_fail_r ? _GEN_1615 : valid_558; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2641 = ~sc_fail_r ? _GEN_1616 : valid_559; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2642 = ~sc_fail_r ? _GEN_1617 : valid_560; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2643 = ~sc_fail_r ? _GEN_1618 : valid_561; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2644 = ~sc_fail_r ? _GEN_1619 : valid_562; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2645 = ~sc_fail_r ? _GEN_1620 : valid_563; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2646 = ~sc_fail_r ? _GEN_1621 : valid_564; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2647 = ~sc_fail_r ? _GEN_1622 : valid_565; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2648 = ~sc_fail_r ? _GEN_1623 : valid_566; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2649 = ~sc_fail_r ? _GEN_1624 : valid_567; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2650 = ~sc_fail_r ? _GEN_1625 : valid_568; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2651 = ~sc_fail_r ? _GEN_1626 : valid_569; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2652 = ~sc_fail_r ? _GEN_1627 : valid_570; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2653 = ~sc_fail_r ? _GEN_1628 : valid_571; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2654 = ~sc_fail_r ? _GEN_1629 : valid_572; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2655 = ~sc_fail_r ? _GEN_1630 : valid_573; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2656 = ~sc_fail_r ? _GEN_1631 : valid_574; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2657 = ~sc_fail_r ? _GEN_1632 : valid_575; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2658 = ~sc_fail_r ? _GEN_1633 : valid_576; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2659 = ~sc_fail_r ? _GEN_1634 : valid_577; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2660 = ~sc_fail_r ? _GEN_1635 : valid_578; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2661 = ~sc_fail_r ? _GEN_1636 : valid_579; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2662 = ~sc_fail_r ? _GEN_1637 : valid_580; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2663 = ~sc_fail_r ? _GEN_1638 : valid_581; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2664 = ~sc_fail_r ? _GEN_1639 : valid_582; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2665 = ~sc_fail_r ? _GEN_1640 : valid_583; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2666 = ~sc_fail_r ? _GEN_1641 : valid_584; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2667 = ~sc_fail_r ? _GEN_1642 : valid_585; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2668 = ~sc_fail_r ? _GEN_1643 : valid_586; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2669 = ~sc_fail_r ? _GEN_1644 : valid_587; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2670 = ~sc_fail_r ? _GEN_1645 : valid_588; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2671 = ~sc_fail_r ? _GEN_1646 : valid_589; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2672 = ~sc_fail_r ? _GEN_1647 : valid_590; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2673 = ~sc_fail_r ? _GEN_1648 : valid_591; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2674 = ~sc_fail_r ? _GEN_1649 : valid_592; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2675 = ~sc_fail_r ? _GEN_1650 : valid_593; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2676 = ~sc_fail_r ? _GEN_1651 : valid_594; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2677 = ~sc_fail_r ? _GEN_1652 : valid_595; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2678 = ~sc_fail_r ? _GEN_1653 : valid_596; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2679 = ~sc_fail_r ? _GEN_1654 : valid_597; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2680 = ~sc_fail_r ? _GEN_1655 : valid_598; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2681 = ~sc_fail_r ? _GEN_1656 : valid_599; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2682 = ~sc_fail_r ? _GEN_1657 : valid_600; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2683 = ~sc_fail_r ? _GEN_1658 : valid_601; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2684 = ~sc_fail_r ? _GEN_1659 : valid_602; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2685 = ~sc_fail_r ? _GEN_1660 : valid_603; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2686 = ~sc_fail_r ? _GEN_1661 : valid_604; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2687 = ~sc_fail_r ? _GEN_1662 : valid_605; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2688 = ~sc_fail_r ? _GEN_1663 : valid_606; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2689 = ~sc_fail_r ? _GEN_1664 : valid_607; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2690 = ~sc_fail_r ? _GEN_1665 : valid_608; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2691 = ~sc_fail_r ? _GEN_1666 : valid_609; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2692 = ~sc_fail_r ? _GEN_1667 : valid_610; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2693 = ~sc_fail_r ? _GEN_1668 : valid_611; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2694 = ~sc_fail_r ? _GEN_1669 : valid_612; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2695 = ~sc_fail_r ? _GEN_1670 : valid_613; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2696 = ~sc_fail_r ? _GEN_1671 : valid_614; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2697 = ~sc_fail_r ? _GEN_1672 : valid_615; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2698 = ~sc_fail_r ? _GEN_1673 : valid_616; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2699 = ~sc_fail_r ? _GEN_1674 : valid_617; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2700 = ~sc_fail_r ? _GEN_1675 : valid_618; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2701 = ~sc_fail_r ? _GEN_1676 : valid_619; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2702 = ~sc_fail_r ? _GEN_1677 : valid_620; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2703 = ~sc_fail_r ? _GEN_1678 : valid_621; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2704 = ~sc_fail_r ? _GEN_1679 : valid_622; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2705 = ~sc_fail_r ? _GEN_1680 : valid_623; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2706 = ~sc_fail_r ? _GEN_1681 : valid_624; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2707 = ~sc_fail_r ? _GEN_1682 : valid_625; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2708 = ~sc_fail_r ? _GEN_1683 : valid_626; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2709 = ~sc_fail_r ? _GEN_1684 : valid_627; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2710 = ~sc_fail_r ? _GEN_1685 : valid_628; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2711 = ~sc_fail_r ? _GEN_1686 : valid_629; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2712 = ~sc_fail_r ? _GEN_1687 : valid_630; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2713 = ~sc_fail_r ? _GEN_1688 : valid_631; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2714 = ~sc_fail_r ? _GEN_1689 : valid_632; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2715 = ~sc_fail_r ? _GEN_1690 : valid_633; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2716 = ~sc_fail_r ? _GEN_1691 : valid_634; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2717 = ~sc_fail_r ? _GEN_1692 : valid_635; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2718 = ~sc_fail_r ? _GEN_1693 : valid_636; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2719 = ~sc_fail_r ? _GEN_1694 : valid_637; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2720 = ~sc_fail_r ? _GEN_1695 : valid_638; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2721 = ~sc_fail_r ? _GEN_1696 : valid_639; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2722 = ~sc_fail_r ? _GEN_1697 : valid_640; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2723 = ~sc_fail_r ? _GEN_1698 : valid_641; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2724 = ~sc_fail_r ? _GEN_1699 : valid_642; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2725 = ~sc_fail_r ? _GEN_1700 : valid_643; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2726 = ~sc_fail_r ? _GEN_1701 : valid_644; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2727 = ~sc_fail_r ? _GEN_1702 : valid_645; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2728 = ~sc_fail_r ? _GEN_1703 : valid_646; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2729 = ~sc_fail_r ? _GEN_1704 : valid_647; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2730 = ~sc_fail_r ? _GEN_1705 : valid_648; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2731 = ~sc_fail_r ? _GEN_1706 : valid_649; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2732 = ~sc_fail_r ? _GEN_1707 : valid_650; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2733 = ~sc_fail_r ? _GEN_1708 : valid_651; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2734 = ~sc_fail_r ? _GEN_1709 : valid_652; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2735 = ~sc_fail_r ? _GEN_1710 : valid_653; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2736 = ~sc_fail_r ? _GEN_1711 : valid_654; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2737 = ~sc_fail_r ? _GEN_1712 : valid_655; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2738 = ~sc_fail_r ? _GEN_1713 : valid_656; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2739 = ~sc_fail_r ? _GEN_1714 : valid_657; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2740 = ~sc_fail_r ? _GEN_1715 : valid_658; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2741 = ~sc_fail_r ? _GEN_1716 : valid_659; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2742 = ~sc_fail_r ? _GEN_1717 : valid_660; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2743 = ~sc_fail_r ? _GEN_1718 : valid_661; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2744 = ~sc_fail_r ? _GEN_1719 : valid_662; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2745 = ~sc_fail_r ? _GEN_1720 : valid_663; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2746 = ~sc_fail_r ? _GEN_1721 : valid_664; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2747 = ~sc_fail_r ? _GEN_1722 : valid_665; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2748 = ~sc_fail_r ? _GEN_1723 : valid_666; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2749 = ~sc_fail_r ? _GEN_1724 : valid_667; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2750 = ~sc_fail_r ? _GEN_1725 : valid_668; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2751 = ~sc_fail_r ? _GEN_1726 : valid_669; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2752 = ~sc_fail_r ? _GEN_1727 : valid_670; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2753 = ~sc_fail_r ? _GEN_1728 : valid_671; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2754 = ~sc_fail_r ? _GEN_1729 : valid_672; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2755 = ~sc_fail_r ? _GEN_1730 : valid_673; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2756 = ~sc_fail_r ? _GEN_1731 : valid_674; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2757 = ~sc_fail_r ? _GEN_1732 : valid_675; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2758 = ~sc_fail_r ? _GEN_1733 : valid_676; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2759 = ~sc_fail_r ? _GEN_1734 : valid_677; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2760 = ~sc_fail_r ? _GEN_1735 : valid_678; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2761 = ~sc_fail_r ? _GEN_1736 : valid_679; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2762 = ~sc_fail_r ? _GEN_1737 : valid_680; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2763 = ~sc_fail_r ? _GEN_1738 : valid_681; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2764 = ~sc_fail_r ? _GEN_1739 : valid_682; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2765 = ~sc_fail_r ? _GEN_1740 : valid_683; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2766 = ~sc_fail_r ? _GEN_1741 : valid_684; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2767 = ~sc_fail_r ? _GEN_1742 : valid_685; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2768 = ~sc_fail_r ? _GEN_1743 : valid_686; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2769 = ~sc_fail_r ? _GEN_1744 : valid_687; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2770 = ~sc_fail_r ? _GEN_1745 : valid_688; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2771 = ~sc_fail_r ? _GEN_1746 : valid_689; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2772 = ~sc_fail_r ? _GEN_1747 : valid_690; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2773 = ~sc_fail_r ? _GEN_1748 : valid_691; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2774 = ~sc_fail_r ? _GEN_1749 : valid_692; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2775 = ~sc_fail_r ? _GEN_1750 : valid_693; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2776 = ~sc_fail_r ? _GEN_1751 : valid_694; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2777 = ~sc_fail_r ? _GEN_1752 : valid_695; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2778 = ~sc_fail_r ? _GEN_1753 : valid_696; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2779 = ~sc_fail_r ? _GEN_1754 : valid_697; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2780 = ~sc_fail_r ? _GEN_1755 : valid_698; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2781 = ~sc_fail_r ? _GEN_1756 : valid_699; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2782 = ~sc_fail_r ? _GEN_1757 : valid_700; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2783 = ~sc_fail_r ? _GEN_1758 : valid_701; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2784 = ~sc_fail_r ? _GEN_1759 : valid_702; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2785 = ~sc_fail_r ? _GEN_1760 : valid_703; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2786 = ~sc_fail_r ? _GEN_1761 : valid_704; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2787 = ~sc_fail_r ? _GEN_1762 : valid_705; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2788 = ~sc_fail_r ? _GEN_1763 : valid_706; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2789 = ~sc_fail_r ? _GEN_1764 : valid_707; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2790 = ~sc_fail_r ? _GEN_1765 : valid_708; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2791 = ~sc_fail_r ? _GEN_1766 : valid_709; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2792 = ~sc_fail_r ? _GEN_1767 : valid_710; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2793 = ~sc_fail_r ? _GEN_1768 : valid_711; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2794 = ~sc_fail_r ? _GEN_1769 : valid_712; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2795 = ~sc_fail_r ? _GEN_1770 : valid_713; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2796 = ~sc_fail_r ? _GEN_1771 : valid_714; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2797 = ~sc_fail_r ? _GEN_1772 : valid_715; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2798 = ~sc_fail_r ? _GEN_1773 : valid_716; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2799 = ~sc_fail_r ? _GEN_1774 : valid_717; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2800 = ~sc_fail_r ? _GEN_1775 : valid_718; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2801 = ~sc_fail_r ? _GEN_1776 : valid_719; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2802 = ~sc_fail_r ? _GEN_1777 : valid_720; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2803 = ~sc_fail_r ? _GEN_1778 : valid_721; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2804 = ~sc_fail_r ? _GEN_1779 : valid_722; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2805 = ~sc_fail_r ? _GEN_1780 : valid_723; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2806 = ~sc_fail_r ? _GEN_1781 : valid_724; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2807 = ~sc_fail_r ? _GEN_1782 : valid_725; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2808 = ~sc_fail_r ? _GEN_1783 : valid_726; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2809 = ~sc_fail_r ? _GEN_1784 : valid_727; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2810 = ~sc_fail_r ? _GEN_1785 : valid_728; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2811 = ~sc_fail_r ? _GEN_1786 : valid_729; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2812 = ~sc_fail_r ? _GEN_1787 : valid_730; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2813 = ~sc_fail_r ? _GEN_1788 : valid_731; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2814 = ~sc_fail_r ? _GEN_1789 : valid_732; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2815 = ~sc_fail_r ? _GEN_1790 : valid_733; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2816 = ~sc_fail_r ? _GEN_1791 : valid_734; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2817 = ~sc_fail_r ? _GEN_1792 : valid_735; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2818 = ~sc_fail_r ? _GEN_1793 : valid_736; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2819 = ~sc_fail_r ? _GEN_1794 : valid_737; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2820 = ~sc_fail_r ? _GEN_1795 : valid_738; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2821 = ~sc_fail_r ? _GEN_1796 : valid_739; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2822 = ~sc_fail_r ? _GEN_1797 : valid_740; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2823 = ~sc_fail_r ? _GEN_1798 : valid_741; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2824 = ~sc_fail_r ? _GEN_1799 : valid_742; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2825 = ~sc_fail_r ? _GEN_1800 : valid_743; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2826 = ~sc_fail_r ? _GEN_1801 : valid_744; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2827 = ~sc_fail_r ? _GEN_1802 : valid_745; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2828 = ~sc_fail_r ? _GEN_1803 : valid_746; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2829 = ~sc_fail_r ? _GEN_1804 : valid_747; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2830 = ~sc_fail_r ? _GEN_1805 : valid_748; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2831 = ~sc_fail_r ? _GEN_1806 : valid_749; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2832 = ~sc_fail_r ? _GEN_1807 : valid_750; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2833 = ~sc_fail_r ? _GEN_1808 : valid_751; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2834 = ~sc_fail_r ? _GEN_1809 : valid_752; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2835 = ~sc_fail_r ? _GEN_1810 : valid_753; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2836 = ~sc_fail_r ? _GEN_1811 : valid_754; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2837 = ~sc_fail_r ? _GEN_1812 : valid_755; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2838 = ~sc_fail_r ? _GEN_1813 : valid_756; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2839 = ~sc_fail_r ? _GEN_1814 : valid_757; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2840 = ~sc_fail_r ? _GEN_1815 : valid_758; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2841 = ~sc_fail_r ? _GEN_1816 : valid_759; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2842 = ~sc_fail_r ? _GEN_1817 : valid_760; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2843 = ~sc_fail_r ? _GEN_1818 : valid_761; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2844 = ~sc_fail_r ? _GEN_1819 : valid_762; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2845 = ~sc_fail_r ? _GEN_1820 : valid_763; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2846 = ~sc_fail_r ? _GEN_1821 : valid_764; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2847 = ~sc_fail_r ? _GEN_1822 : valid_765; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2848 = ~sc_fail_r ? _GEN_1823 : valid_766; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2849 = ~sc_fail_r ? _GEN_1824 : valid_767; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2850 = ~sc_fail_r ? _GEN_1825 : valid_768; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2851 = ~sc_fail_r ? _GEN_1826 : valid_769; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2852 = ~sc_fail_r ? _GEN_1827 : valid_770; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2853 = ~sc_fail_r ? _GEN_1828 : valid_771; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2854 = ~sc_fail_r ? _GEN_1829 : valid_772; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2855 = ~sc_fail_r ? _GEN_1830 : valid_773; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2856 = ~sc_fail_r ? _GEN_1831 : valid_774; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2857 = ~sc_fail_r ? _GEN_1832 : valid_775; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2858 = ~sc_fail_r ? _GEN_1833 : valid_776; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2859 = ~sc_fail_r ? _GEN_1834 : valid_777; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2860 = ~sc_fail_r ? _GEN_1835 : valid_778; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2861 = ~sc_fail_r ? _GEN_1836 : valid_779; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2862 = ~sc_fail_r ? _GEN_1837 : valid_780; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2863 = ~sc_fail_r ? _GEN_1838 : valid_781; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2864 = ~sc_fail_r ? _GEN_1839 : valid_782; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2865 = ~sc_fail_r ? _GEN_1840 : valid_783; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2866 = ~sc_fail_r ? _GEN_1841 : valid_784; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2867 = ~sc_fail_r ? _GEN_1842 : valid_785; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2868 = ~sc_fail_r ? _GEN_1843 : valid_786; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2869 = ~sc_fail_r ? _GEN_1844 : valid_787; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2870 = ~sc_fail_r ? _GEN_1845 : valid_788; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2871 = ~sc_fail_r ? _GEN_1846 : valid_789; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2872 = ~sc_fail_r ? _GEN_1847 : valid_790; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2873 = ~sc_fail_r ? _GEN_1848 : valid_791; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2874 = ~sc_fail_r ? _GEN_1849 : valid_792; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2875 = ~sc_fail_r ? _GEN_1850 : valid_793; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2876 = ~sc_fail_r ? _GEN_1851 : valid_794; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2877 = ~sc_fail_r ? _GEN_1852 : valid_795; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2878 = ~sc_fail_r ? _GEN_1853 : valid_796; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2879 = ~sc_fail_r ? _GEN_1854 : valid_797; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2880 = ~sc_fail_r ? _GEN_1855 : valid_798; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2881 = ~sc_fail_r ? _GEN_1856 : valid_799; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2882 = ~sc_fail_r ? _GEN_1857 : valid_800; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2883 = ~sc_fail_r ? _GEN_1858 : valid_801; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2884 = ~sc_fail_r ? _GEN_1859 : valid_802; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2885 = ~sc_fail_r ? _GEN_1860 : valid_803; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2886 = ~sc_fail_r ? _GEN_1861 : valid_804; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2887 = ~sc_fail_r ? _GEN_1862 : valid_805; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2888 = ~sc_fail_r ? _GEN_1863 : valid_806; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2889 = ~sc_fail_r ? _GEN_1864 : valid_807; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2890 = ~sc_fail_r ? _GEN_1865 : valid_808; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2891 = ~sc_fail_r ? _GEN_1866 : valid_809; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2892 = ~sc_fail_r ? _GEN_1867 : valid_810; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2893 = ~sc_fail_r ? _GEN_1868 : valid_811; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2894 = ~sc_fail_r ? _GEN_1869 : valid_812; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2895 = ~sc_fail_r ? _GEN_1870 : valid_813; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2896 = ~sc_fail_r ? _GEN_1871 : valid_814; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2897 = ~sc_fail_r ? _GEN_1872 : valid_815; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2898 = ~sc_fail_r ? _GEN_1873 : valid_816; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2899 = ~sc_fail_r ? _GEN_1874 : valid_817; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2900 = ~sc_fail_r ? _GEN_1875 : valid_818; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2901 = ~sc_fail_r ? _GEN_1876 : valid_819; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2902 = ~sc_fail_r ? _GEN_1877 : valid_820; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2903 = ~sc_fail_r ? _GEN_1878 : valid_821; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2904 = ~sc_fail_r ? _GEN_1879 : valid_822; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2905 = ~sc_fail_r ? _GEN_1880 : valid_823; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2906 = ~sc_fail_r ? _GEN_1881 : valid_824; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2907 = ~sc_fail_r ? _GEN_1882 : valid_825; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2908 = ~sc_fail_r ? _GEN_1883 : valid_826; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2909 = ~sc_fail_r ? _GEN_1884 : valid_827; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2910 = ~sc_fail_r ? _GEN_1885 : valid_828; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2911 = ~sc_fail_r ? _GEN_1886 : valid_829; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2912 = ~sc_fail_r ? _GEN_1887 : valid_830; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2913 = ~sc_fail_r ? _GEN_1888 : valid_831; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2914 = ~sc_fail_r ? _GEN_1889 : valid_832; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2915 = ~sc_fail_r ? _GEN_1890 : valid_833; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2916 = ~sc_fail_r ? _GEN_1891 : valid_834; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2917 = ~sc_fail_r ? _GEN_1892 : valid_835; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2918 = ~sc_fail_r ? _GEN_1893 : valid_836; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2919 = ~sc_fail_r ? _GEN_1894 : valid_837; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2920 = ~sc_fail_r ? _GEN_1895 : valid_838; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2921 = ~sc_fail_r ? _GEN_1896 : valid_839; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2922 = ~sc_fail_r ? _GEN_1897 : valid_840; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2923 = ~sc_fail_r ? _GEN_1898 : valid_841; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2924 = ~sc_fail_r ? _GEN_1899 : valid_842; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2925 = ~sc_fail_r ? _GEN_1900 : valid_843; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2926 = ~sc_fail_r ? _GEN_1901 : valid_844; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2927 = ~sc_fail_r ? _GEN_1902 : valid_845; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2928 = ~sc_fail_r ? _GEN_1903 : valid_846; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2929 = ~sc_fail_r ? _GEN_1904 : valid_847; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2930 = ~sc_fail_r ? _GEN_1905 : valid_848; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2931 = ~sc_fail_r ? _GEN_1906 : valid_849; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2932 = ~sc_fail_r ? _GEN_1907 : valid_850; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2933 = ~sc_fail_r ? _GEN_1908 : valid_851; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2934 = ~sc_fail_r ? _GEN_1909 : valid_852; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2935 = ~sc_fail_r ? _GEN_1910 : valid_853; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2936 = ~sc_fail_r ? _GEN_1911 : valid_854; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2937 = ~sc_fail_r ? _GEN_1912 : valid_855; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2938 = ~sc_fail_r ? _GEN_1913 : valid_856; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2939 = ~sc_fail_r ? _GEN_1914 : valid_857; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2940 = ~sc_fail_r ? _GEN_1915 : valid_858; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2941 = ~sc_fail_r ? _GEN_1916 : valid_859; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2942 = ~sc_fail_r ? _GEN_1917 : valid_860; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2943 = ~sc_fail_r ? _GEN_1918 : valid_861; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2944 = ~sc_fail_r ? _GEN_1919 : valid_862; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2945 = ~sc_fail_r ? _GEN_1920 : valid_863; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2946 = ~sc_fail_r ? _GEN_1921 : valid_864; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2947 = ~sc_fail_r ? _GEN_1922 : valid_865; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2948 = ~sc_fail_r ? _GEN_1923 : valid_866; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2949 = ~sc_fail_r ? _GEN_1924 : valid_867; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2950 = ~sc_fail_r ? _GEN_1925 : valid_868; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2951 = ~sc_fail_r ? _GEN_1926 : valid_869; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2952 = ~sc_fail_r ? _GEN_1927 : valid_870; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2953 = ~sc_fail_r ? _GEN_1928 : valid_871; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2954 = ~sc_fail_r ? _GEN_1929 : valid_872; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2955 = ~sc_fail_r ? _GEN_1930 : valid_873; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2956 = ~sc_fail_r ? _GEN_1931 : valid_874; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2957 = ~sc_fail_r ? _GEN_1932 : valid_875; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2958 = ~sc_fail_r ? _GEN_1933 : valid_876; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2959 = ~sc_fail_r ? _GEN_1934 : valid_877; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2960 = ~sc_fail_r ? _GEN_1935 : valid_878; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2961 = ~sc_fail_r ? _GEN_1936 : valid_879; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2962 = ~sc_fail_r ? _GEN_1937 : valid_880; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2963 = ~sc_fail_r ? _GEN_1938 : valid_881; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2964 = ~sc_fail_r ? _GEN_1939 : valid_882; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2965 = ~sc_fail_r ? _GEN_1940 : valid_883; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2966 = ~sc_fail_r ? _GEN_1941 : valid_884; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2967 = ~sc_fail_r ? _GEN_1942 : valid_885; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2968 = ~sc_fail_r ? _GEN_1943 : valid_886; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2969 = ~sc_fail_r ? _GEN_1944 : valid_887; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2970 = ~sc_fail_r ? _GEN_1945 : valid_888; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2971 = ~sc_fail_r ? _GEN_1946 : valid_889; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2972 = ~sc_fail_r ? _GEN_1947 : valid_890; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2973 = ~sc_fail_r ? _GEN_1948 : valid_891; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2974 = ~sc_fail_r ? _GEN_1949 : valid_892; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2975 = ~sc_fail_r ? _GEN_1950 : valid_893; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2976 = ~sc_fail_r ? _GEN_1951 : valid_894; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2977 = ~sc_fail_r ? _GEN_1952 : valid_895; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2978 = ~sc_fail_r ? _GEN_1953 : valid_896; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2979 = ~sc_fail_r ? _GEN_1954 : valid_897; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2980 = ~sc_fail_r ? _GEN_1955 : valid_898; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2981 = ~sc_fail_r ? _GEN_1956 : valid_899; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2982 = ~sc_fail_r ? _GEN_1957 : valid_900; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2983 = ~sc_fail_r ? _GEN_1958 : valid_901; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2984 = ~sc_fail_r ? _GEN_1959 : valid_902; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2985 = ~sc_fail_r ? _GEN_1960 : valid_903; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2986 = ~sc_fail_r ? _GEN_1961 : valid_904; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2987 = ~sc_fail_r ? _GEN_1962 : valid_905; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2988 = ~sc_fail_r ? _GEN_1963 : valid_906; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2989 = ~sc_fail_r ? _GEN_1964 : valid_907; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2990 = ~sc_fail_r ? _GEN_1965 : valid_908; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2991 = ~sc_fail_r ? _GEN_1966 : valid_909; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2992 = ~sc_fail_r ? _GEN_1967 : valid_910; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2993 = ~sc_fail_r ? _GEN_1968 : valid_911; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2994 = ~sc_fail_r ? _GEN_1969 : valid_912; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2995 = ~sc_fail_r ? _GEN_1970 : valid_913; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2996 = ~sc_fail_r ? _GEN_1971 : valid_914; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2997 = ~sc_fail_r ? _GEN_1972 : valid_915; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2998 = ~sc_fail_r ? _GEN_1973 : valid_916; // @[DCache.scala 171:24 56:22]
  wire  _GEN_2999 = ~sc_fail_r ? _GEN_1974 : valid_917; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3000 = ~sc_fail_r ? _GEN_1975 : valid_918; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3001 = ~sc_fail_r ? _GEN_1976 : valid_919; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3002 = ~sc_fail_r ? _GEN_1977 : valid_920; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3003 = ~sc_fail_r ? _GEN_1978 : valid_921; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3004 = ~sc_fail_r ? _GEN_1979 : valid_922; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3005 = ~sc_fail_r ? _GEN_1980 : valid_923; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3006 = ~sc_fail_r ? _GEN_1981 : valid_924; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3007 = ~sc_fail_r ? _GEN_1982 : valid_925; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3008 = ~sc_fail_r ? _GEN_1983 : valid_926; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3009 = ~sc_fail_r ? _GEN_1984 : valid_927; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3010 = ~sc_fail_r ? _GEN_1985 : valid_928; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3011 = ~sc_fail_r ? _GEN_1986 : valid_929; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3012 = ~sc_fail_r ? _GEN_1987 : valid_930; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3013 = ~sc_fail_r ? _GEN_1988 : valid_931; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3014 = ~sc_fail_r ? _GEN_1989 : valid_932; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3015 = ~sc_fail_r ? _GEN_1990 : valid_933; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3016 = ~sc_fail_r ? _GEN_1991 : valid_934; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3017 = ~sc_fail_r ? _GEN_1992 : valid_935; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3018 = ~sc_fail_r ? _GEN_1993 : valid_936; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3019 = ~sc_fail_r ? _GEN_1994 : valid_937; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3020 = ~sc_fail_r ? _GEN_1995 : valid_938; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3021 = ~sc_fail_r ? _GEN_1996 : valid_939; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3022 = ~sc_fail_r ? _GEN_1997 : valid_940; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3023 = ~sc_fail_r ? _GEN_1998 : valid_941; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3024 = ~sc_fail_r ? _GEN_1999 : valid_942; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3025 = ~sc_fail_r ? _GEN_2000 : valid_943; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3026 = ~sc_fail_r ? _GEN_2001 : valid_944; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3027 = ~sc_fail_r ? _GEN_2002 : valid_945; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3028 = ~sc_fail_r ? _GEN_2003 : valid_946; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3029 = ~sc_fail_r ? _GEN_2004 : valid_947; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3030 = ~sc_fail_r ? _GEN_2005 : valid_948; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3031 = ~sc_fail_r ? _GEN_2006 : valid_949; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3032 = ~sc_fail_r ? _GEN_2007 : valid_950; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3033 = ~sc_fail_r ? _GEN_2008 : valid_951; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3034 = ~sc_fail_r ? _GEN_2009 : valid_952; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3035 = ~sc_fail_r ? _GEN_2010 : valid_953; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3036 = ~sc_fail_r ? _GEN_2011 : valid_954; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3037 = ~sc_fail_r ? _GEN_2012 : valid_955; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3038 = ~sc_fail_r ? _GEN_2013 : valid_956; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3039 = ~sc_fail_r ? _GEN_2014 : valid_957; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3040 = ~sc_fail_r ? _GEN_2015 : valid_958; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3041 = ~sc_fail_r ? _GEN_2016 : valid_959; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3042 = ~sc_fail_r ? _GEN_2017 : valid_960; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3043 = ~sc_fail_r ? _GEN_2018 : valid_961; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3044 = ~sc_fail_r ? _GEN_2019 : valid_962; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3045 = ~sc_fail_r ? _GEN_2020 : valid_963; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3046 = ~sc_fail_r ? _GEN_2021 : valid_964; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3047 = ~sc_fail_r ? _GEN_2022 : valid_965; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3048 = ~sc_fail_r ? _GEN_2023 : valid_966; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3049 = ~sc_fail_r ? _GEN_2024 : valid_967; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3050 = ~sc_fail_r ? _GEN_2025 : valid_968; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3051 = ~sc_fail_r ? _GEN_2026 : valid_969; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3052 = ~sc_fail_r ? _GEN_2027 : valid_970; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3053 = ~sc_fail_r ? _GEN_2028 : valid_971; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3054 = ~sc_fail_r ? _GEN_2029 : valid_972; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3055 = ~sc_fail_r ? _GEN_2030 : valid_973; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3056 = ~sc_fail_r ? _GEN_2031 : valid_974; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3057 = ~sc_fail_r ? _GEN_2032 : valid_975; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3058 = ~sc_fail_r ? _GEN_2033 : valid_976; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3059 = ~sc_fail_r ? _GEN_2034 : valid_977; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3060 = ~sc_fail_r ? _GEN_2035 : valid_978; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3061 = ~sc_fail_r ? _GEN_2036 : valid_979; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3062 = ~sc_fail_r ? _GEN_2037 : valid_980; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3063 = ~sc_fail_r ? _GEN_2038 : valid_981; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3064 = ~sc_fail_r ? _GEN_2039 : valid_982; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3065 = ~sc_fail_r ? _GEN_2040 : valid_983; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3066 = ~sc_fail_r ? _GEN_2041 : valid_984; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3067 = ~sc_fail_r ? _GEN_2042 : valid_985; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3068 = ~sc_fail_r ? _GEN_2043 : valid_986; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3069 = ~sc_fail_r ? _GEN_2044 : valid_987; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3070 = ~sc_fail_r ? _GEN_2045 : valid_988; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3071 = ~sc_fail_r ? _GEN_2046 : valid_989; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3072 = ~sc_fail_r ? _GEN_2047 : valid_990; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3073 = ~sc_fail_r ? _GEN_2048 : valid_991; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3074 = ~sc_fail_r ? _GEN_2049 : valid_992; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3075 = ~sc_fail_r ? _GEN_2050 : valid_993; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3076 = ~sc_fail_r ? _GEN_2051 : valid_994; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3077 = ~sc_fail_r ? _GEN_2052 : valid_995; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3078 = ~sc_fail_r ? _GEN_2053 : valid_996; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3079 = ~sc_fail_r ? _GEN_2054 : valid_997; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3080 = ~sc_fail_r ? _GEN_2055 : valid_998; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3081 = ~sc_fail_r ? _GEN_2056 : valid_999; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3082 = ~sc_fail_r ? _GEN_2057 : valid_1000; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3083 = ~sc_fail_r ? _GEN_2058 : valid_1001; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3084 = ~sc_fail_r ? _GEN_2059 : valid_1002; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3085 = ~sc_fail_r ? _GEN_2060 : valid_1003; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3086 = ~sc_fail_r ? _GEN_2061 : valid_1004; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3087 = ~sc_fail_r ? _GEN_2062 : valid_1005; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3088 = ~sc_fail_r ? _GEN_2063 : valid_1006; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3089 = ~sc_fail_r ? _GEN_2064 : valid_1007; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3090 = ~sc_fail_r ? _GEN_2065 : valid_1008; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3091 = ~sc_fail_r ? _GEN_2066 : valid_1009; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3092 = ~sc_fail_r ? _GEN_2067 : valid_1010; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3093 = ~sc_fail_r ? _GEN_2068 : valid_1011; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3094 = ~sc_fail_r ? _GEN_2069 : valid_1012; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3095 = ~sc_fail_r ? _GEN_2070 : valid_1013; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3096 = ~sc_fail_r ? _GEN_2071 : valid_1014; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3097 = ~sc_fail_r ? _GEN_2072 : valid_1015; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3098 = ~sc_fail_r ? _GEN_2073 : valid_1016; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3099 = ~sc_fail_r ? _GEN_2074 : valid_1017; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3100 = ~sc_fail_r ? _GEN_2075 : valid_1018; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3101 = ~sc_fail_r ? _GEN_2076 : valid_1019; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3102 = ~sc_fail_r ? _GEN_2077 : valid_1020; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3103 = ~sc_fail_r ? _GEN_2078 : valid_1021; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3104 = ~sc_fail_r ? _GEN_2079 : valid_1022; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3105 = ~sc_fail_r ? _GEN_2080 : valid_1023; // @[DCache.scala 171:24 56:22]
  wire  _GEN_3107 = state == 3'h7 ? _T_12 : req_r_wen & array_hit; // @[DCache.scala 165:26 177:24]
  wire  _GEN_3108 = state == 3'h7 ? _GEN_2082 : valid_0; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3109 = state == 3'h7 ? _GEN_2083 : valid_1; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3110 = state == 3'h7 ? _GEN_2084 : valid_2; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3111 = state == 3'h7 ? _GEN_2085 : valid_3; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3112 = state == 3'h7 ? _GEN_2086 : valid_4; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3113 = state == 3'h7 ? _GEN_2087 : valid_5; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3114 = state == 3'h7 ? _GEN_2088 : valid_6; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3115 = state == 3'h7 ? _GEN_2089 : valid_7; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3116 = state == 3'h7 ? _GEN_2090 : valid_8; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3117 = state == 3'h7 ? _GEN_2091 : valid_9; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3118 = state == 3'h7 ? _GEN_2092 : valid_10; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3119 = state == 3'h7 ? _GEN_2093 : valid_11; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3120 = state == 3'h7 ? _GEN_2094 : valid_12; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3121 = state == 3'h7 ? _GEN_2095 : valid_13; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3122 = state == 3'h7 ? _GEN_2096 : valid_14; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3123 = state == 3'h7 ? _GEN_2097 : valid_15; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3124 = state == 3'h7 ? _GEN_2098 : valid_16; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3125 = state == 3'h7 ? _GEN_2099 : valid_17; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3126 = state == 3'h7 ? _GEN_2100 : valid_18; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3127 = state == 3'h7 ? _GEN_2101 : valid_19; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3128 = state == 3'h7 ? _GEN_2102 : valid_20; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3129 = state == 3'h7 ? _GEN_2103 : valid_21; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3130 = state == 3'h7 ? _GEN_2104 : valid_22; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3131 = state == 3'h7 ? _GEN_2105 : valid_23; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3132 = state == 3'h7 ? _GEN_2106 : valid_24; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3133 = state == 3'h7 ? _GEN_2107 : valid_25; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3134 = state == 3'h7 ? _GEN_2108 : valid_26; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3135 = state == 3'h7 ? _GEN_2109 : valid_27; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3136 = state == 3'h7 ? _GEN_2110 : valid_28; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3137 = state == 3'h7 ? _GEN_2111 : valid_29; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3138 = state == 3'h7 ? _GEN_2112 : valid_30; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3139 = state == 3'h7 ? _GEN_2113 : valid_31; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3140 = state == 3'h7 ? _GEN_2114 : valid_32; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3141 = state == 3'h7 ? _GEN_2115 : valid_33; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3142 = state == 3'h7 ? _GEN_2116 : valid_34; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3143 = state == 3'h7 ? _GEN_2117 : valid_35; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3144 = state == 3'h7 ? _GEN_2118 : valid_36; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3145 = state == 3'h7 ? _GEN_2119 : valid_37; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3146 = state == 3'h7 ? _GEN_2120 : valid_38; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3147 = state == 3'h7 ? _GEN_2121 : valid_39; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3148 = state == 3'h7 ? _GEN_2122 : valid_40; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3149 = state == 3'h7 ? _GEN_2123 : valid_41; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3150 = state == 3'h7 ? _GEN_2124 : valid_42; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3151 = state == 3'h7 ? _GEN_2125 : valid_43; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3152 = state == 3'h7 ? _GEN_2126 : valid_44; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3153 = state == 3'h7 ? _GEN_2127 : valid_45; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3154 = state == 3'h7 ? _GEN_2128 : valid_46; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3155 = state == 3'h7 ? _GEN_2129 : valid_47; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3156 = state == 3'h7 ? _GEN_2130 : valid_48; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3157 = state == 3'h7 ? _GEN_2131 : valid_49; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3158 = state == 3'h7 ? _GEN_2132 : valid_50; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3159 = state == 3'h7 ? _GEN_2133 : valid_51; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3160 = state == 3'h7 ? _GEN_2134 : valid_52; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3161 = state == 3'h7 ? _GEN_2135 : valid_53; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3162 = state == 3'h7 ? _GEN_2136 : valid_54; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3163 = state == 3'h7 ? _GEN_2137 : valid_55; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3164 = state == 3'h7 ? _GEN_2138 : valid_56; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3165 = state == 3'h7 ? _GEN_2139 : valid_57; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3166 = state == 3'h7 ? _GEN_2140 : valid_58; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3167 = state == 3'h7 ? _GEN_2141 : valid_59; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3168 = state == 3'h7 ? _GEN_2142 : valid_60; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3169 = state == 3'h7 ? _GEN_2143 : valid_61; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3170 = state == 3'h7 ? _GEN_2144 : valid_62; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3171 = state == 3'h7 ? _GEN_2145 : valid_63; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3172 = state == 3'h7 ? _GEN_2146 : valid_64; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3173 = state == 3'h7 ? _GEN_2147 : valid_65; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3174 = state == 3'h7 ? _GEN_2148 : valid_66; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3175 = state == 3'h7 ? _GEN_2149 : valid_67; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3176 = state == 3'h7 ? _GEN_2150 : valid_68; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3177 = state == 3'h7 ? _GEN_2151 : valid_69; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3178 = state == 3'h7 ? _GEN_2152 : valid_70; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3179 = state == 3'h7 ? _GEN_2153 : valid_71; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3180 = state == 3'h7 ? _GEN_2154 : valid_72; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3181 = state == 3'h7 ? _GEN_2155 : valid_73; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3182 = state == 3'h7 ? _GEN_2156 : valid_74; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3183 = state == 3'h7 ? _GEN_2157 : valid_75; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3184 = state == 3'h7 ? _GEN_2158 : valid_76; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3185 = state == 3'h7 ? _GEN_2159 : valid_77; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3186 = state == 3'h7 ? _GEN_2160 : valid_78; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3187 = state == 3'h7 ? _GEN_2161 : valid_79; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3188 = state == 3'h7 ? _GEN_2162 : valid_80; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3189 = state == 3'h7 ? _GEN_2163 : valid_81; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3190 = state == 3'h7 ? _GEN_2164 : valid_82; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3191 = state == 3'h7 ? _GEN_2165 : valid_83; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3192 = state == 3'h7 ? _GEN_2166 : valid_84; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3193 = state == 3'h7 ? _GEN_2167 : valid_85; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3194 = state == 3'h7 ? _GEN_2168 : valid_86; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3195 = state == 3'h7 ? _GEN_2169 : valid_87; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3196 = state == 3'h7 ? _GEN_2170 : valid_88; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3197 = state == 3'h7 ? _GEN_2171 : valid_89; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3198 = state == 3'h7 ? _GEN_2172 : valid_90; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3199 = state == 3'h7 ? _GEN_2173 : valid_91; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3200 = state == 3'h7 ? _GEN_2174 : valid_92; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3201 = state == 3'h7 ? _GEN_2175 : valid_93; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3202 = state == 3'h7 ? _GEN_2176 : valid_94; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3203 = state == 3'h7 ? _GEN_2177 : valid_95; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3204 = state == 3'h7 ? _GEN_2178 : valid_96; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3205 = state == 3'h7 ? _GEN_2179 : valid_97; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3206 = state == 3'h7 ? _GEN_2180 : valid_98; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3207 = state == 3'h7 ? _GEN_2181 : valid_99; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3208 = state == 3'h7 ? _GEN_2182 : valid_100; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3209 = state == 3'h7 ? _GEN_2183 : valid_101; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3210 = state == 3'h7 ? _GEN_2184 : valid_102; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3211 = state == 3'h7 ? _GEN_2185 : valid_103; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3212 = state == 3'h7 ? _GEN_2186 : valid_104; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3213 = state == 3'h7 ? _GEN_2187 : valid_105; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3214 = state == 3'h7 ? _GEN_2188 : valid_106; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3215 = state == 3'h7 ? _GEN_2189 : valid_107; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3216 = state == 3'h7 ? _GEN_2190 : valid_108; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3217 = state == 3'h7 ? _GEN_2191 : valid_109; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3218 = state == 3'h7 ? _GEN_2192 : valid_110; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3219 = state == 3'h7 ? _GEN_2193 : valid_111; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3220 = state == 3'h7 ? _GEN_2194 : valid_112; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3221 = state == 3'h7 ? _GEN_2195 : valid_113; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3222 = state == 3'h7 ? _GEN_2196 : valid_114; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3223 = state == 3'h7 ? _GEN_2197 : valid_115; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3224 = state == 3'h7 ? _GEN_2198 : valid_116; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3225 = state == 3'h7 ? _GEN_2199 : valid_117; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3226 = state == 3'h7 ? _GEN_2200 : valid_118; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3227 = state == 3'h7 ? _GEN_2201 : valid_119; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3228 = state == 3'h7 ? _GEN_2202 : valid_120; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3229 = state == 3'h7 ? _GEN_2203 : valid_121; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3230 = state == 3'h7 ? _GEN_2204 : valid_122; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3231 = state == 3'h7 ? _GEN_2205 : valid_123; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3232 = state == 3'h7 ? _GEN_2206 : valid_124; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3233 = state == 3'h7 ? _GEN_2207 : valid_125; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3234 = state == 3'h7 ? _GEN_2208 : valid_126; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3235 = state == 3'h7 ? _GEN_2209 : valid_127; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3236 = state == 3'h7 ? _GEN_2210 : valid_128; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3237 = state == 3'h7 ? _GEN_2211 : valid_129; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3238 = state == 3'h7 ? _GEN_2212 : valid_130; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3239 = state == 3'h7 ? _GEN_2213 : valid_131; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3240 = state == 3'h7 ? _GEN_2214 : valid_132; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3241 = state == 3'h7 ? _GEN_2215 : valid_133; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3242 = state == 3'h7 ? _GEN_2216 : valid_134; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3243 = state == 3'h7 ? _GEN_2217 : valid_135; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3244 = state == 3'h7 ? _GEN_2218 : valid_136; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3245 = state == 3'h7 ? _GEN_2219 : valid_137; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3246 = state == 3'h7 ? _GEN_2220 : valid_138; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3247 = state == 3'h7 ? _GEN_2221 : valid_139; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3248 = state == 3'h7 ? _GEN_2222 : valid_140; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3249 = state == 3'h7 ? _GEN_2223 : valid_141; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3250 = state == 3'h7 ? _GEN_2224 : valid_142; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3251 = state == 3'h7 ? _GEN_2225 : valid_143; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3252 = state == 3'h7 ? _GEN_2226 : valid_144; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3253 = state == 3'h7 ? _GEN_2227 : valid_145; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3254 = state == 3'h7 ? _GEN_2228 : valid_146; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3255 = state == 3'h7 ? _GEN_2229 : valid_147; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3256 = state == 3'h7 ? _GEN_2230 : valid_148; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3257 = state == 3'h7 ? _GEN_2231 : valid_149; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3258 = state == 3'h7 ? _GEN_2232 : valid_150; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3259 = state == 3'h7 ? _GEN_2233 : valid_151; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3260 = state == 3'h7 ? _GEN_2234 : valid_152; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3261 = state == 3'h7 ? _GEN_2235 : valid_153; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3262 = state == 3'h7 ? _GEN_2236 : valid_154; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3263 = state == 3'h7 ? _GEN_2237 : valid_155; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3264 = state == 3'h7 ? _GEN_2238 : valid_156; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3265 = state == 3'h7 ? _GEN_2239 : valid_157; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3266 = state == 3'h7 ? _GEN_2240 : valid_158; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3267 = state == 3'h7 ? _GEN_2241 : valid_159; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3268 = state == 3'h7 ? _GEN_2242 : valid_160; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3269 = state == 3'h7 ? _GEN_2243 : valid_161; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3270 = state == 3'h7 ? _GEN_2244 : valid_162; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3271 = state == 3'h7 ? _GEN_2245 : valid_163; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3272 = state == 3'h7 ? _GEN_2246 : valid_164; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3273 = state == 3'h7 ? _GEN_2247 : valid_165; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3274 = state == 3'h7 ? _GEN_2248 : valid_166; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3275 = state == 3'h7 ? _GEN_2249 : valid_167; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3276 = state == 3'h7 ? _GEN_2250 : valid_168; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3277 = state == 3'h7 ? _GEN_2251 : valid_169; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3278 = state == 3'h7 ? _GEN_2252 : valid_170; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3279 = state == 3'h7 ? _GEN_2253 : valid_171; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3280 = state == 3'h7 ? _GEN_2254 : valid_172; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3281 = state == 3'h7 ? _GEN_2255 : valid_173; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3282 = state == 3'h7 ? _GEN_2256 : valid_174; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3283 = state == 3'h7 ? _GEN_2257 : valid_175; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3284 = state == 3'h7 ? _GEN_2258 : valid_176; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3285 = state == 3'h7 ? _GEN_2259 : valid_177; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3286 = state == 3'h7 ? _GEN_2260 : valid_178; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3287 = state == 3'h7 ? _GEN_2261 : valid_179; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3288 = state == 3'h7 ? _GEN_2262 : valid_180; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3289 = state == 3'h7 ? _GEN_2263 : valid_181; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3290 = state == 3'h7 ? _GEN_2264 : valid_182; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3291 = state == 3'h7 ? _GEN_2265 : valid_183; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3292 = state == 3'h7 ? _GEN_2266 : valid_184; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3293 = state == 3'h7 ? _GEN_2267 : valid_185; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3294 = state == 3'h7 ? _GEN_2268 : valid_186; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3295 = state == 3'h7 ? _GEN_2269 : valid_187; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3296 = state == 3'h7 ? _GEN_2270 : valid_188; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3297 = state == 3'h7 ? _GEN_2271 : valid_189; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3298 = state == 3'h7 ? _GEN_2272 : valid_190; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3299 = state == 3'h7 ? _GEN_2273 : valid_191; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3300 = state == 3'h7 ? _GEN_2274 : valid_192; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3301 = state == 3'h7 ? _GEN_2275 : valid_193; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3302 = state == 3'h7 ? _GEN_2276 : valid_194; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3303 = state == 3'h7 ? _GEN_2277 : valid_195; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3304 = state == 3'h7 ? _GEN_2278 : valid_196; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3305 = state == 3'h7 ? _GEN_2279 : valid_197; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3306 = state == 3'h7 ? _GEN_2280 : valid_198; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3307 = state == 3'h7 ? _GEN_2281 : valid_199; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3308 = state == 3'h7 ? _GEN_2282 : valid_200; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3309 = state == 3'h7 ? _GEN_2283 : valid_201; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3310 = state == 3'h7 ? _GEN_2284 : valid_202; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3311 = state == 3'h7 ? _GEN_2285 : valid_203; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3312 = state == 3'h7 ? _GEN_2286 : valid_204; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3313 = state == 3'h7 ? _GEN_2287 : valid_205; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3314 = state == 3'h7 ? _GEN_2288 : valid_206; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3315 = state == 3'h7 ? _GEN_2289 : valid_207; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3316 = state == 3'h7 ? _GEN_2290 : valid_208; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3317 = state == 3'h7 ? _GEN_2291 : valid_209; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3318 = state == 3'h7 ? _GEN_2292 : valid_210; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3319 = state == 3'h7 ? _GEN_2293 : valid_211; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3320 = state == 3'h7 ? _GEN_2294 : valid_212; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3321 = state == 3'h7 ? _GEN_2295 : valid_213; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3322 = state == 3'h7 ? _GEN_2296 : valid_214; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3323 = state == 3'h7 ? _GEN_2297 : valid_215; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3324 = state == 3'h7 ? _GEN_2298 : valid_216; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3325 = state == 3'h7 ? _GEN_2299 : valid_217; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3326 = state == 3'h7 ? _GEN_2300 : valid_218; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3327 = state == 3'h7 ? _GEN_2301 : valid_219; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3328 = state == 3'h7 ? _GEN_2302 : valid_220; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3329 = state == 3'h7 ? _GEN_2303 : valid_221; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3330 = state == 3'h7 ? _GEN_2304 : valid_222; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3331 = state == 3'h7 ? _GEN_2305 : valid_223; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3332 = state == 3'h7 ? _GEN_2306 : valid_224; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3333 = state == 3'h7 ? _GEN_2307 : valid_225; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3334 = state == 3'h7 ? _GEN_2308 : valid_226; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3335 = state == 3'h7 ? _GEN_2309 : valid_227; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3336 = state == 3'h7 ? _GEN_2310 : valid_228; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3337 = state == 3'h7 ? _GEN_2311 : valid_229; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3338 = state == 3'h7 ? _GEN_2312 : valid_230; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3339 = state == 3'h7 ? _GEN_2313 : valid_231; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3340 = state == 3'h7 ? _GEN_2314 : valid_232; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3341 = state == 3'h7 ? _GEN_2315 : valid_233; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3342 = state == 3'h7 ? _GEN_2316 : valid_234; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3343 = state == 3'h7 ? _GEN_2317 : valid_235; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3344 = state == 3'h7 ? _GEN_2318 : valid_236; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3345 = state == 3'h7 ? _GEN_2319 : valid_237; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3346 = state == 3'h7 ? _GEN_2320 : valid_238; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3347 = state == 3'h7 ? _GEN_2321 : valid_239; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3348 = state == 3'h7 ? _GEN_2322 : valid_240; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3349 = state == 3'h7 ? _GEN_2323 : valid_241; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3350 = state == 3'h7 ? _GEN_2324 : valid_242; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3351 = state == 3'h7 ? _GEN_2325 : valid_243; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3352 = state == 3'h7 ? _GEN_2326 : valid_244; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3353 = state == 3'h7 ? _GEN_2327 : valid_245; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3354 = state == 3'h7 ? _GEN_2328 : valid_246; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3355 = state == 3'h7 ? _GEN_2329 : valid_247; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3356 = state == 3'h7 ? _GEN_2330 : valid_248; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3357 = state == 3'h7 ? _GEN_2331 : valid_249; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3358 = state == 3'h7 ? _GEN_2332 : valid_250; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3359 = state == 3'h7 ? _GEN_2333 : valid_251; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3360 = state == 3'h7 ? _GEN_2334 : valid_252; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3361 = state == 3'h7 ? _GEN_2335 : valid_253; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3362 = state == 3'h7 ? _GEN_2336 : valid_254; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3363 = state == 3'h7 ? _GEN_2337 : valid_255; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3364 = state == 3'h7 ? _GEN_2338 : valid_256; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3365 = state == 3'h7 ? _GEN_2339 : valid_257; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3366 = state == 3'h7 ? _GEN_2340 : valid_258; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3367 = state == 3'h7 ? _GEN_2341 : valid_259; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3368 = state == 3'h7 ? _GEN_2342 : valid_260; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3369 = state == 3'h7 ? _GEN_2343 : valid_261; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3370 = state == 3'h7 ? _GEN_2344 : valid_262; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3371 = state == 3'h7 ? _GEN_2345 : valid_263; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3372 = state == 3'h7 ? _GEN_2346 : valid_264; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3373 = state == 3'h7 ? _GEN_2347 : valid_265; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3374 = state == 3'h7 ? _GEN_2348 : valid_266; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3375 = state == 3'h7 ? _GEN_2349 : valid_267; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3376 = state == 3'h7 ? _GEN_2350 : valid_268; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3377 = state == 3'h7 ? _GEN_2351 : valid_269; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3378 = state == 3'h7 ? _GEN_2352 : valid_270; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3379 = state == 3'h7 ? _GEN_2353 : valid_271; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3380 = state == 3'h7 ? _GEN_2354 : valid_272; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3381 = state == 3'h7 ? _GEN_2355 : valid_273; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3382 = state == 3'h7 ? _GEN_2356 : valid_274; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3383 = state == 3'h7 ? _GEN_2357 : valid_275; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3384 = state == 3'h7 ? _GEN_2358 : valid_276; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3385 = state == 3'h7 ? _GEN_2359 : valid_277; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3386 = state == 3'h7 ? _GEN_2360 : valid_278; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3387 = state == 3'h7 ? _GEN_2361 : valid_279; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3388 = state == 3'h7 ? _GEN_2362 : valid_280; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3389 = state == 3'h7 ? _GEN_2363 : valid_281; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3390 = state == 3'h7 ? _GEN_2364 : valid_282; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3391 = state == 3'h7 ? _GEN_2365 : valid_283; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3392 = state == 3'h7 ? _GEN_2366 : valid_284; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3393 = state == 3'h7 ? _GEN_2367 : valid_285; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3394 = state == 3'h7 ? _GEN_2368 : valid_286; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3395 = state == 3'h7 ? _GEN_2369 : valid_287; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3396 = state == 3'h7 ? _GEN_2370 : valid_288; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3397 = state == 3'h7 ? _GEN_2371 : valid_289; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3398 = state == 3'h7 ? _GEN_2372 : valid_290; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3399 = state == 3'h7 ? _GEN_2373 : valid_291; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3400 = state == 3'h7 ? _GEN_2374 : valid_292; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3401 = state == 3'h7 ? _GEN_2375 : valid_293; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3402 = state == 3'h7 ? _GEN_2376 : valid_294; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3403 = state == 3'h7 ? _GEN_2377 : valid_295; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3404 = state == 3'h7 ? _GEN_2378 : valid_296; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3405 = state == 3'h7 ? _GEN_2379 : valid_297; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3406 = state == 3'h7 ? _GEN_2380 : valid_298; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3407 = state == 3'h7 ? _GEN_2381 : valid_299; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3408 = state == 3'h7 ? _GEN_2382 : valid_300; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3409 = state == 3'h7 ? _GEN_2383 : valid_301; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3410 = state == 3'h7 ? _GEN_2384 : valid_302; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3411 = state == 3'h7 ? _GEN_2385 : valid_303; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3412 = state == 3'h7 ? _GEN_2386 : valid_304; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3413 = state == 3'h7 ? _GEN_2387 : valid_305; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3414 = state == 3'h7 ? _GEN_2388 : valid_306; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3415 = state == 3'h7 ? _GEN_2389 : valid_307; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3416 = state == 3'h7 ? _GEN_2390 : valid_308; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3417 = state == 3'h7 ? _GEN_2391 : valid_309; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3418 = state == 3'h7 ? _GEN_2392 : valid_310; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3419 = state == 3'h7 ? _GEN_2393 : valid_311; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3420 = state == 3'h7 ? _GEN_2394 : valid_312; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3421 = state == 3'h7 ? _GEN_2395 : valid_313; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3422 = state == 3'h7 ? _GEN_2396 : valid_314; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3423 = state == 3'h7 ? _GEN_2397 : valid_315; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3424 = state == 3'h7 ? _GEN_2398 : valid_316; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3425 = state == 3'h7 ? _GEN_2399 : valid_317; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3426 = state == 3'h7 ? _GEN_2400 : valid_318; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3427 = state == 3'h7 ? _GEN_2401 : valid_319; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3428 = state == 3'h7 ? _GEN_2402 : valid_320; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3429 = state == 3'h7 ? _GEN_2403 : valid_321; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3430 = state == 3'h7 ? _GEN_2404 : valid_322; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3431 = state == 3'h7 ? _GEN_2405 : valid_323; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3432 = state == 3'h7 ? _GEN_2406 : valid_324; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3433 = state == 3'h7 ? _GEN_2407 : valid_325; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3434 = state == 3'h7 ? _GEN_2408 : valid_326; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3435 = state == 3'h7 ? _GEN_2409 : valid_327; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3436 = state == 3'h7 ? _GEN_2410 : valid_328; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3437 = state == 3'h7 ? _GEN_2411 : valid_329; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3438 = state == 3'h7 ? _GEN_2412 : valid_330; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3439 = state == 3'h7 ? _GEN_2413 : valid_331; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3440 = state == 3'h7 ? _GEN_2414 : valid_332; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3441 = state == 3'h7 ? _GEN_2415 : valid_333; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3442 = state == 3'h7 ? _GEN_2416 : valid_334; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3443 = state == 3'h7 ? _GEN_2417 : valid_335; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3444 = state == 3'h7 ? _GEN_2418 : valid_336; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3445 = state == 3'h7 ? _GEN_2419 : valid_337; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3446 = state == 3'h7 ? _GEN_2420 : valid_338; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3447 = state == 3'h7 ? _GEN_2421 : valid_339; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3448 = state == 3'h7 ? _GEN_2422 : valid_340; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3449 = state == 3'h7 ? _GEN_2423 : valid_341; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3450 = state == 3'h7 ? _GEN_2424 : valid_342; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3451 = state == 3'h7 ? _GEN_2425 : valid_343; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3452 = state == 3'h7 ? _GEN_2426 : valid_344; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3453 = state == 3'h7 ? _GEN_2427 : valid_345; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3454 = state == 3'h7 ? _GEN_2428 : valid_346; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3455 = state == 3'h7 ? _GEN_2429 : valid_347; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3456 = state == 3'h7 ? _GEN_2430 : valid_348; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3457 = state == 3'h7 ? _GEN_2431 : valid_349; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3458 = state == 3'h7 ? _GEN_2432 : valid_350; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3459 = state == 3'h7 ? _GEN_2433 : valid_351; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3460 = state == 3'h7 ? _GEN_2434 : valid_352; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3461 = state == 3'h7 ? _GEN_2435 : valid_353; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3462 = state == 3'h7 ? _GEN_2436 : valid_354; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3463 = state == 3'h7 ? _GEN_2437 : valid_355; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3464 = state == 3'h7 ? _GEN_2438 : valid_356; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3465 = state == 3'h7 ? _GEN_2439 : valid_357; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3466 = state == 3'h7 ? _GEN_2440 : valid_358; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3467 = state == 3'h7 ? _GEN_2441 : valid_359; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3468 = state == 3'h7 ? _GEN_2442 : valid_360; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3469 = state == 3'h7 ? _GEN_2443 : valid_361; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3470 = state == 3'h7 ? _GEN_2444 : valid_362; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3471 = state == 3'h7 ? _GEN_2445 : valid_363; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3472 = state == 3'h7 ? _GEN_2446 : valid_364; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3473 = state == 3'h7 ? _GEN_2447 : valid_365; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3474 = state == 3'h7 ? _GEN_2448 : valid_366; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3475 = state == 3'h7 ? _GEN_2449 : valid_367; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3476 = state == 3'h7 ? _GEN_2450 : valid_368; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3477 = state == 3'h7 ? _GEN_2451 : valid_369; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3478 = state == 3'h7 ? _GEN_2452 : valid_370; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3479 = state == 3'h7 ? _GEN_2453 : valid_371; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3480 = state == 3'h7 ? _GEN_2454 : valid_372; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3481 = state == 3'h7 ? _GEN_2455 : valid_373; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3482 = state == 3'h7 ? _GEN_2456 : valid_374; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3483 = state == 3'h7 ? _GEN_2457 : valid_375; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3484 = state == 3'h7 ? _GEN_2458 : valid_376; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3485 = state == 3'h7 ? _GEN_2459 : valid_377; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3486 = state == 3'h7 ? _GEN_2460 : valid_378; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3487 = state == 3'h7 ? _GEN_2461 : valid_379; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3488 = state == 3'h7 ? _GEN_2462 : valid_380; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3489 = state == 3'h7 ? _GEN_2463 : valid_381; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3490 = state == 3'h7 ? _GEN_2464 : valid_382; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3491 = state == 3'h7 ? _GEN_2465 : valid_383; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3492 = state == 3'h7 ? _GEN_2466 : valid_384; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3493 = state == 3'h7 ? _GEN_2467 : valid_385; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3494 = state == 3'h7 ? _GEN_2468 : valid_386; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3495 = state == 3'h7 ? _GEN_2469 : valid_387; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3496 = state == 3'h7 ? _GEN_2470 : valid_388; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3497 = state == 3'h7 ? _GEN_2471 : valid_389; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3498 = state == 3'h7 ? _GEN_2472 : valid_390; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3499 = state == 3'h7 ? _GEN_2473 : valid_391; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3500 = state == 3'h7 ? _GEN_2474 : valid_392; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3501 = state == 3'h7 ? _GEN_2475 : valid_393; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3502 = state == 3'h7 ? _GEN_2476 : valid_394; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3503 = state == 3'h7 ? _GEN_2477 : valid_395; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3504 = state == 3'h7 ? _GEN_2478 : valid_396; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3505 = state == 3'h7 ? _GEN_2479 : valid_397; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3506 = state == 3'h7 ? _GEN_2480 : valid_398; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3507 = state == 3'h7 ? _GEN_2481 : valid_399; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3508 = state == 3'h7 ? _GEN_2482 : valid_400; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3509 = state == 3'h7 ? _GEN_2483 : valid_401; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3510 = state == 3'h7 ? _GEN_2484 : valid_402; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3511 = state == 3'h7 ? _GEN_2485 : valid_403; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3512 = state == 3'h7 ? _GEN_2486 : valid_404; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3513 = state == 3'h7 ? _GEN_2487 : valid_405; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3514 = state == 3'h7 ? _GEN_2488 : valid_406; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3515 = state == 3'h7 ? _GEN_2489 : valid_407; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3516 = state == 3'h7 ? _GEN_2490 : valid_408; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3517 = state == 3'h7 ? _GEN_2491 : valid_409; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3518 = state == 3'h7 ? _GEN_2492 : valid_410; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3519 = state == 3'h7 ? _GEN_2493 : valid_411; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3520 = state == 3'h7 ? _GEN_2494 : valid_412; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3521 = state == 3'h7 ? _GEN_2495 : valid_413; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3522 = state == 3'h7 ? _GEN_2496 : valid_414; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3523 = state == 3'h7 ? _GEN_2497 : valid_415; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3524 = state == 3'h7 ? _GEN_2498 : valid_416; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3525 = state == 3'h7 ? _GEN_2499 : valid_417; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3526 = state == 3'h7 ? _GEN_2500 : valid_418; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3527 = state == 3'h7 ? _GEN_2501 : valid_419; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3528 = state == 3'h7 ? _GEN_2502 : valid_420; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3529 = state == 3'h7 ? _GEN_2503 : valid_421; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3530 = state == 3'h7 ? _GEN_2504 : valid_422; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3531 = state == 3'h7 ? _GEN_2505 : valid_423; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3532 = state == 3'h7 ? _GEN_2506 : valid_424; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3533 = state == 3'h7 ? _GEN_2507 : valid_425; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3534 = state == 3'h7 ? _GEN_2508 : valid_426; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3535 = state == 3'h7 ? _GEN_2509 : valid_427; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3536 = state == 3'h7 ? _GEN_2510 : valid_428; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3537 = state == 3'h7 ? _GEN_2511 : valid_429; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3538 = state == 3'h7 ? _GEN_2512 : valid_430; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3539 = state == 3'h7 ? _GEN_2513 : valid_431; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3540 = state == 3'h7 ? _GEN_2514 : valid_432; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3541 = state == 3'h7 ? _GEN_2515 : valid_433; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3542 = state == 3'h7 ? _GEN_2516 : valid_434; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3543 = state == 3'h7 ? _GEN_2517 : valid_435; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3544 = state == 3'h7 ? _GEN_2518 : valid_436; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3545 = state == 3'h7 ? _GEN_2519 : valid_437; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3546 = state == 3'h7 ? _GEN_2520 : valid_438; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3547 = state == 3'h7 ? _GEN_2521 : valid_439; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3548 = state == 3'h7 ? _GEN_2522 : valid_440; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3549 = state == 3'h7 ? _GEN_2523 : valid_441; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3550 = state == 3'h7 ? _GEN_2524 : valid_442; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3551 = state == 3'h7 ? _GEN_2525 : valid_443; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3552 = state == 3'h7 ? _GEN_2526 : valid_444; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3553 = state == 3'h7 ? _GEN_2527 : valid_445; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3554 = state == 3'h7 ? _GEN_2528 : valid_446; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3555 = state == 3'h7 ? _GEN_2529 : valid_447; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3556 = state == 3'h7 ? _GEN_2530 : valid_448; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3557 = state == 3'h7 ? _GEN_2531 : valid_449; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3558 = state == 3'h7 ? _GEN_2532 : valid_450; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3559 = state == 3'h7 ? _GEN_2533 : valid_451; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3560 = state == 3'h7 ? _GEN_2534 : valid_452; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3561 = state == 3'h7 ? _GEN_2535 : valid_453; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3562 = state == 3'h7 ? _GEN_2536 : valid_454; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3563 = state == 3'h7 ? _GEN_2537 : valid_455; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3564 = state == 3'h7 ? _GEN_2538 : valid_456; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3565 = state == 3'h7 ? _GEN_2539 : valid_457; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3566 = state == 3'h7 ? _GEN_2540 : valid_458; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3567 = state == 3'h7 ? _GEN_2541 : valid_459; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3568 = state == 3'h7 ? _GEN_2542 : valid_460; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3569 = state == 3'h7 ? _GEN_2543 : valid_461; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3570 = state == 3'h7 ? _GEN_2544 : valid_462; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3571 = state == 3'h7 ? _GEN_2545 : valid_463; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3572 = state == 3'h7 ? _GEN_2546 : valid_464; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3573 = state == 3'h7 ? _GEN_2547 : valid_465; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3574 = state == 3'h7 ? _GEN_2548 : valid_466; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3575 = state == 3'h7 ? _GEN_2549 : valid_467; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3576 = state == 3'h7 ? _GEN_2550 : valid_468; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3577 = state == 3'h7 ? _GEN_2551 : valid_469; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3578 = state == 3'h7 ? _GEN_2552 : valid_470; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3579 = state == 3'h7 ? _GEN_2553 : valid_471; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3580 = state == 3'h7 ? _GEN_2554 : valid_472; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3581 = state == 3'h7 ? _GEN_2555 : valid_473; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3582 = state == 3'h7 ? _GEN_2556 : valid_474; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3583 = state == 3'h7 ? _GEN_2557 : valid_475; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3584 = state == 3'h7 ? _GEN_2558 : valid_476; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3585 = state == 3'h7 ? _GEN_2559 : valid_477; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3586 = state == 3'h7 ? _GEN_2560 : valid_478; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3587 = state == 3'h7 ? _GEN_2561 : valid_479; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3588 = state == 3'h7 ? _GEN_2562 : valid_480; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3589 = state == 3'h7 ? _GEN_2563 : valid_481; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3590 = state == 3'h7 ? _GEN_2564 : valid_482; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3591 = state == 3'h7 ? _GEN_2565 : valid_483; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3592 = state == 3'h7 ? _GEN_2566 : valid_484; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3593 = state == 3'h7 ? _GEN_2567 : valid_485; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3594 = state == 3'h7 ? _GEN_2568 : valid_486; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3595 = state == 3'h7 ? _GEN_2569 : valid_487; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3596 = state == 3'h7 ? _GEN_2570 : valid_488; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3597 = state == 3'h7 ? _GEN_2571 : valid_489; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3598 = state == 3'h7 ? _GEN_2572 : valid_490; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3599 = state == 3'h7 ? _GEN_2573 : valid_491; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3600 = state == 3'h7 ? _GEN_2574 : valid_492; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3601 = state == 3'h7 ? _GEN_2575 : valid_493; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3602 = state == 3'h7 ? _GEN_2576 : valid_494; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3603 = state == 3'h7 ? _GEN_2577 : valid_495; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3604 = state == 3'h7 ? _GEN_2578 : valid_496; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3605 = state == 3'h7 ? _GEN_2579 : valid_497; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3606 = state == 3'h7 ? _GEN_2580 : valid_498; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3607 = state == 3'h7 ? _GEN_2581 : valid_499; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3608 = state == 3'h7 ? _GEN_2582 : valid_500; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3609 = state == 3'h7 ? _GEN_2583 : valid_501; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3610 = state == 3'h7 ? _GEN_2584 : valid_502; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3611 = state == 3'h7 ? _GEN_2585 : valid_503; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3612 = state == 3'h7 ? _GEN_2586 : valid_504; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3613 = state == 3'h7 ? _GEN_2587 : valid_505; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3614 = state == 3'h7 ? _GEN_2588 : valid_506; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3615 = state == 3'h7 ? _GEN_2589 : valid_507; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3616 = state == 3'h7 ? _GEN_2590 : valid_508; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3617 = state == 3'h7 ? _GEN_2591 : valid_509; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3618 = state == 3'h7 ? _GEN_2592 : valid_510; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3619 = state == 3'h7 ? _GEN_2593 : valid_511; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3620 = state == 3'h7 ? _GEN_2594 : valid_512; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3621 = state == 3'h7 ? _GEN_2595 : valid_513; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3622 = state == 3'h7 ? _GEN_2596 : valid_514; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3623 = state == 3'h7 ? _GEN_2597 : valid_515; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3624 = state == 3'h7 ? _GEN_2598 : valid_516; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3625 = state == 3'h7 ? _GEN_2599 : valid_517; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3626 = state == 3'h7 ? _GEN_2600 : valid_518; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3627 = state == 3'h7 ? _GEN_2601 : valid_519; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3628 = state == 3'h7 ? _GEN_2602 : valid_520; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3629 = state == 3'h7 ? _GEN_2603 : valid_521; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3630 = state == 3'h7 ? _GEN_2604 : valid_522; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3631 = state == 3'h7 ? _GEN_2605 : valid_523; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3632 = state == 3'h7 ? _GEN_2606 : valid_524; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3633 = state == 3'h7 ? _GEN_2607 : valid_525; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3634 = state == 3'h7 ? _GEN_2608 : valid_526; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3635 = state == 3'h7 ? _GEN_2609 : valid_527; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3636 = state == 3'h7 ? _GEN_2610 : valid_528; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3637 = state == 3'h7 ? _GEN_2611 : valid_529; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3638 = state == 3'h7 ? _GEN_2612 : valid_530; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3639 = state == 3'h7 ? _GEN_2613 : valid_531; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3640 = state == 3'h7 ? _GEN_2614 : valid_532; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3641 = state == 3'h7 ? _GEN_2615 : valid_533; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3642 = state == 3'h7 ? _GEN_2616 : valid_534; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3643 = state == 3'h7 ? _GEN_2617 : valid_535; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3644 = state == 3'h7 ? _GEN_2618 : valid_536; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3645 = state == 3'h7 ? _GEN_2619 : valid_537; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3646 = state == 3'h7 ? _GEN_2620 : valid_538; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3647 = state == 3'h7 ? _GEN_2621 : valid_539; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3648 = state == 3'h7 ? _GEN_2622 : valid_540; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3649 = state == 3'h7 ? _GEN_2623 : valid_541; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3650 = state == 3'h7 ? _GEN_2624 : valid_542; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3651 = state == 3'h7 ? _GEN_2625 : valid_543; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3652 = state == 3'h7 ? _GEN_2626 : valid_544; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3653 = state == 3'h7 ? _GEN_2627 : valid_545; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3654 = state == 3'h7 ? _GEN_2628 : valid_546; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3655 = state == 3'h7 ? _GEN_2629 : valid_547; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3656 = state == 3'h7 ? _GEN_2630 : valid_548; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3657 = state == 3'h7 ? _GEN_2631 : valid_549; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3658 = state == 3'h7 ? _GEN_2632 : valid_550; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3659 = state == 3'h7 ? _GEN_2633 : valid_551; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3660 = state == 3'h7 ? _GEN_2634 : valid_552; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3661 = state == 3'h7 ? _GEN_2635 : valid_553; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3662 = state == 3'h7 ? _GEN_2636 : valid_554; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3663 = state == 3'h7 ? _GEN_2637 : valid_555; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3664 = state == 3'h7 ? _GEN_2638 : valid_556; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3665 = state == 3'h7 ? _GEN_2639 : valid_557; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3666 = state == 3'h7 ? _GEN_2640 : valid_558; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3667 = state == 3'h7 ? _GEN_2641 : valid_559; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3668 = state == 3'h7 ? _GEN_2642 : valid_560; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3669 = state == 3'h7 ? _GEN_2643 : valid_561; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3670 = state == 3'h7 ? _GEN_2644 : valid_562; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3671 = state == 3'h7 ? _GEN_2645 : valid_563; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3672 = state == 3'h7 ? _GEN_2646 : valid_564; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3673 = state == 3'h7 ? _GEN_2647 : valid_565; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3674 = state == 3'h7 ? _GEN_2648 : valid_566; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3675 = state == 3'h7 ? _GEN_2649 : valid_567; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3676 = state == 3'h7 ? _GEN_2650 : valid_568; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3677 = state == 3'h7 ? _GEN_2651 : valid_569; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3678 = state == 3'h7 ? _GEN_2652 : valid_570; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3679 = state == 3'h7 ? _GEN_2653 : valid_571; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3680 = state == 3'h7 ? _GEN_2654 : valid_572; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3681 = state == 3'h7 ? _GEN_2655 : valid_573; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3682 = state == 3'h7 ? _GEN_2656 : valid_574; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3683 = state == 3'h7 ? _GEN_2657 : valid_575; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3684 = state == 3'h7 ? _GEN_2658 : valid_576; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3685 = state == 3'h7 ? _GEN_2659 : valid_577; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3686 = state == 3'h7 ? _GEN_2660 : valid_578; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3687 = state == 3'h7 ? _GEN_2661 : valid_579; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3688 = state == 3'h7 ? _GEN_2662 : valid_580; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3689 = state == 3'h7 ? _GEN_2663 : valid_581; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3690 = state == 3'h7 ? _GEN_2664 : valid_582; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3691 = state == 3'h7 ? _GEN_2665 : valid_583; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3692 = state == 3'h7 ? _GEN_2666 : valid_584; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3693 = state == 3'h7 ? _GEN_2667 : valid_585; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3694 = state == 3'h7 ? _GEN_2668 : valid_586; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3695 = state == 3'h7 ? _GEN_2669 : valid_587; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3696 = state == 3'h7 ? _GEN_2670 : valid_588; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3697 = state == 3'h7 ? _GEN_2671 : valid_589; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3698 = state == 3'h7 ? _GEN_2672 : valid_590; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3699 = state == 3'h7 ? _GEN_2673 : valid_591; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3700 = state == 3'h7 ? _GEN_2674 : valid_592; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3701 = state == 3'h7 ? _GEN_2675 : valid_593; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3702 = state == 3'h7 ? _GEN_2676 : valid_594; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3703 = state == 3'h7 ? _GEN_2677 : valid_595; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3704 = state == 3'h7 ? _GEN_2678 : valid_596; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3705 = state == 3'h7 ? _GEN_2679 : valid_597; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3706 = state == 3'h7 ? _GEN_2680 : valid_598; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3707 = state == 3'h7 ? _GEN_2681 : valid_599; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3708 = state == 3'h7 ? _GEN_2682 : valid_600; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3709 = state == 3'h7 ? _GEN_2683 : valid_601; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3710 = state == 3'h7 ? _GEN_2684 : valid_602; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3711 = state == 3'h7 ? _GEN_2685 : valid_603; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3712 = state == 3'h7 ? _GEN_2686 : valid_604; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3713 = state == 3'h7 ? _GEN_2687 : valid_605; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3714 = state == 3'h7 ? _GEN_2688 : valid_606; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3715 = state == 3'h7 ? _GEN_2689 : valid_607; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3716 = state == 3'h7 ? _GEN_2690 : valid_608; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3717 = state == 3'h7 ? _GEN_2691 : valid_609; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3718 = state == 3'h7 ? _GEN_2692 : valid_610; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3719 = state == 3'h7 ? _GEN_2693 : valid_611; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3720 = state == 3'h7 ? _GEN_2694 : valid_612; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3721 = state == 3'h7 ? _GEN_2695 : valid_613; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3722 = state == 3'h7 ? _GEN_2696 : valid_614; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3723 = state == 3'h7 ? _GEN_2697 : valid_615; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3724 = state == 3'h7 ? _GEN_2698 : valid_616; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3725 = state == 3'h7 ? _GEN_2699 : valid_617; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3726 = state == 3'h7 ? _GEN_2700 : valid_618; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3727 = state == 3'h7 ? _GEN_2701 : valid_619; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3728 = state == 3'h7 ? _GEN_2702 : valid_620; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3729 = state == 3'h7 ? _GEN_2703 : valid_621; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3730 = state == 3'h7 ? _GEN_2704 : valid_622; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3731 = state == 3'h7 ? _GEN_2705 : valid_623; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3732 = state == 3'h7 ? _GEN_2706 : valid_624; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3733 = state == 3'h7 ? _GEN_2707 : valid_625; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3734 = state == 3'h7 ? _GEN_2708 : valid_626; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3735 = state == 3'h7 ? _GEN_2709 : valid_627; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3736 = state == 3'h7 ? _GEN_2710 : valid_628; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3737 = state == 3'h7 ? _GEN_2711 : valid_629; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3738 = state == 3'h7 ? _GEN_2712 : valid_630; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3739 = state == 3'h7 ? _GEN_2713 : valid_631; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3740 = state == 3'h7 ? _GEN_2714 : valid_632; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3741 = state == 3'h7 ? _GEN_2715 : valid_633; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3742 = state == 3'h7 ? _GEN_2716 : valid_634; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3743 = state == 3'h7 ? _GEN_2717 : valid_635; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3744 = state == 3'h7 ? _GEN_2718 : valid_636; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3745 = state == 3'h7 ? _GEN_2719 : valid_637; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3746 = state == 3'h7 ? _GEN_2720 : valid_638; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3747 = state == 3'h7 ? _GEN_2721 : valid_639; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3748 = state == 3'h7 ? _GEN_2722 : valid_640; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3749 = state == 3'h7 ? _GEN_2723 : valid_641; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3750 = state == 3'h7 ? _GEN_2724 : valid_642; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3751 = state == 3'h7 ? _GEN_2725 : valid_643; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3752 = state == 3'h7 ? _GEN_2726 : valid_644; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3753 = state == 3'h7 ? _GEN_2727 : valid_645; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3754 = state == 3'h7 ? _GEN_2728 : valid_646; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3755 = state == 3'h7 ? _GEN_2729 : valid_647; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3756 = state == 3'h7 ? _GEN_2730 : valid_648; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3757 = state == 3'h7 ? _GEN_2731 : valid_649; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3758 = state == 3'h7 ? _GEN_2732 : valid_650; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3759 = state == 3'h7 ? _GEN_2733 : valid_651; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3760 = state == 3'h7 ? _GEN_2734 : valid_652; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3761 = state == 3'h7 ? _GEN_2735 : valid_653; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3762 = state == 3'h7 ? _GEN_2736 : valid_654; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3763 = state == 3'h7 ? _GEN_2737 : valid_655; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3764 = state == 3'h7 ? _GEN_2738 : valid_656; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3765 = state == 3'h7 ? _GEN_2739 : valid_657; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3766 = state == 3'h7 ? _GEN_2740 : valid_658; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3767 = state == 3'h7 ? _GEN_2741 : valid_659; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3768 = state == 3'h7 ? _GEN_2742 : valid_660; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3769 = state == 3'h7 ? _GEN_2743 : valid_661; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3770 = state == 3'h7 ? _GEN_2744 : valid_662; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3771 = state == 3'h7 ? _GEN_2745 : valid_663; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3772 = state == 3'h7 ? _GEN_2746 : valid_664; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3773 = state == 3'h7 ? _GEN_2747 : valid_665; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3774 = state == 3'h7 ? _GEN_2748 : valid_666; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3775 = state == 3'h7 ? _GEN_2749 : valid_667; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3776 = state == 3'h7 ? _GEN_2750 : valid_668; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3777 = state == 3'h7 ? _GEN_2751 : valid_669; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3778 = state == 3'h7 ? _GEN_2752 : valid_670; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3779 = state == 3'h7 ? _GEN_2753 : valid_671; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3780 = state == 3'h7 ? _GEN_2754 : valid_672; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3781 = state == 3'h7 ? _GEN_2755 : valid_673; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3782 = state == 3'h7 ? _GEN_2756 : valid_674; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3783 = state == 3'h7 ? _GEN_2757 : valid_675; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3784 = state == 3'h7 ? _GEN_2758 : valid_676; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3785 = state == 3'h7 ? _GEN_2759 : valid_677; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3786 = state == 3'h7 ? _GEN_2760 : valid_678; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3787 = state == 3'h7 ? _GEN_2761 : valid_679; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3788 = state == 3'h7 ? _GEN_2762 : valid_680; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3789 = state == 3'h7 ? _GEN_2763 : valid_681; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3790 = state == 3'h7 ? _GEN_2764 : valid_682; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3791 = state == 3'h7 ? _GEN_2765 : valid_683; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3792 = state == 3'h7 ? _GEN_2766 : valid_684; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3793 = state == 3'h7 ? _GEN_2767 : valid_685; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3794 = state == 3'h7 ? _GEN_2768 : valid_686; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3795 = state == 3'h7 ? _GEN_2769 : valid_687; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3796 = state == 3'h7 ? _GEN_2770 : valid_688; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3797 = state == 3'h7 ? _GEN_2771 : valid_689; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3798 = state == 3'h7 ? _GEN_2772 : valid_690; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3799 = state == 3'h7 ? _GEN_2773 : valid_691; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3800 = state == 3'h7 ? _GEN_2774 : valid_692; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3801 = state == 3'h7 ? _GEN_2775 : valid_693; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3802 = state == 3'h7 ? _GEN_2776 : valid_694; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3803 = state == 3'h7 ? _GEN_2777 : valid_695; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3804 = state == 3'h7 ? _GEN_2778 : valid_696; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3805 = state == 3'h7 ? _GEN_2779 : valid_697; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3806 = state == 3'h7 ? _GEN_2780 : valid_698; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3807 = state == 3'h7 ? _GEN_2781 : valid_699; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3808 = state == 3'h7 ? _GEN_2782 : valid_700; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3809 = state == 3'h7 ? _GEN_2783 : valid_701; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3810 = state == 3'h7 ? _GEN_2784 : valid_702; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3811 = state == 3'h7 ? _GEN_2785 : valid_703; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3812 = state == 3'h7 ? _GEN_2786 : valid_704; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3813 = state == 3'h7 ? _GEN_2787 : valid_705; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3814 = state == 3'h7 ? _GEN_2788 : valid_706; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3815 = state == 3'h7 ? _GEN_2789 : valid_707; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3816 = state == 3'h7 ? _GEN_2790 : valid_708; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3817 = state == 3'h7 ? _GEN_2791 : valid_709; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3818 = state == 3'h7 ? _GEN_2792 : valid_710; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3819 = state == 3'h7 ? _GEN_2793 : valid_711; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3820 = state == 3'h7 ? _GEN_2794 : valid_712; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3821 = state == 3'h7 ? _GEN_2795 : valid_713; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3822 = state == 3'h7 ? _GEN_2796 : valid_714; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3823 = state == 3'h7 ? _GEN_2797 : valid_715; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3824 = state == 3'h7 ? _GEN_2798 : valid_716; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3825 = state == 3'h7 ? _GEN_2799 : valid_717; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3826 = state == 3'h7 ? _GEN_2800 : valid_718; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3827 = state == 3'h7 ? _GEN_2801 : valid_719; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3828 = state == 3'h7 ? _GEN_2802 : valid_720; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3829 = state == 3'h7 ? _GEN_2803 : valid_721; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3830 = state == 3'h7 ? _GEN_2804 : valid_722; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3831 = state == 3'h7 ? _GEN_2805 : valid_723; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3832 = state == 3'h7 ? _GEN_2806 : valid_724; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3833 = state == 3'h7 ? _GEN_2807 : valid_725; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3834 = state == 3'h7 ? _GEN_2808 : valid_726; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3835 = state == 3'h7 ? _GEN_2809 : valid_727; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3836 = state == 3'h7 ? _GEN_2810 : valid_728; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3837 = state == 3'h7 ? _GEN_2811 : valid_729; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3838 = state == 3'h7 ? _GEN_2812 : valid_730; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3839 = state == 3'h7 ? _GEN_2813 : valid_731; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3840 = state == 3'h7 ? _GEN_2814 : valid_732; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3841 = state == 3'h7 ? _GEN_2815 : valid_733; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3842 = state == 3'h7 ? _GEN_2816 : valid_734; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3843 = state == 3'h7 ? _GEN_2817 : valid_735; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3844 = state == 3'h7 ? _GEN_2818 : valid_736; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3845 = state == 3'h7 ? _GEN_2819 : valid_737; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3846 = state == 3'h7 ? _GEN_2820 : valid_738; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3847 = state == 3'h7 ? _GEN_2821 : valid_739; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3848 = state == 3'h7 ? _GEN_2822 : valid_740; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3849 = state == 3'h7 ? _GEN_2823 : valid_741; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3850 = state == 3'h7 ? _GEN_2824 : valid_742; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3851 = state == 3'h7 ? _GEN_2825 : valid_743; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3852 = state == 3'h7 ? _GEN_2826 : valid_744; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3853 = state == 3'h7 ? _GEN_2827 : valid_745; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3854 = state == 3'h7 ? _GEN_2828 : valid_746; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3855 = state == 3'h7 ? _GEN_2829 : valid_747; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3856 = state == 3'h7 ? _GEN_2830 : valid_748; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3857 = state == 3'h7 ? _GEN_2831 : valid_749; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3858 = state == 3'h7 ? _GEN_2832 : valid_750; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3859 = state == 3'h7 ? _GEN_2833 : valid_751; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3860 = state == 3'h7 ? _GEN_2834 : valid_752; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3861 = state == 3'h7 ? _GEN_2835 : valid_753; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3862 = state == 3'h7 ? _GEN_2836 : valid_754; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3863 = state == 3'h7 ? _GEN_2837 : valid_755; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3864 = state == 3'h7 ? _GEN_2838 : valid_756; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3865 = state == 3'h7 ? _GEN_2839 : valid_757; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3866 = state == 3'h7 ? _GEN_2840 : valid_758; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3867 = state == 3'h7 ? _GEN_2841 : valid_759; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3868 = state == 3'h7 ? _GEN_2842 : valid_760; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3869 = state == 3'h7 ? _GEN_2843 : valid_761; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3870 = state == 3'h7 ? _GEN_2844 : valid_762; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3871 = state == 3'h7 ? _GEN_2845 : valid_763; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3872 = state == 3'h7 ? _GEN_2846 : valid_764; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3873 = state == 3'h7 ? _GEN_2847 : valid_765; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3874 = state == 3'h7 ? _GEN_2848 : valid_766; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3875 = state == 3'h7 ? _GEN_2849 : valid_767; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3876 = state == 3'h7 ? _GEN_2850 : valid_768; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3877 = state == 3'h7 ? _GEN_2851 : valid_769; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3878 = state == 3'h7 ? _GEN_2852 : valid_770; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3879 = state == 3'h7 ? _GEN_2853 : valid_771; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3880 = state == 3'h7 ? _GEN_2854 : valid_772; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3881 = state == 3'h7 ? _GEN_2855 : valid_773; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3882 = state == 3'h7 ? _GEN_2856 : valid_774; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3883 = state == 3'h7 ? _GEN_2857 : valid_775; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3884 = state == 3'h7 ? _GEN_2858 : valid_776; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3885 = state == 3'h7 ? _GEN_2859 : valid_777; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3886 = state == 3'h7 ? _GEN_2860 : valid_778; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3887 = state == 3'h7 ? _GEN_2861 : valid_779; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3888 = state == 3'h7 ? _GEN_2862 : valid_780; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3889 = state == 3'h7 ? _GEN_2863 : valid_781; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3890 = state == 3'h7 ? _GEN_2864 : valid_782; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3891 = state == 3'h7 ? _GEN_2865 : valid_783; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3892 = state == 3'h7 ? _GEN_2866 : valid_784; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3893 = state == 3'h7 ? _GEN_2867 : valid_785; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3894 = state == 3'h7 ? _GEN_2868 : valid_786; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3895 = state == 3'h7 ? _GEN_2869 : valid_787; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3896 = state == 3'h7 ? _GEN_2870 : valid_788; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3897 = state == 3'h7 ? _GEN_2871 : valid_789; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3898 = state == 3'h7 ? _GEN_2872 : valid_790; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3899 = state == 3'h7 ? _GEN_2873 : valid_791; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3900 = state == 3'h7 ? _GEN_2874 : valid_792; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3901 = state == 3'h7 ? _GEN_2875 : valid_793; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3902 = state == 3'h7 ? _GEN_2876 : valid_794; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3903 = state == 3'h7 ? _GEN_2877 : valid_795; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3904 = state == 3'h7 ? _GEN_2878 : valid_796; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3905 = state == 3'h7 ? _GEN_2879 : valid_797; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3906 = state == 3'h7 ? _GEN_2880 : valid_798; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3907 = state == 3'h7 ? _GEN_2881 : valid_799; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3908 = state == 3'h7 ? _GEN_2882 : valid_800; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3909 = state == 3'h7 ? _GEN_2883 : valid_801; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3910 = state == 3'h7 ? _GEN_2884 : valid_802; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3911 = state == 3'h7 ? _GEN_2885 : valid_803; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3912 = state == 3'h7 ? _GEN_2886 : valid_804; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3913 = state == 3'h7 ? _GEN_2887 : valid_805; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3914 = state == 3'h7 ? _GEN_2888 : valid_806; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3915 = state == 3'h7 ? _GEN_2889 : valid_807; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3916 = state == 3'h7 ? _GEN_2890 : valid_808; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3917 = state == 3'h7 ? _GEN_2891 : valid_809; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3918 = state == 3'h7 ? _GEN_2892 : valid_810; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3919 = state == 3'h7 ? _GEN_2893 : valid_811; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3920 = state == 3'h7 ? _GEN_2894 : valid_812; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3921 = state == 3'h7 ? _GEN_2895 : valid_813; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3922 = state == 3'h7 ? _GEN_2896 : valid_814; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3923 = state == 3'h7 ? _GEN_2897 : valid_815; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3924 = state == 3'h7 ? _GEN_2898 : valid_816; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3925 = state == 3'h7 ? _GEN_2899 : valid_817; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3926 = state == 3'h7 ? _GEN_2900 : valid_818; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3927 = state == 3'h7 ? _GEN_2901 : valid_819; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3928 = state == 3'h7 ? _GEN_2902 : valid_820; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3929 = state == 3'h7 ? _GEN_2903 : valid_821; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3930 = state == 3'h7 ? _GEN_2904 : valid_822; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3931 = state == 3'h7 ? _GEN_2905 : valid_823; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3932 = state == 3'h7 ? _GEN_2906 : valid_824; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3933 = state == 3'h7 ? _GEN_2907 : valid_825; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3934 = state == 3'h7 ? _GEN_2908 : valid_826; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3935 = state == 3'h7 ? _GEN_2909 : valid_827; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3936 = state == 3'h7 ? _GEN_2910 : valid_828; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3937 = state == 3'h7 ? _GEN_2911 : valid_829; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3938 = state == 3'h7 ? _GEN_2912 : valid_830; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3939 = state == 3'h7 ? _GEN_2913 : valid_831; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3940 = state == 3'h7 ? _GEN_2914 : valid_832; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3941 = state == 3'h7 ? _GEN_2915 : valid_833; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3942 = state == 3'h7 ? _GEN_2916 : valid_834; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3943 = state == 3'h7 ? _GEN_2917 : valid_835; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3944 = state == 3'h7 ? _GEN_2918 : valid_836; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3945 = state == 3'h7 ? _GEN_2919 : valid_837; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3946 = state == 3'h7 ? _GEN_2920 : valid_838; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3947 = state == 3'h7 ? _GEN_2921 : valid_839; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3948 = state == 3'h7 ? _GEN_2922 : valid_840; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3949 = state == 3'h7 ? _GEN_2923 : valid_841; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3950 = state == 3'h7 ? _GEN_2924 : valid_842; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3951 = state == 3'h7 ? _GEN_2925 : valid_843; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3952 = state == 3'h7 ? _GEN_2926 : valid_844; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3953 = state == 3'h7 ? _GEN_2927 : valid_845; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3954 = state == 3'h7 ? _GEN_2928 : valid_846; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3955 = state == 3'h7 ? _GEN_2929 : valid_847; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3956 = state == 3'h7 ? _GEN_2930 : valid_848; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3957 = state == 3'h7 ? _GEN_2931 : valid_849; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3958 = state == 3'h7 ? _GEN_2932 : valid_850; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3959 = state == 3'h7 ? _GEN_2933 : valid_851; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3960 = state == 3'h7 ? _GEN_2934 : valid_852; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3961 = state == 3'h7 ? _GEN_2935 : valid_853; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3962 = state == 3'h7 ? _GEN_2936 : valid_854; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3963 = state == 3'h7 ? _GEN_2937 : valid_855; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3964 = state == 3'h7 ? _GEN_2938 : valid_856; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3965 = state == 3'h7 ? _GEN_2939 : valid_857; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3966 = state == 3'h7 ? _GEN_2940 : valid_858; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3967 = state == 3'h7 ? _GEN_2941 : valid_859; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3968 = state == 3'h7 ? _GEN_2942 : valid_860; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3969 = state == 3'h7 ? _GEN_2943 : valid_861; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3970 = state == 3'h7 ? _GEN_2944 : valid_862; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3971 = state == 3'h7 ? _GEN_2945 : valid_863; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3972 = state == 3'h7 ? _GEN_2946 : valid_864; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3973 = state == 3'h7 ? _GEN_2947 : valid_865; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3974 = state == 3'h7 ? _GEN_2948 : valid_866; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3975 = state == 3'h7 ? _GEN_2949 : valid_867; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3976 = state == 3'h7 ? _GEN_2950 : valid_868; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3977 = state == 3'h7 ? _GEN_2951 : valid_869; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3978 = state == 3'h7 ? _GEN_2952 : valid_870; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3979 = state == 3'h7 ? _GEN_2953 : valid_871; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3980 = state == 3'h7 ? _GEN_2954 : valid_872; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3981 = state == 3'h7 ? _GEN_2955 : valid_873; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3982 = state == 3'h7 ? _GEN_2956 : valid_874; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3983 = state == 3'h7 ? _GEN_2957 : valid_875; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3984 = state == 3'h7 ? _GEN_2958 : valid_876; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3985 = state == 3'h7 ? _GEN_2959 : valid_877; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3986 = state == 3'h7 ? _GEN_2960 : valid_878; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3987 = state == 3'h7 ? _GEN_2961 : valid_879; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3988 = state == 3'h7 ? _GEN_2962 : valid_880; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3989 = state == 3'h7 ? _GEN_2963 : valid_881; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3990 = state == 3'h7 ? _GEN_2964 : valid_882; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3991 = state == 3'h7 ? _GEN_2965 : valid_883; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3992 = state == 3'h7 ? _GEN_2966 : valid_884; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3993 = state == 3'h7 ? _GEN_2967 : valid_885; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3994 = state == 3'h7 ? _GEN_2968 : valid_886; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3995 = state == 3'h7 ? _GEN_2969 : valid_887; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3996 = state == 3'h7 ? _GEN_2970 : valid_888; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3997 = state == 3'h7 ? _GEN_2971 : valid_889; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3998 = state == 3'h7 ? _GEN_2972 : valid_890; // @[DCache.scala 165:26 56:22]
  wire  _GEN_3999 = state == 3'h7 ? _GEN_2973 : valid_891; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4000 = state == 3'h7 ? _GEN_2974 : valid_892; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4001 = state == 3'h7 ? _GEN_2975 : valid_893; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4002 = state == 3'h7 ? _GEN_2976 : valid_894; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4003 = state == 3'h7 ? _GEN_2977 : valid_895; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4004 = state == 3'h7 ? _GEN_2978 : valid_896; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4005 = state == 3'h7 ? _GEN_2979 : valid_897; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4006 = state == 3'h7 ? _GEN_2980 : valid_898; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4007 = state == 3'h7 ? _GEN_2981 : valid_899; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4008 = state == 3'h7 ? _GEN_2982 : valid_900; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4009 = state == 3'h7 ? _GEN_2983 : valid_901; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4010 = state == 3'h7 ? _GEN_2984 : valid_902; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4011 = state == 3'h7 ? _GEN_2985 : valid_903; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4012 = state == 3'h7 ? _GEN_2986 : valid_904; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4013 = state == 3'h7 ? _GEN_2987 : valid_905; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4014 = state == 3'h7 ? _GEN_2988 : valid_906; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4015 = state == 3'h7 ? _GEN_2989 : valid_907; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4016 = state == 3'h7 ? _GEN_2990 : valid_908; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4017 = state == 3'h7 ? _GEN_2991 : valid_909; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4018 = state == 3'h7 ? _GEN_2992 : valid_910; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4019 = state == 3'h7 ? _GEN_2993 : valid_911; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4020 = state == 3'h7 ? _GEN_2994 : valid_912; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4021 = state == 3'h7 ? _GEN_2995 : valid_913; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4022 = state == 3'h7 ? _GEN_2996 : valid_914; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4023 = state == 3'h7 ? _GEN_2997 : valid_915; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4024 = state == 3'h7 ? _GEN_2998 : valid_916; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4025 = state == 3'h7 ? _GEN_2999 : valid_917; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4026 = state == 3'h7 ? _GEN_3000 : valid_918; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4027 = state == 3'h7 ? _GEN_3001 : valid_919; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4028 = state == 3'h7 ? _GEN_3002 : valid_920; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4029 = state == 3'h7 ? _GEN_3003 : valid_921; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4030 = state == 3'h7 ? _GEN_3004 : valid_922; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4031 = state == 3'h7 ? _GEN_3005 : valid_923; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4032 = state == 3'h7 ? _GEN_3006 : valid_924; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4033 = state == 3'h7 ? _GEN_3007 : valid_925; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4034 = state == 3'h7 ? _GEN_3008 : valid_926; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4035 = state == 3'h7 ? _GEN_3009 : valid_927; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4036 = state == 3'h7 ? _GEN_3010 : valid_928; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4037 = state == 3'h7 ? _GEN_3011 : valid_929; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4038 = state == 3'h7 ? _GEN_3012 : valid_930; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4039 = state == 3'h7 ? _GEN_3013 : valid_931; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4040 = state == 3'h7 ? _GEN_3014 : valid_932; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4041 = state == 3'h7 ? _GEN_3015 : valid_933; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4042 = state == 3'h7 ? _GEN_3016 : valid_934; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4043 = state == 3'h7 ? _GEN_3017 : valid_935; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4044 = state == 3'h7 ? _GEN_3018 : valid_936; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4045 = state == 3'h7 ? _GEN_3019 : valid_937; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4046 = state == 3'h7 ? _GEN_3020 : valid_938; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4047 = state == 3'h7 ? _GEN_3021 : valid_939; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4048 = state == 3'h7 ? _GEN_3022 : valid_940; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4049 = state == 3'h7 ? _GEN_3023 : valid_941; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4050 = state == 3'h7 ? _GEN_3024 : valid_942; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4051 = state == 3'h7 ? _GEN_3025 : valid_943; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4052 = state == 3'h7 ? _GEN_3026 : valid_944; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4053 = state == 3'h7 ? _GEN_3027 : valid_945; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4054 = state == 3'h7 ? _GEN_3028 : valid_946; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4055 = state == 3'h7 ? _GEN_3029 : valid_947; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4056 = state == 3'h7 ? _GEN_3030 : valid_948; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4057 = state == 3'h7 ? _GEN_3031 : valid_949; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4058 = state == 3'h7 ? _GEN_3032 : valid_950; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4059 = state == 3'h7 ? _GEN_3033 : valid_951; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4060 = state == 3'h7 ? _GEN_3034 : valid_952; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4061 = state == 3'h7 ? _GEN_3035 : valid_953; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4062 = state == 3'h7 ? _GEN_3036 : valid_954; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4063 = state == 3'h7 ? _GEN_3037 : valid_955; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4064 = state == 3'h7 ? _GEN_3038 : valid_956; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4065 = state == 3'h7 ? _GEN_3039 : valid_957; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4066 = state == 3'h7 ? _GEN_3040 : valid_958; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4067 = state == 3'h7 ? _GEN_3041 : valid_959; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4068 = state == 3'h7 ? _GEN_3042 : valid_960; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4069 = state == 3'h7 ? _GEN_3043 : valid_961; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4070 = state == 3'h7 ? _GEN_3044 : valid_962; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4071 = state == 3'h7 ? _GEN_3045 : valid_963; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4072 = state == 3'h7 ? _GEN_3046 : valid_964; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4073 = state == 3'h7 ? _GEN_3047 : valid_965; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4074 = state == 3'h7 ? _GEN_3048 : valid_966; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4075 = state == 3'h7 ? _GEN_3049 : valid_967; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4076 = state == 3'h7 ? _GEN_3050 : valid_968; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4077 = state == 3'h7 ? _GEN_3051 : valid_969; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4078 = state == 3'h7 ? _GEN_3052 : valid_970; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4079 = state == 3'h7 ? _GEN_3053 : valid_971; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4080 = state == 3'h7 ? _GEN_3054 : valid_972; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4081 = state == 3'h7 ? _GEN_3055 : valid_973; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4082 = state == 3'h7 ? _GEN_3056 : valid_974; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4083 = state == 3'h7 ? _GEN_3057 : valid_975; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4084 = state == 3'h7 ? _GEN_3058 : valid_976; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4085 = state == 3'h7 ? _GEN_3059 : valid_977; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4086 = state == 3'h7 ? _GEN_3060 : valid_978; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4087 = state == 3'h7 ? _GEN_3061 : valid_979; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4088 = state == 3'h7 ? _GEN_3062 : valid_980; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4089 = state == 3'h7 ? _GEN_3063 : valid_981; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4090 = state == 3'h7 ? _GEN_3064 : valid_982; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4091 = state == 3'h7 ? _GEN_3065 : valid_983; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4092 = state == 3'h7 ? _GEN_3066 : valid_984; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4093 = state == 3'h7 ? _GEN_3067 : valid_985; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4094 = state == 3'h7 ? _GEN_3068 : valid_986; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4095 = state == 3'h7 ? _GEN_3069 : valid_987; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4096 = state == 3'h7 ? _GEN_3070 : valid_988; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4097 = state == 3'h7 ? _GEN_3071 : valid_989; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4098 = state == 3'h7 ? _GEN_3072 : valid_990; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4099 = state == 3'h7 ? _GEN_3073 : valid_991; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4100 = state == 3'h7 ? _GEN_3074 : valid_992; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4101 = state == 3'h7 ? _GEN_3075 : valid_993; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4102 = state == 3'h7 ? _GEN_3076 : valid_994; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4103 = state == 3'h7 ? _GEN_3077 : valid_995; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4104 = state == 3'h7 ? _GEN_3078 : valid_996; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4105 = state == 3'h7 ? _GEN_3079 : valid_997; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4106 = state == 3'h7 ? _GEN_3080 : valid_998; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4107 = state == 3'h7 ? _GEN_3081 : valid_999; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4108 = state == 3'h7 ? _GEN_3082 : valid_1000; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4109 = state == 3'h7 ? _GEN_3083 : valid_1001; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4110 = state == 3'h7 ? _GEN_3084 : valid_1002; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4111 = state == 3'h7 ? _GEN_3085 : valid_1003; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4112 = state == 3'h7 ? _GEN_3086 : valid_1004; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4113 = state == 3'h7 ? _GEN_3087 : valid_1005; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4114 = state == 3'h7 ? _GEN_3088 : valid_1006; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4115 = state == 3'h7 ? _GEN_3089 : valid_1007; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4116 = state == 3'h7 ? _GEN_3090 : valid_1008; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4117 = state == 3'h7 ? _GEN_3091 : valid_1009; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4118 = state == 3'h7 ? _GEN_3092 : valid_1010; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4119 = state == 3'h7 ? _GEN_3093 : valid_1011; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4120 = state == 3'h7 ? _GEN_3094 : valid_1012; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4121 = state == 3'h7 ? _GEN_3095 : valid_1013; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4122 = state == 3'h7 ? _GEN_3096 : valid_1014; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4123 = state == 3'h7 ? _GEN_3097 : valid_1015; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4124 = state == 3'h7 ? _GEN_3098 : valid_1016; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4125 = state == 3'h7 ? _GEN_3099 : valid_1017; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4126 = state == 3'h7 ? _GEN_3100 : valid_1018; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4127 = state == 3'h7 ? _GEN_3101 : valid_1019; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4128 = state == 3'h7 ? _GEN_3102 : valid_1020; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4129 = state == 3'h7 ? _GEN_3103 : valid_1021; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4130 = state == 3'h7 ? _GEN_3104 : valid_1022; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4131 = state == 3'h7 ? _GEN_3105 : valid_1023; // @[DCache.scala 165:26 56:22]
  wire  _GEN_4134 = _array_io_en_T_1 ? _GEN_3108 : valid_0; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4135 = _array_io_en_T_1 ? _GEN_3109 : valid_1; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4136 = _array_io_en_T_1 ? _GEN_3110 : valid_2; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4137 = _array_io_en_T_1 ? _GEN_3111 : valid_3; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4138 = _array_io_en_T_1 ? _GEN_3112 : valid_4; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4139 = _array_io_en_T_1 ? _GEN_3113 : valid_5; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4140 = _array_io_en_T_1 ? _GEN_3114 : valid_6; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4141 = _array_io_en_T_1 ? _GEN_3115 : valid_7; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4142 = _array_io_en_T_1 ? _GEN_3116 : valid_8; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4143 = _array_io_en_T_1 ? _GEN_3117 : valid_9; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4144 = _array_io_en_T_1 ? _GEN_3118 : valid_10; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4145 = _array_io_en_T_1 ? _GEN_3119 : valid_11; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4146 = _array_io_en_T_1 ? _GEN_3120 : valid_12; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4147 = _array_io_en_T_1 ? _GEN_3121 : valid_13; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4148 = _array_io_en_T_1 ? _GEN_3122 : valid_14; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4149 = _array_io_en_T_1 ? _GEN_3123 : valid_15; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4150 = _array_io_en_T_1 ? _GEN_3124 : valid_16; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4151 = _array_io_en_T_1 ? _GEN_3125 : valid_17; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4152 = _array_io_en_T_1 ? _GEN_3126 : valid_18; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4153 = _array_io_en_T_1 ? _GEN_3127 : valid_19; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4154 = _array_io_en_T_1 ? _GEN_3128 : valid_20; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4155 = _array_io_en_T_1 ? _GEN_3129 : valid_21; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4156 = _array_io_en_T_1 ? _GEN_3130 : valid_22; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4157 = _array_io_en_T_1 ? _GEN_3131 : valid_23; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4158 = _array_io_en_T_1 ? _GEN_3132 : valid_24; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4159 = _array_io_en_T_1 ? _GEN_3133 : valid_25; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4160 = _array_io_en_T_1 ? _GEN_3134 : valid_26; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4161 = _array_io_en_T_1 ? _GEN_3135 : valid_27; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4162 = _array_io_en_T_1 ? _GEN_3136 : valid_28; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4163 = _array_io_en_T_1 ? _GEN_3137 : valid_29; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4164 = _array_io_en_T_1 ? _GEN_3138 : valid_30; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4165 = _array_io_en_T_1 ? _GEN_3139 : valid_31; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4166 = _array_io_en_T_1 ? _GEN_3140 : valid_32; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4167 = _array_io_en_T_1 ? _GEN_3141 : valid_33; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4168 = _array_io_en_T_1 ? _GEN_3142 : valid_34; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4169 = _array_io_en_T_1 ? _GEN_3143 : valid_35; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4170 = _array_io_en_T_1 ? _GEN_3144 : valid_36; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4171 = _array_io_en_T_1 ? _GEN_3145 : valid_37; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4172 = _array_io_en_T_1 ? _GEN_3146 : valid_38; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4173 = _array_io_en_T_1 ? _GEN_3147 : valid_39; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4174 = _array_io_en_T_1 ? _GEN_3148 : valid_40; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4175 = _array_io_en_T_1 ? _GEN_3149 : valid_41; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4176 = _array_io_en_T_1 ? _GEN_3150 : valid_42; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4177 = _array_io_en_T_1 ? _GEN_3151 : valid_43; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4178 = _array_io_en_T_1 ? _GEN_3152 : valid_44; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4179 = _array_io_en_T_1 ? _GEN_3153 : valid_45; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4180 = _array_io_en_T_1 ? _GEN_3154 : valid_46; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4181 = _array_io_en_T_1 ? _GEN_3155 : valid_47; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4182 = _array_io_en_T_1 ? _GEN_3156 : valid_48; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4183 = _array_io_en_T_1 ? _GEN_3157 : valid_49; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4184 = _array_io_en_T_1 ? _GEN_3158 : valid_50; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4185 = _array_io_en_T_1 ? _GEN_3159 : valid_51; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4186 = _array_io_en_T_1 ? _GEN_3160 : valid_52; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4187 = _array_io_en_T_1 ? _GEN_3161 : valid_53; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4188 = _array_io_en_T_1 ? _GEN_3162 : valid_54; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4189 = _array_io_en_T_1 ? _GEN_3163 : valid_55; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4190 = _array_io_en_T_1 ? _GEN_3164 : valid_56; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4191 = _array_io_en_T_1 ? _GEN_3165 : valid_57; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4192 = _array_io_en_T_1 ? _GEN_3166 : valid_58; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4193 = _array_io_en_T_1 ? _GEN_3167 : valid_59; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4194 = _array_io_en_T_1 ? _GEN_3168 : valid_60; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4195 = _array_io_en_T_1 ? _GEN_3169 : valid_61; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4196 = _array_io_en_T_1 ? _GEN_3170 : valid_62; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4197 = _array_io_en_T_1 ? _GEN_3171 : valid_63; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4198 = _array_io_en_T_1 ? _GEN_3172 : valid_64; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4199 = _array_io_en_T_1 ? _GEN_3173 : valid_65; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4200 = _array_io_en_T_1 ? _GEN_3174 : valid_66; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4201 = _array_io_en_T_1 ? _GEN_3175 : valid_67; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4202 = _array_io_en_T_1 ? _GEN_3176 : valid_68; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4203 = _array_io_en_T_1 ? _GEN_3177 : valid_69; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4204 = _array_io_en_T_1 ? _GEN_3178 : valid_70; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4205 = _array_io_en_T_1 ? _GEN_3179 : valid_71; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4206 = _array_io_en_T_1 ? _GEN_3180 : valid_72; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4207 = _array_io_en_T_1 ? _GEN_3181 : valid_73; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4208 = _array_io_en_T_1 ? _GEN_3182 : valid_74; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4209 = _array_io_en_T_1 ? _GEN_3183 : valid_75; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4210 = _array_io_en_T_1 ? _GEN_3184 : valid_76; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4211 = _array_io_en_T_1 ? _GEN_3185 : valid_77; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4212 = _array_io_en_T_1 ? _GEN_3186 : valid_78; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4213 = _array_io_en_T_1 ? _GEN_3187 : valid_79; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4214 = _array_io_en_T_1 ? _GEN_3188 : valid_80; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4215 = _array_io_en_T_1 ? _GEN_3189 : valid_81; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4216 = _array_io_en_T_1 ? _GEN_3190 : valid_82; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4217 = _array_io_en_T_1 ? _GEN_3191 : valid_83; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4218 = _array_io_en_T_1 ? _GEN_3192 : valid_84; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4219 = _array_io_en_T_1 ? _GEN_3193 : valid_85; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4220 = _array_io_en_T_1 ? _GEN_3194 : valid_86; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4221 = _array_io_en_T_1 ? _GEN_3195 : valid_87; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4222 = _array_io_en_T_1 ? _GEN_3196 : valid_88; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4223 = _array_io_en_T_1 ? _GEN_3197 : valid_89; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4224 = _array_io_en_T_1 ? _GEN_3198 : valid_90; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4225 = _array_io_en_T_1 ? _GEN_3199 : valid_91; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4226 = _array_io_en_T_1 ? _GEN_3200 : valid_92; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4227 = _array_io_en_T_1 ? _GEN_3201 : valid_93; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4228 = _array_io_en_T_1 ? _GEN_3202 : valid_94; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4229 = _array_io_en_T_1 ? _GEN_3203 : valid_95; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4230 = _array_io_en_T_1 ? _GEN_3204 : valid_96; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4231 = _array_io_en_T_1 ? _GEN_3205 : valid_97; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4232 = _array_io_en_T_1 ? _GEN_3206 : valid_98; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4233 = _array_io_en_T_1 ? _GEN_3207 : valid_99; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4234 = _array_io_en_T_1 ? _GEN_3208 : valid_100; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4235 = _array_io_en_T_1 ? _GEN_3209 : valid_101; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4236 = _array_io_en_T_1 ? _GEN_3210 : valid_102; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4237 = _array_io_en_T_1 ? _GEN_3211 : valid_103; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4238 = _array_io_en_T_1 ? _GEN_3212 : valid_104; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4239 = _array_io_en_T_1 ? _GEN_3213 : valid_105; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4240 = _array_io_en_T_1 ? _GEN_3214 : valid_106; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4241 = _array_io_en_T_1 ? _GEN_3215 : valid_107; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4242 = _array_io_en_T_1 ? _GEN_3216 : valid_108; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4243 = _array_io_en_T_1 ? _GEN_3217 : valid_109; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4244 = _array_io_en_T_1 ? _GEN_3218 : valid_110; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4245 = _array_io_en_T_1 ? _GEN_3219 : valid_111; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4246 = _array_io_en_T_1 ? _GEN_3220 : valid_112; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4247 = _array_io_en_T_1 ? _GEN_3221 : valid_113; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4248 = _array_io_en_T_1 ? _GEN_3222 : valid_114; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4249 = _array_io_en_T_1 ? _GEN_3223 : valid_115; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4250 = _array_io_en_T_1 ? _GEN_3224 : valid_116; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4251 = _array_io_en_T_1 ? _GEN_3225 : valid_117; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4252 = _array_io_en_T_1 ? _GEN_3226 : valid_118; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4253 = _array_io_en_T_1 ? _GEN_3227 : valid_119; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4254 = _array_io_en_T_1 ? _GEN_3228 : valid_120; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4255 = _array_io_en_T_1 ? _GEN_3229 : valid_121; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4256 = _array_io_en_T_1 ? _GEN_3230 : valid_122; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4257 = _array_io_en_T_1 ? _GEN_3231 : valid_123; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4258 = _array_io_en_T_1 ? _GEN_3232 : valid_124; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4259 = _array_io_en_T_1 ? _GEN_3233 : valid_125; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4260 = _array_io_en_T_1 ? _GEN_3234 : valid_126; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4261 = _array_io_en_T_1 ? _GEN_3235 : valid_127; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4262 = _array_io_en_T_1 ? _GEN_3236 : valid_128; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4263 = _array_io_en_T_1 ? _GEN_3237 : valid_129; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4264 = _array_io_en_T_1 ? _GEN_3238 : valid_130; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4265 = _array_io_en_T_1 ? _GEN_3239 : valid_131; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4266 = _array_io_en_T_1 ? _GEN_3240 : valid_132; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4267 = _array_io_en_T_1 ? _GEN_3241 : valid_133; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4268 = _array_io_en_T_1 ? _GEN_3242 : valid_134; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4269 = _array_io_en_T_1 ? _GEN_3243 : valid_135; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4270 = _array_io_en_T_1 ? _GEN_3244 : valid_136; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4271 = _array_io_en_T_1 ? _GEN_3245 : valid_137; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4272 = _array_io_en_T_1 ? _GEN_3246 : valid_138; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4273 = _array_io_en_T_1 ? _GEN_3247 : valid_139; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4274 = _array_io_en_T_1 ? _GEN_3248 : valid_140; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4275 = _array_io_en_T_1 ? _GEN_3249 : valid_141; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4276 = _array_io_en_T_1 ? _GEN_3250 : valid_142; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4277 = _array_io_en_T_1 ? _GEN_3251 : valid_143; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4278 = _array_io_en_T_1 ? _GEN_3252 : valid_144; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4279 = _array_io_en_T_1 ? _GEN_3253 : valid_145; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4280 = _array_io_en_T_1 ? _GEN_3254 : valid_146; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4281 = _array_io_en_T_1 ? _GEN_3255 : valid_147; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4282 = _array_io_en_T_1 ? _GEN_3256 : valid_148; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4283 = _array_io_en_T_1 ? _GEN_3257 : valid_149; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4284 = _array_io_en_T_1 ? _GEN_3258 : valid_150; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4285 = _array_io_en_T_1 ? _GEN_3259 : valid_151; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4286 = _array_io_en_T_1 ? _GEN_3260 : valid_152; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4287 = _array_io_en_T_1 ? _GEN_3261 : valid_153; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4288 = _array_io_en_T_1 ? _GEN_3262 : valid_154; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4289 = _array_io_en_T_1 ? _GEN_3263 : valid_155; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4290 = _array_io_en_T_1 ? _GEN_3264 : valid_156; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4291 = _array_io_en_T_1 ? _GEN_3265 : valid_157; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4292 = _array_io_en_T_1 ? _GEN_3266 : valid_158; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4293 = _array_io_en_T_1 ? _GEN_3267 : valid_159; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4294 = _array_io_en_T_1 ? _GEN_3268 : valid_160; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4295 = _array_io_en_T_1 ? _GEN_3269 : valid_161; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4296 = _array_io_en_T_1 ? _GEN_3270 : valid_162; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4297 = _array_io_en_T_1 ? _GEN_3271 : valid_163; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4298 = _array_io_en_T_1 ? _GEN_3272 : valid_164; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4299 = _array_io_en_T_1 ? _GEN_3273 : valid_165; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4300 = _array_io_en_T_1 ? _GEN_3274 : valid_166; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4301 = _array_io_en_T_1 ? _GEN_3275 : valid_167; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4302 = _array_io_en_T_1 ? _GEN_3276 : valid_168; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4303 = _array_io_en_T_1 ? _GEN_3277 : valid_169; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4304 = _array_io_en_T_1 ? _GEN_3278 : valid_170; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4305 = _array_io_en_T_1 ? _GEN_3279 : valid_171; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4306 = _array_io_en_T_1 ? _GEN_3280 : valid_172; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4307 = _array_io_en_T_1 ? _GEN_3281 : valid_173; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4308 = _array_io_en_T_1 ? _GEN_3282 : valid_174; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4309 = _array_io_en_T_1 ? _GEN_3283 : valid_175; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4310 = _array_io_en_T_1 ? _GEN_3284 : valid_176; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4311 = _array_io_en_T_1 ? _GEN_3285 : valid_177; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4312 = _array_io_en_T_1 ? _GEN_3286 : valid_178; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4313 = _array_io_en_T_1 ? _GEN_3287 : valid_179; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4314 = _array_io_en_T_1 ? _GEN_3288 : valid_180; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4315 = _array_io_en_T_1 ? _GEN_3289 : valid_181; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4316 = _array_io_en_T_1 ? _GEN_3290 : valid_182; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4317 = _array_io_en_T_1 ? _GEN_3291 : valid_183; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4318 = _array_io_en_T_1 ? _GEN_3292 : valid_184; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4319 = _array_io_en_T_1 ? _GEN_3293 : valid_185; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4320 = _array_io_en_T_1 ? _GEN_3294 : valid_186; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4321 = _array_io_en_T_1 ? _GEN_3295 : valid_187; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4322 = _array_io_en_T_1 ? _GEN_3296 : valid_188; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4323 = _array_io_en_T_1 ? _GEN_3297 : valid_189; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4324 = _array_io_en_T_1 ? _GEN_3298 : valid_190; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4325 = _array_io_en_T_1 ? _GEN_3299 : valid_191; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4326 = _array_io_en_T_1 ? _GEN_3300 : valid_192; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4327 = _array_io_en_T_1 ? _GEN_3301 : valid_193; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4328 = _array_io_en_T_1 ? _GEN_3302 : valid_194; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4329 = _array_io_en_T_1 ? _GEN_3303 : valid_195; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4330 = _array_io_en_T_1 ? _GEN_3304 : valid_196; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4331 = _array_io_en_T_1 ? _GEN_3305 : valid_197; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4332 = _array_io_en_T_1 ? _GEN_3306 : valid_198; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4333 = _array_io_en_T_1 ? _GEN_3307 : valid_199; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4334 = _array_io_en_T_1 ? _GEN_3308 : valid_200; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4335 = _array_io_en_T_1 ? _GEN_3309 : valid_201; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4336 = _array_io_en_T_1 ? _GEN_3310 : valid_202; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4337 = _array_io_en_T_1 ? _GEN_3311 : valid_203; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4338 = _array_io_en_T_1 ? _GEN_3312 : valid_204; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4339 = _array_io_en_T_1 ? _GEN_3313 : valid_205; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4340 = _array_io_en_T_1 ? _GEN_3314 : valid_206; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4341 = _array_io_en_T_1 ? _GEN_3315 : valid_207; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4342 = _array_io_en_T_1 ? _GEN_3316 : valid_208; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4343 = _array_io_en_T_1 ? _GEN_3317 : valid_209; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4344 = _array_io_en_T_1 ? _GEN_3318 : valid_210; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4345 = _array_io_en_T_1 ? _GEN_3319 : valid_211; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4346 = _array_io_en_T_1 ? _GEN_3320 : valid_212; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4347 = _array_io_en_T_1 ? _GEN_3321 : valid_213; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4348 = _array_io_en_T_1 ? _GEN_3322 : valid_214; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4349 = _array_io_en_T_1 ? _GEN_3323 : valid_215; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4350 = _array_io_en_T_1 ? _GEN_3324 : valid_216; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4351 = _array_io_en_T_1 ? _GEN_3325 : valid_217; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4352 = _array_io_en_T_1 ? _GEN_3326 : valid_218; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4353 = _array_io_en_T_1 ? _GEN_3327 : valid_219; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4354 = _array_io_en_T_1 ? _GEN_3328 : valid_220; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4355 = _array_io_en_T_1 ? _GEN_3329 : valid_221; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4356 = _array_io_en_T_1 ? _GEN_3330 : valid_222; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4357 = _array_io_en_T_1 ? _GEN_3331 : valid_223; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4358 = _array_io_en_T_1 ? _GEN_3332 : valid_224; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4359 = _array_io_en_T_1 ? _GEN_3333 : valid_225; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4360 = _array_io_en_T_1 ? _GEN_3334 : valid_226; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4361 = _array_io_en_T_1 ? _GEN_3335 : valid_227; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4362 = _array_io_en_T_1 ? _GEN_3336 : valid_228; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4363 = _array_io_en_T_1 ? _GEN_3337 : valid_229; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4364 = _array_io_en_T_1 ? _GEN_3338 : valid_230; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4365 = _array_io_en_T_1 ? _GEN_3339 : valid_231; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4366 = _array_io_en_T_1 ? _GEN_3340 : valid_232; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4367 = _array_io_en_T_1 ? _GEN_3341 : valid_233; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4368 = _array_io_en_T_1 ? _GEN_3342 : valid_234; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4369 = _array_io_en_T_1 ? _GEN_3343 : valid_235; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4370 = _array_io_en_T_1 ? _GEN_3344 : valid_236; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4371 = _array_io_en_T_1 ? _GEN_3345 : valid_237; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4372 = _array_io_en_T_1 ? _GEN_3346 : valid_238; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4373 = _array_io_en_T_1 ? _GEN_3347 : valid_239; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4374 = _array_io_en_T_1 ? _GEN_3348 : valid_240; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4375 = _array_io_en_T_1 ? _GEN_3349 : valid_241; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4376 = _array_io_en_T_1 ? _GEN_3350 : valid_242; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4377 = _array_io_en_T_1 ? _GEN_3351 : valid_243; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4378 = _array_io_en_T_1 ? _GEN_3352 : valid_244; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4379 = _array_io_en_T_1 ? _GEN_3353 : valid_245; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4380 = _array_io_en_T_1 ? _GEN_3354 : valid_246; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4381 = _array_io_en_T_1 ? _GEN_3355 : valid_247; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4382 = _array_io_en_T_1 ? _GEN_3356 : valid_248; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4383 = _array_io_en_T_1 ? _GEN_3357 : valid_249; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4384 = _array_io_en_T_1 ? _GEN_3358 : valid_250; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4385 = _array_io_en_T_1 ? _GEN_3359 : valid_251; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4386 = _array_io_en_T_1 ? _GEN_3360 : valid_252; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4387 = _array_io_en_T_1 ? _GEN_3361 : valid_253; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4388 = _array_io_en_T_1 ? _GEN_3362 : valid_254; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4389 = _array_io_en_T_1 ? _GEN_3363 : valid_255; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4390 = _array_io_en_T_1 ? _GEN_3364 : valid_256; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4391 = _array_io_en_T_1 ? _GEN_3365 : valid_257; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4392 = _array_io_en_T_1 ? _GEN_3366 : valid_258; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4393 = _array_io_en_T_1 ? _GEN_3367 : valid_259; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4394 = _array_io_en_T_1 ? _GEN_3368 : valid_260; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4395 = _array_io_en_T_1 ? _GEN_3369 : valid_261; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4396 = _array_io_en_T_1 ? _GEN_3370 : valid_262; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4397 = _array_io_en_T_1 ? _GEN_3371 : valid_263; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4398 = _array_io_en_T_1 ? _GEN_3372 : valid_264; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4399 = _array_io_en_T_1 ? _GEN_3373 : valid_265; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4400 = _array_io_en_T_1 ? _GEN_3374 : valid_266; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4401 = _array_io_en_T_1 ? _GEN_3375 : valid_267; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4402 = _array_io_en_T_1 ? _GEN_3376 : valid_268; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4403 = _array_io_en_T_1 ? _GEN_3377 : valid_269; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4404 = _array_io_en_T_1 ? _GEN_3378 : valid_270; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4405 = _array_io_en_T_1 ? _GEN_3379 : valid_271; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4406 = _array_io_en_T_1 ? _GEN_3380 : valid_272; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4407 = _array_io_en_T_1 ? _GEN_3381 : valid_273; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4408 = _array_io_en_T_1 ? _GEN_3382 : valid_274; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4409 = _array_io_en_T_1 ? _GEN_3383 : valid_275; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4410 = _array_io_en_T_1 ? _GEN_3384 : valid_276; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4411 = _array_io_en_T_1 ? _GEN_3385 : valid_277; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4412 = _array_io_en_T_1 ? _GEN_3386 : valid_278; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4413 = _array_io_en_T_1 ? _GEN_3387 : valid_279; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4414 = _array_io_en_T_1 ? _GEN_3388 : valid_280; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4415 = _array_io_en_T_1 ? _GEN_3389 : valid_281; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4416 = _array_io_en_T_1 ? _GEN_3390 : valid_282; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4417 = _array_io_en_T_1 ? _GEN_3391 : valid_283; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4418 = _array_io_en_T_1 ? _GEN_3392 : valid_284; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4419 = _array_io_en_T_1 ? _GEN_3393 : valid_285; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4420 = _array_io_en_T_1 ? _GEN_3394 : valid_286; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4421 = _array_io_en_T_1 ? _GEN_3395 : valid_287; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4422 = _array_io_en_T_1 ? _GEN_3396 : valid_288; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4423 = _array_io_en_T_1 ? _GEN_3397 : valid_289; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4424 = _array_io_en_T_1 ? _GEN_3398 : valid_290; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4425 = _array_io_en_T_1 ? _GEN_3399 : valid_291; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4426 = _array_io_en_T_1 ? _GEN_3400 : valid_292; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4427 = _array_io_en_T_1 ? _GEN_3401 : valid_293; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4428 = _array_io_en_T_1 ? _GEN_3402 : valid_294; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4429 = _array_io_en_T_1 ? _GEN_3403 : valid_295; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4430 = _array_io_en_T_1 ? _GEN_3404 : valid_296; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4431 = _array_io_en_T_1 ? _GEN_3405 : valid_297; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4432 = _array_io_en_T_1 ? _GEN_3406 : valid_298; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4433 = _array_io_en_T_1 ? _GEN_3407 : valid_299; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4434 = _array_io_en_T_1 ? _GEN_3408 : valid_300; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4435 = _array_io_en_T_1 ? _GEN_3409 : valid_301; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4436 = _array_io_en_T_1 ? _GEN_3410 : valid_302; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4437 = _array_io_en_T_1 ? _GEN_3411 : valid_303; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4438 = _array_io_en_T_1 ? _GEN_3412 : valid_304; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4439 = _array_io_en_T_1 ? _GEN_3413 : valid_305; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4440 = _array_io_en_T_1 ? _GEN_3414 : valid_306; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4441 = _array_io_en_T_1 ? _GEN_3415 : valid_307; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4442 = _array_io_en_T_1 ? _GEN_3416 : valid_308; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4443 = _array_io_en_T_1 ? _GEN_3417 : valid_309; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4444 = _array_io_en_T_1 ? _GEN_3418 : valid_310; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4445 = _array_io_en_T_1 ? _GEN_3419 : valid_311; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4446 = _array_io_en_T_1 ? _GEN_3420 : valid_312; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4447 = _array_io_en_T_1 ? _GEN_3421 : valid_313; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4448 = _array_io_en_T_1 ? _GEN_3422 : valid_314; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4449 = _array_io_en_T_1 ? _GEN_3423 : valid_315; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4450 = _array_io_en_T_1 ? _GEN_3424 : valid_316; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4451 = _array_io_en_T_1 ? _GEN_3425 : valid_317; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4452 = _array_io_en_T_1 ? _GEN_3426 : valid_318; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4453 = _array_io_en_T_1 ? _GEN_3427 : valid_319; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4454 = _array_io_en_T_1 ? _GEN_3428 : valid_320; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4455 = _array_io_en_T_1 ? _GEN_3429 : valid_321; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4456 = _array_io_en_T_1 ? _GEN_3430 : valid_322; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4457 = _array_io_en_T_1 ? _GEN_3431 : valid_323; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4458 = _array_io_en_T_1 ? _GEN_3432 : valid_324; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4459 = _array_io_en_T_1 ? _GEN_3433 : valid_325; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4460 = _array_io_en_T_1 ? _GEN_3434 : valid_326; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4461 = _array_io_en_T_1 ? _GEN_3435 : valid_327; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4462 = _array_io_en_T_1 ? _GEN_3436 : valid_328; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4463 = _array_io_en_T_1 ? _GEN_3437 : valid_329; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4464 = _array_io_en_T_1 ? _GEN_3438 : valid_330; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4465 = _array_io_en_T_1 ? _GEN_3439 : valid_331; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4466 = _array_io_en_T_1 ? _GEN_3440 : valid_332; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4467 = _array_io_en_T_1 ? _GEN_3441 : valid_333; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4468 = _array_io_en_T_1 ? _GEN_3442 : valid_334; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4469 = _array_io_en_T_1 ? _GEN_3443 : valid_335; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4470 = _array_io_en_T_1 ? _GEN_3444 : valid_336; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4471 = _array_io_en_T_1 ? _GEN_3445 : valid_337; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4472 = _array_io_en_T_1 ? _GEN_3446 : valid_338; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4473 = _array_io_en_T_1 ? _GEN_3447 : valid_339; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4474 = _array_io_en_T_1 ? _GEN_3448 : valid_340; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4475 = _array_io_en_T_1 ? _GEN_3449 : valid_341; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4476 = _array_io_en_T_1 ? _GEN_3450 : valid_342; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4477 = _array_io_en_T_1 ? _GEN_3451 : valid_343; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4478 = _array_io_en_T_1 ? _GEN_3452 : valid_344; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4479 = _array_io_en_T_1 ? _GEN_3453 : valid_345; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4480 = _array_io_en_T_1 ? _GEN_3454 : valid_346; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4481 = _array_io_en_T_1 ? _GEN_3455 : valid_347; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4482 = _array_io_en_T_1 ? _GEN_3456 : valid_348; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4483 = _array_io_en_T_1 ? _GEN_3457 : valid_349; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4484 = _array_io_en_T_1 ? _GEN_3458 : valid_350; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4485 = _array_io_en_T_1 ? _GEN_3459 : valid_351; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4486 = _array_io_en_T_1 ? _GEN_3460 : valid_352; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4487 = _array_io_en_T_1 ? _GEN_3461 : valid_353; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4488 = _array_io_en_T_1 ? _GEN_3462 : valid_354; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4489 = _array_io_en_T_1 ? _GEN_3463 : valid_355; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4490 = _array_io_en_T_1 ? _GEN_3464 : valid_356; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4491 = _array_io_en_T_1 ? _GEN_3465 : valid_357; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4492 = _array_io_en_T_1 ? _GEN_3466 : valid_358; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4493 = _array_io_en_T_1 ? _GEN_3467 : valid_359; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4494 = _array_io_en_T_1 ? _GEN_3468 : valid_360; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4495 = _array_io_en_T_1 ? _GEN_3469 : valid_361; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4496 = _array_io_en_T_1 ? _GEN_3470 : valid_362; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4497 = _array_io_en_T_1 ? _GEN_3471 : valid_363; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4498 = _array_io_en_T_1 ? _GEN_3472 : valid_364; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4499 = _array_io_en_T_1 ? _GEN_3473 : valid_365; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4500 = _array_io_en_T_1 ? _GEN_3474 : valid_366; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4501 = _array_io_en_T_1 ? _GEN_3475 : valid_367; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4502 = _array_io_en_T_1 ? _GEN_3476 : valid_368; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4503 = _array_io_en_T_1 ? _GEN_3477 : valid_369; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4504 = _array_io_en_T_1 ? _GEN_3478 : valid_370; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4505 = _array_io_en_T_1 ? _GEN_3479 : valid_371; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4506 = _array_io_en_T_1 ? _GEN_3480 : valid_372; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4507 = _array_io_en_T_1 ? _GEN_3481 : valid_373; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4508 = _array_io_en_T_1 ? _GEN_3482 : valid_374; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4509 = _array_io_en_T_1 ? _GEN_3483 : valid_375; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4510 = _array_io_en_T_1 ? _GEN_3484 : valid_376; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4511 = _array_io_en_T_1 ? _GEN_3485 : valid_377; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4512 = _array_io_en_T_1 ? _GEN_3486 : valid_378; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4513 = _array_io_en_T_1 ? _GEN_3487 : valid_379; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4514 = _array_io_en_T_1 ? _GEN_3488 : valid_380; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4515 = _array_io_en_T_1 ? _GEN_3489 : valid_381; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4516 = _array_io_en_T_1 ? _GEN_3490 : valid_382; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4517 = _array_io_en_T_1 ? _GEN_3491 : valid_383; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4518 = _array_io_en_T_1 ? _GEN_3492 : valid_384; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4519 = _array_io_en_T_1 ? _GEN_3493 : valid_385; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4520 = _array_io_en_T_1 ? _GEN_3494 : valid_386; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4521 = _array_io_en_T_1 ? _GEN_3495 : valid_387; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4522 = _array_io_en_T_1 ? _GEN_3496 : valid_388; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4523 = _array_io_en_T_1 ? _GEN_3497 : valid_389; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4524 = _array_io_en_T_1 ? _GEN_3498 : valid_390; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4525 = _array_io_en_T_1 ? _GEN_3499 : valid_391; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4526 = _array_io_en_T_1 ? _GEN_3500 : valid_392; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4527 = _array_io_en_T_1 ? _GEN_3501 : valid_393; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4528 = _array_io_en_T_1 ? _GEN_3502 : valid_394; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4529 = _array_io_en_T_1 ? _GEN_3503 : valid_395; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4530 = _array_io_en_T_1 ? _GEN_3504 : valid_396; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4531 = _array_io_en_T_1 ? _GEN_3505 : valid_397; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4532 = _array_io_en_T_1 ? _GEN_3506 : valid_398; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4533 = _array_io_en_T_1 ? _GEN_3507 : valid_399; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4534 = _array_io_en_T_1 ? _GEN_3508 : valid_400; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4535 = _array_io_en_T_1 ? _GEN_3509 : valid_401; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4536 = _array_io_en_T_1 ? _GEN_3510 : valid_402; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4537 = _array_io_en_T_1 ? _GEN_3511 : valid_403; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4538 = _array_io_en_T_1 ? _GEN_3512 : valid_404; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4539 = _array_io_en_T_1 ? _GEN_3513 : valid_405; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4540 = _array_io_en_T_1 ? _GEN_3514 : valid_406; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4541 = _array_io_en_T_1 ? _GEN_3515 : valid_407; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4542 = _array_io_en_T_1 ? _GEN_3516 : valid_408; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4543 = _array_io_en_T_1 ? _GEN_3517 : valid_409; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4544 = _array_io_en_T_1 ? _GEN_3518 : valid_410; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4545 = _array_io_en_T_1 ? _GEN_3519 : valid_411; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4546 = _array_io_en_T_1 ? _GEN_3520 : valid_412; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4547 = _array_io_en_T_1 ? _GEN_3521 : valid_413; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4548 = _array_io_en_T_1 ? _GEN_3522 : valid_414; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4549 = _array_io_en_T_1 ? _GEN_3523 : valid_415; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4550 = _array_io_en_T_1 ? _GEN_3524 : valid_416; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4551 = _array_io_en_T_1 ? _GEN_3525 : valid_417; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4552 = _array_io_en_T_1 ? _GEN_3526 : valid_418; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4553 = _array_io_en_T_1 ? _GEN_3527 : valid_419; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4554 = _array_io_en_T_1 ? _GEN_3528 : valid_420; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4555 = _array_io_en_T_1 ? _GEN_3529 : valid_421; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4556 = _array_io_en_T_1 ? _GEN_3530 : valid_422; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4557 = _array_io_en_T_1 ? _GEN_3531 : valid_423; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4558 = _array_io_en_T_1 ? _GEN_3532 : valid_424; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4559 = _array_io_en_T_1 ? _GEN_3533 : valid_425; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4560 = _array_io_en_T_1 ? _GEN_3534 : valid_426; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4561 = _array_io_en_T_1 ? _GEN_3535 : valid_427; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4562 = _array_io_en_T_1 ? _GEN_3536 : valid_428; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4563 = _array_io_en_T_1 ? _GEN_3537 : valid_429; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4564 = _array_io_en_T_1 ? _GEN_3538 : valid_430; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4565 = _array_io_en_T_1 ? _GEN_3539 : valid_431; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4566 = _array_io_en_T_1 ? _GEN_3540 : valid_432; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4567 = _array_io_en_T_1 ? _GEN_3541 : valid_433; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4568 = _array_io_en_T_1 ? _GEN_3542 : valid_434; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4569 = _array_io_en_T_1 ? _GEN_3543 : valid_435; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4570 = _array_io_en_T_1 ? _GEN_3544 : valid_436; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4571 = _array_io_en_T_1 ? _GEN_3545 : valid_437; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4572 = _array_io_en_T_1 ? _GEN_3546 : valid_438; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4573 = _array_io_en_T_1 ? _GEN_3547 : valid_439; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4574 = _array_io_en_T_1 ? _GEN_3548 : valid_440; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4575 = _array_io_en_T_1 ? _GEN_3549 : valid_441; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4576 = _array_io_en_T_1 ? _GEN_3550 : valid_442; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4577 = _array_io_en_T_1 ? _GEN_3551 : valid_443; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4578 = _array_io_en_T_1 ? _GEN_3552 : valid_444; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4579 = _array_io_en_T_1 ? _GEN_3553 : valid_445; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4580 = _array_io_en_T_1 ? _GEN_3554 : valid_446; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4581 = _array_io_en_T_1 ? _GEN_3555 : valid_447; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4582 = _array_io_en_T_1 ? _GEN_3556 : valid_448; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4583 = _array_io_en_T_1 ? _GEN_3557 : valid_449; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4584 = _array_io_en_T_1 ? _GEN_3558 : valid_450; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4585 = _array_io_en_T_1 ? _GEN_3559 : valid_451; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4586 = _array_io_en_T_1 ? _GEN_3560 : valid_452; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4587 = _array_io_en_T_1 ? _GEN_3561 : valid_453; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4588 = _array_io_en_T_1 ? _GEN_3562 : valid_454; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4589 = _array_io_en_T_1 ? _GEN_3563 : valid_455; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4590 = _array_io_en_T_1 ? _GEN_3564 : valid_456; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4591 = _array_io_en_T_1 ? _GEN_3565 : valid_457; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4592 = _array_io_en_T_1 ? _GEN_3566 : valid_458; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4593 = _array_io_en_T_1 ? _GEN_3567 : valid_459; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4594 = _array_io_en_T_1 ? _GEN_3568 : valid_460; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4595 = _array_io_en_T_1 ? _GEN_3569 : valid_461; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4596 = _array_io_en_T_1 ? _GEN_3570 : valid_462; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4597 = _array_io_en_T_1 ? _GEN_3571 : valid_463; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4598 = _array_io_en_T_1 ? _GEN_3572 : valid_464; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4599 = _array_io_en_T_1 ? _GEN_3573 : valid_465; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4600 = _array_io_en_T_1 ? _GEN_3574 : valid_466; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4601 = _array_io_en_T_1 ? _GEN_3575 : valid_467; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4602 = _array_io_en_T_1 ? _GEN_3576 : valid_468; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4603 = _array_io_en_T_1 ? _GEN_3577 : valid_469; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4604 = _array_io_en_T_1 ? _GEN_3578 : valid_470; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4605 = _array_io_en_T_1 ? _GEN_3579 : valid_471; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4606 = _array_io_en_T_1 ? _GEN_3580 : valid_472; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4607 = _array_io_en_T_1 ? _GEN_3581 : valid_473; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4608 = _array_io_en_T_1 ? _GEN_3582 : valid_474; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4609 = _array_io_en_T_1 ? _GEN_3583 : valid_475; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4610 = _array_io_en_T_1 ? _GEN_3584 : valid_476; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4611 = _array_io_en_T_1 ? _GEN_3585 : valid_477; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4612 = _array_io_en_T_1 ? _GEN_3586 : valid_478; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4613 = _array_io_en_T_1 ? _GEN_3587 : valid_479; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4614 = _array_io_en_T_1 ? _GEN_3588 : valid_480; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4615 = _array_io_en_T_1 ? _GEN_3589 : valid_481; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4616 = _array_io_en_T_1 ? _GEN_3590 : valid_482; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4617 = _array_io_en_T_1 ? _GEN_3591 : valid_483; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4618 = _array_io_en_T_1 ? _GEN_3592 : valid_484; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4619 = _array_io_en_T_1 ? _GEN_3593 : valid_485; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4620 = _array_io_en_T_1 ? _GEN_3594 : valid_486; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4621 = _array_io_en_T_1 ? _GEN_3595 : valid_487; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4622 = _array_io_en_T_1 ? _GEN_3596 : valid_488; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4623 = _array_io_en_T_1 ? _GEN_3597 : valid_489; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4624 = _array_io_en_T_1 ? _GEN_3598 : valid_490; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4625 = _array_io_en_T_1 ? _GEN_3599 : valid_491; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4626 = _array_io_en_T_1 ? _GEN_3600 : valid_492; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4627 = _array_io_en_T_1 ? _GEN_3601 : valid_493; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4628 = _array_io_en_T_1 ? _GEN_3602 : valid_494; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4629 = _array_io_en_T_1 ? _GEN_3603 : valid_495; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4630 = _array_io_en_T_1 ? _GEN_3604 : valid_496; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4631 = _array_io_en_T_1 ? _GEN_3605 : valid_497; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4632 = _array_io_en_T_1 ? _GEN_3606 : valid_498; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4633 = _array_io_en_T_1 ? _GEN_3607 : valid_499; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4634 = _array_io_en_T_1 ? _GEN_3608 : valid_500; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4635 = _array_io_en_T_1 ? _GEN_3609 : valid_501; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4636 = _array_io_en_T_1 ? _GEN_3610 : valid_502; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4637 = _array_io_en_T_1 ? _GEN_3611 : valid_503; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4638 = _array_io_en_T_1 ? _GEN_3612 : valid_504; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4639 = _array_io_en_T_1 ? _GEN_3613 : valid_505; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4640 = _array_io_en_T_1 ? _GEN_3614 : valid_506; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4641 = _array_io_en_T_1 ? _GEN_3615 : valid_507; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4642 = _array_io_en_T_1 ? _GEN_3616 : valid_508; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4643 = _array_io_en_T_1 ? _GEN_3617 : valid_509; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4644 = _array_io_en_T_1 ? _GEN_3618 : valid_510; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4645 = _array_io_en_T_1 ? _GEN_3619 : valid_511; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4646 = _array_io_en_T_1 ? _GEN_3620 : valid_512; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4647 = _array_io_en_T_1 ? _GEN_3621 : valid_513; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4648 = _array_io_en_T_1 ? _GEN_3622 : valid_514; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4649 = _array_io_en_T_1 ? _GEN_3623 : valid_515; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4650 = _array_io_en_T_1 ? _GEN_3624 : valid_516; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4651 = _array_io_en_T_1 ? _GEN_3625 : valid_517; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4652 = _array_io_en_T_1 ? _GEN_3626 : valid_518; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4653 = _array_io_en_T_1 ? _GEN_3627 : valid_519; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4654 = _array_io_en_T_1 ? _GEN_3628 : valid_520; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4655 = _array_io_en_T_1 ? _GEN_3629 : valid_521; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4656 = _array_io_en_T_1 ? _GEN_3630 : valid_522; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4657 = _array_io_en_T_1 ? _GEN_3631 : valid_523; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4658 = _array_io_en_T_1 ? _GEN_3632 : valid_524; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4659 = _array_io_en_T_1 ? _GEN_3633 : valid_525; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4660 = _array_io_en_T_1 ? _GEN_3634 : valid_526; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4661 = _array_io_en_T_1 ? _GEN_3635 : valid_527; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4662 = _array_io_en_T_1 ? _GEN_3636 : valid_528; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4663 = _array_io_en_T_1 ? _GEN_3637 : valid_529; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4664 = _array_io_en_T_1 ? _GEN_3638 : valid_530; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4665 = _array_io_en_T_1 ? _GEN_3639 : valid_531; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4666 = _array_io_en_T_1 ? _GEN_3640 : valid_532; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4667 = _array_io_en_T_1 ? _GEN_3641 : valid_533; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4668 = _array_io_en_T_1 ? _GEN_3642 : valid_534; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4669 = _array_io_en_T_1 ? _GEN_3643 : valid_535; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4670 = _array_io_en_T_1 ? _GEN_3644 : valid_536; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4671 = _array_io_en_T_1 ? _GEN_3645 : valid_537; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4672 = _array_io_en_T_1 ? _GEN_3646 : valid_538; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4673 = _array_io_en_T_1 ? _GEN_3647 : valid_539; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4674 = _array_io_en_T_1 ? _GEN_3648 : valid_540; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4675 = _array_io_en_T_1 ? _GEN_3649 : valid_541; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4676 = _array_io_en_T_1 ? _GEN_3650 : valid_542; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4677 = _array_io_en_T_1 ? _GEN_3651 : valid_543; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4678 = _array_io_en_T_1 ? _GEN_3652 : valid_544; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4679 = _array_io_en_T_1 ? _GEN_3653 : valid_545; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4680 = _array_io_en_T_1 ? _GEN_3654 : valid_546; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4681 = _array_io_en_T_1 ? _GEN_3655 : valid_547; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4682 = _array_io_en_T_1 ? _GEN_3656 : valid_548; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4683 = _array_io_en_T_1 ? _GEN_3657 : valid_549; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4684 = _array_io_en_T_1 ? _GEN_3658 : valid_550; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4685 = _array_io_en_T_1 ? _GEN_3659 : valid_551; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4686 = _array_io_en_T_1 ? _GEN_3660 : valid_552; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4687 = _array_io_en_T_1 ? _GEN_3661 : valid_553; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4688 = _array_io_en_T_1 ? _GEN_3662 : valid_554; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4689 = _array_io_en_T_1 ? _GEN_3663 : valid_555; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4690 = _array_io_en_T_1 ? _GEN_3664 : valid_556; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4691 = _array_io_en_T_1 ? _GEN_3665 : valid_557; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4692 = _array_io_en_T_1 ? _GEN_3666 : valid_558; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4693 = _array_io_en_T_1 ? _GEN_3667 : valid_559; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4694 = _array_io_en_T_1 ? _GEN_3668 : valid_560; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4695 = _array_io_en_T_1 ? _GEN_3669 : valid_561; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4696 = _array_io_en_T_1 ? _GEN_3670 : valid_562; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4697 = _array_io_en_T_1 ? _GEN_3671 : valid_563; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4698 = _array_io_en_T_1 ? _GEN_3672 : valid_564; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4699 = _array_io_en_T_1 ? _GEN_3673 : valid_565; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4700 = _array_io_en_T_1 ? _GEN_3674 : valid_566; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4701 = _array_io_en_T_1 ? _GEN_3675 : valid_567; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4702 = _array_io_en_T_1 ? _GEN_3676 : valid_568; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4703 = _array_io_en_T_1 ? _GEN_3677 : valid_569; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4704 = _array_io_en_T_1 ? _GEN_3678 : valid_570; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4705 = _array_io_en_T_1 ? _GEN_3679 : valid_571; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4706 = _array_io_en_T_1 ? _GEN_3680 : valid_572; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4707 = _array_io_en_T_1 ? _GEN_3681 : valid_573; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4708 = _array_io_en_T_1 ? _GEN_3682 : valid_574; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4709 = _array_io_en_T_1 ? _GEN_3683 : valid_575; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4710 = _array_io_en_T_1 ? _GEN_3684 : valid_576; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4711 = _array_io_en_T_1 ? _GEN_3685 : valid_577; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4712 = _array_io_en_T_1 ? _GEN_3686 : valid_578; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4713 = _array_io_en_T_1 ? _GEN_3687 : valid_579; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4714 = _array_io_en_T_1 ? _GEN_3688 : valid_580; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4715 = _array_io_en_T_1 ? _GEN_3689 : valid_581; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4716 = _array_io_en_T_1 ? _GEN_3690 : valid_582; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4717 = _array_io_en_T_1 ? _GEN_3691 : valid_583; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4718 = _array_io_en_T_1 ? _GEN_3692 : valid_584; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4719 = _array_io_en_T_1 ? _GEN_3693 : valid_585; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4720 = _array_io_en_T_1 ? _GEN_3694 : valid_586; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4721 = _array_io_en_T_1 ? _GEN_3695 : valid_587; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4722 = _array_io_en_T_1 ? _GEN_3696 : valid_588; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4723 = _array_io_en_T_1 ? _GEN_3697 : valid_589; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4724 = _array_io_en_T_1 ? _GEN_3698 : valid_590; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4725 = _array_io_en_T_1 ? _GEN_3699 : valid_591; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4726 = _array_io_en_T_1 ? _GEN_3700 : valid_592; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4727 = _array_io_en_T_1 ? _GEN_3701 : valid_593; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4728 = _array_io_en_T_1 ? _GEN_3702 : valid_594; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4729 = _array_io_en_T_1 ? _GEN_3703 : valid_595; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4730 = _array_io_en_T_1 ? _GEN_3704 : valid_596; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4731 = _array_io_en_T_1 ? _GEN_3705 : valid_597; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4732 = _array_io_en_T_1 ? _GEN_3706 : valid_598; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4733 = _array_io_en_T_1 ? _GEN_3707 : valid_599; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4734 = _array_io_en_T_1 ? _GEN_3708 : valid_600; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4735 = _array_io_en_T_1 ? _GEN_3709 : valid_601; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4736 = _array_io_en_T_1 ? _GEN_3710 : valid_602; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4737 = _array_io_en_T_1 ? _GEN_3711 : valid_603; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4738 = _array_io_en_T_1 ? _GEN_3712 : valid_604; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4739 = _array_io_en_T_1 ? _GEN_3713 : valid_605; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4740 = _array_io_en_T_1 ? _GEN_3714 : valid_606; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4741 = _array_io_en_T_1 ? _GEN_3715 : valid_607; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4742 = _array_io_en_T_1 ? _GEN_3716 : valid_608; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4743 = _array_io_en_T_1 ? _GEN_3717 : valid_609; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4744 = _array_io_en_T_1 ? _GEN_3718 : valid_610; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4745 = _array_io_en_T_1 ? _GEN_3719 : valid_611; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4746 = _array_io_en_T_1 ? _GEN_3720 : valid_612; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4747 = _array_io_en_T_1 ? _GEN_3721 : valid_613; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4748 = _array_io_en_T_1 ? _GEN_3722 : valid_614; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4749 = _array_io_en_T_1 ? _GEN_3723 : valid_615; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4750 = _array_io_en_T_1 ? _GEN_3724 : valid_616; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4751 = _array_io_en_T_1 ? _GEN_3725 : valid_617; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4752 = _array_io_en_T_1 ? _GEN_3726 : valid_618; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4753 = _array_io_en_T_1 ? _GEN_3727 : valid_619; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4754 = _array_io_en_T_1 ? _GEN_3728 : valid_620; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4755 = _array_io_en_T_1 ? _GEN_3729 : valid_621; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4756 = _array_io_en_T_1 ? _GEN_3730 : valid_622; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4757 = _array_io_en_T_1 ? _GEN_3731 : valid_623; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4758 = _array_io_en_T_1 ? _GEN_3732 : valid_624; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4759 = _array_io_en_T_1 ? _GEN_3733 : valid_625; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4760 = _array_io_en_T_1 ? _GEN_3734 : valid_626; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4761 = _array_io_en_T_1 ? _GEN_3735 : valid_627; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4762 = _array_io_en_T_1 ? _GEN_3736 : valid_628; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4763 = _array_io_en_T_1 ? _GEN_3737 : valid_629; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4764 = _array_io_en_T_1 ? _GEN_3738 : valid_630; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4765 = _array_io_en_T_1 ? _GEN_3739 : valid_631; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4766 = _array_io_en_T_1 ? _GEN_3740 : valid_632; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4767 = _array_io_en_T_1 ? _GEN_3741 : valid_633; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4768 = _array_io_en_T_1 ? _GEN_3742 : valid_634; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4769 = _array_io_en_T_1 ? _GEN_3743 : valid_635; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4770 = _array_io_en_T_1 ? _GEN_3744 : valid_636; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4771 = _array_io_en_T_1 ? _GEN_3745 : valid_637; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4772 = _array_io_en_T_1 ? _GEN_3746 : valid_638; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4773 = _array_io_en_T_1 ? _GEN_3747 : valid_639; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4774 = _array_io_en_T_1 ? _GEN_3748 : valid_640; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4775 = _array_io_en_T_1 ? _GEN_3749 : valid_641; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4776 = _array_io_en_T_1 ? _GEN_3750 : valid_642; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4777 = _array_io_en_T_1 ? _GEN_3751 : valid_643; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4778 = _array_io_en_T_1 ? _GEN_3752 : valid_644; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4779 = _array_io_en_T_1 ? _GEN_3753 : valid_645; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4780 = _array_io_en_T_1 ? _GEN_3754 : valid_646; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4781 = _array_io_en_T_1 ? _GEN_3755 : valid_647; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4782 = _array_io_en_T_1 ? _GEN_3756 : valid_648; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4783 = _array_io_en_T_1 ? _GEN_3757 : valid_649; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4784 = _array_io_en_T_1 ? _GEN_3758 : valid_650; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4785 = _array_io_en_T_1 ? _GEN_3759 : valid_651; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4786 = _array_io_en_T_1 ? _GEN_3760 : valid_652; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4787 = _array_io_en_T_1 ? _GEN_3761 : valid_653; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4788 = _array_io_en_T_1 ? _GEN_3762 : valid_654; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4789 = _array_io_en_T_1 ? _GEN_3763 : valid_655; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4790 = _array_io_en_T_1 ? _GEN_3764 : valid_656; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4791 = _array_io_en_T_1 ? _GEN_3765 : valid_657; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4792 = _array_io_en_T_1 ? _GEN_3766 : valid_658; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4793 = _array_io_en_T_1 ? _GEN_3767 : valid_659; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4794 = _array_io_en_T_1 ? _GEN_3768 : valid_660; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4795 = _array_io_en_T_1 ? _GEN_3769 : valid_661; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4796 = _array_io_en_T_1 ? _GEN_3770 : valid_662; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4797 = _array_io_en_T_1 ? _GEN_3771 : valid_663; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4798 = _array_io_en_T_1 ? _GEN_3772 : valid_664; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4799 = _array_io_en_T_1 ? _GEN_3773 : valid_665; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4800 = _array_io_en_T_1 ? _GEN_3774 : valid_666; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4801 = _array_io_en_T_1 ? _GEN_3775 : valid_667; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4802 = _array_io_en_T_1 ? _GEN_3776 : valid_668; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4803 = _array_io_en_T_1 ? _GEN_3777 : valid_669; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4804 = _array_io_en_T_1 ? _GEN_3778 : valid_670; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4805 = _array_io_en_T_1 ? _GEN_3779 : valid_671; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4806 = _array_io_en_T_1 ? _GEN_3780 : valid_672; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4807 = _array_io_en_T_1 ? _GEN_3781 : valid_673; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4808 = _array_io_en_T_1 ? _GEN_3782 : valid_674; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4809 = _array_io_en_T_1 ? _GEN_3783 : valid_675; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4810 = _array_io_en_T_1 ? _GEN_3784 : valid_676; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4811 = _array_io_en_T_1 ? _GEN_3785 : valid_677; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4812 = _array_io_en_T_1 ? _GEN_3786 : valid_678; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4813 = _array_io_en_T_1 ? _GEN_3787 : valid_679; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4814 = _array_io_en_T_1 ? _GEN_3788 : valid_680; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4815 = _array_io_en_T_1 ? _GEN_3789 : valid_681; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4816 = _array_io_en_T_1 ? _GEN_3790 : valid_682; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4817 = _array_io_en_T_1 ? _GEN_3791 : valid_683; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4818 = _array_io_en_T_1 ? _GEN_3792 : valid_684; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4819 = _array_io_en_T_1 ? _GEN_3793 : valid_685; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4820 = _array_io_en_T_1 ? _GEN_3794 : valid_686; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4821 = _array_io_en_T_1 ? _GEN_3795 : valid_687; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4822 = _array_io_en_T_1 ? _GEN_3796 : valid_688; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4823 = _array_io_en_T_1 ? _GEN_3797 : valid_689; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4824 = _array_io_en_T_1 ? _GEN_3798 : valid_690; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4825 = _array_io_en_T_1 ? _GEN_3799 : valid_691; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4826 = _array_io_en_T_1 ? _GEN_3800 : valid_692; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4827 = _array_io_en_T_1 ? _GEN_3801 : valid_693; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4828 = _array_io_en_T_1 ? _GEN_3802 : valid_694; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4829 = _array_io_en_T_1 ? _GEN_3803 : valid_695; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4830 = _array_io_en_T_1 ? _GEN_3804 : valid_696; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4831 = _array_io_en_T_1 ? _GEN_3805 : valid_697; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4832 = _array_io_en_T_1 ? _GEN_3806 : valid_698; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4833 = _array_io_en_T_1 ? _GEN_3807 : valid_699; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4834 = _array_io_en_T_1 ? _GEN_3808 : valid_700; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4835 = _array_io_en_T_1 ? _GEN_3809 : valid_701; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4836 = _array_io_en_T_1 ? _GEN_3810 : valid_702; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4837 = _array_io_en_T_1 ? _GEN_3811 : valid_703; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4838 = _array_io_en_T_1 ? _GEN_3812 : valid_704; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4839 = _array_io_en_T_1 ? _GEN_3813 : valid_705; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4840 = _array_io_en_T_1 ? _GEN_3814 : valid_706; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4841 = _array_io_en_T_1 ? _GEN_3815 : valid_707; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4842 = _array_io_en_T_1 ? _GEN_3816 : valid_708; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4843 = _array_io_en_T_1 ? _GEN_3817 : valid_709; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4844 = _array_io_en_T_1 ? _GEN_3818 : valid_710; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4845 = _array_io_en_T_1 ? _GEN_3819 : valid_711; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4846 = _array_io_en_T_1 ? _GEN_3820 : valid_712; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4847 = _array_io_en_T_1 ? _GEN_3821 : valid_713; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4848 = _array_io_en_T_1 ? _GEN_3822 : valid_714; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4849 = _array_io_en_T_1 ? _GEN_3823 : valid_715; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4850 = _array_io_en_T_1 ? _GEN_3824 : valid_716; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4851 = _array_io_en_T_1 ? _GEN_3825 : valid_717; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4852 = _array_io_en_T_1 ? _GEN_3826 : valid_718; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4853 = _array_io_en_T_1 ? _GEN_3827 : valid_719; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4854 = _array_io_en_T_1 ? _GEN_3828 : valid_720; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4855 = _array_io_en_T_1 ? _GEN_3829 : valid_721; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4856 = _array_io_en_T_1 ? _GEN_3830 : valid_722; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4857 = _array_io_en_T_1 ? _GEN_3831 : valid_723; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4858 = _array_io_en_T_1 ? _GEN_3832 : valid_724; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4859 = _array_io_en_T_1 ? _GEN_3833 : valid_725; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4860 = _array_io_en_T_1 ? _GEN_3834 : valid_726; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4861 = _array_io_en_T_1 ? _GEN_3835 : valid_727; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4862 = _array_io_en_T_1 ? _GEN_3836 : valid_728; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4863 = _array_io_en_T_1 ? _GEN_3837 : valid_729; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4864 = _array_io_en_T_1 ? _GEN_3838 : valid_730; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4865 = _array_io_en_T_1 ? _GEN_3839 : valid_731; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4866 = _array_io_en_T_1 ? _GEN_3840 : valid_732; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4867 = _array_io_en_T_1 ? _GEN_3841 : valid_733; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4868 = _array_io_en_T_1 ? _GEN_3842 : valid_734; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4869 = _array_io_en_T_1 ? _GEN_3843 : valid_735; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4870 = _array_io_en_T_1 ? _GEN_3844 : valid_736; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4871 = _array_io_en_T_1 ? _GEN_3845 : valid_737; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4872 = _array_io_en_T_1 ? _GEN_3846 : valid_738; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4873 = _array_io_en_T_1 ? _GEN_3847 : valid_739; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4874 = _array_io_en_T_1 ? _GEN_3848 : valid_740; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4875 = _array_io_en_T_1 ? _GEN_3849 : valid_741; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4876 = _array_io_en_T_1 ? _GEN_3850 : valid_742; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4877 = _array_io_en_T_1 ? _GEN_3851 : valid_743; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4878 = _array_io_en_T_1 ? _GEN_3852 : valid_744; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4879 = _array_io_en_T_1 ? _GEN_3853 : valid_745; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4880 = _array_io_en_T_1 ? _GEN_3854 : valid_746; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4881 = _array_io_en_T_1 ? _GEN_3855 : valid_747; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4882 = _array_io_en_T_1 ? _GEN_3856 : valid_748; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4883 = _array_io_en_T_1 ? _GEN_3857 : valid_749; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4884 = _array_io_en_T_1 ? _GEN_3858 : valid_750; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4885 = _array_io_en_T_1 ? _GEN_3859 : valid_751; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4886 = _array_io_en_T_1 ? _GEN_3860 : valid_752; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4887 = _array_io_en_T_1 ? _GEN_3861 : valid_753; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4888 = _array_io_en_T_1 ? _GEN_3862 : valid_754; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4889 = _array_io_en_T_1 ? _GEN_3863 : valid_755; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4890 = _array_io_en_T_1 ? _GEN_3864 : valid_756; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4891 = _array_io_en_T_1 ? _GEN_3865 : valid_757; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4892 = _array_io_en_T_1 ? _GEN_3866 : valid_758; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4893 = _array_io_en_T_1 ? _GEN_3867 : valid_759; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4894 = _array_io_en_T_1 ? _GEN_3868 : valid_760; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4895 = _array_io_en_T_1 ? _GEN_3869 : valid_761; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4896 = _array_io_en_T_1 ? _GEN_3870 : valid_762; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4897 = _array_io_en_T_1 ? _GEN_3871 : valid_763; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4898 = _array_io_en_T_1 ? _GEN_3872 : valid_764; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4899 = _array_io_en_T_1 ? _GEN_3873 : valid_765; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4900 = _array_io_en_T_1 ? _GEN_3874 : valid_766; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4901 = _array_io_en_T_1 ? _GEN_3875 : valid_767; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4902 = _array_io_en_T_1 ? _GEN_3876 : valid_768; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4903 = _array_io_en_T_1 ? _GEN_3877 : valid_769; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4904 = _array_io_en_T_1 ? _GEN_3878 : valid_770; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4905 = _array_io_en_T_1 ? _GEN_3879 : valid_771; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4906 = _array_io_en_T_1 ? _GEN_3880 : valid_772; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4907 = _array_io_en_T_1 ? _GEN_3881 : valid_773; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4908 = _array_io_en_T_1 ? _GEN_3882 : valid_774; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4909 = _array_io_en_T_1 ? _GEN_3883 : valid_775; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4910 = _array_io_en_T_1 ? _GEN_3884 : valid_776; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4911 = _array_io_en_T_1 ? _GEN_3885 : valid_777; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4912 = _array_io_en_T_1 ? _GEN_3886 : valid_778; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4913 = _array_io_en_T_1 ? _GEN_3887 : valid_779; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4914 = _array_io_en_T_1 ? _GEN_3888 : valid_780; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4915 = _array_io_en_T_1 ? _GEN_3889 : valid_781; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4916 = _array_io_en_T_1 ? _GEN_3890 : valid_782; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4917 = _array_io_en_T_1 ? _GEN_3891 : valid_783; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4918 = _array_io_en_T_1 ? _GEN_3892 : valid_784; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4919 = _array_io_en_T_1 ? _GEN_3893 : valid_785; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4920 = _array_io_en_T_1 ? _GEN_3894 : valid_786; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4921 = _array_io_en_T_1 ? _GEN_3895 : valid_787; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4922 = _array_io_en_T_1 ? _GEN_3896 : valid_788; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4923 = _array_io_en_T_1 ? _GEN_3897 : valid_789; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4924 = _array_io_en_T_1 ? _GEN_3898 : valid_790; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4925 = _array_io_en_T_1 ? _GEN_3899 : valid_791; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4926 = _array_io_en_T_1 ? _GEN_3900 : valid_792; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4927 = _array_io_en_T_1 ? _GEN_3901 : valid_793; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4928 = _array_io_en_T_1 ? _GEN_3902 : valid_794; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4929 = _array_io_en_T_1 ? _GEN_3903 : valid_795; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4930 = _array_io_en_T_1 ? _GEN_3904 : valid_796; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4931 = _array_io_en_T_1 ? _GEN_3905 : valid_797; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4932 = _array_io_en_T_1 ? _GEN_3906 : valid_798; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4933 = _array_io_en_T_1 ? _GEN_3907 : valid_799; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4934 = _array_io_en_T_1 ? _GEN_3908 : valid_800; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4935 = _array_io_en_T_1 ? _GEN_3909 : valid_801; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4936 = _array_io_en_T_1 ? _GEN_3910 : valid_802; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4937 = _array_io_en_T_1 ? _GEN_3911 : valid_803; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4938 = _array_io_en_T_1 ? _GEN_3912 : valid_804; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4939 = _array_io_en_T_1 ? _GEN_3913 : valid_805; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4940 = _array_io_en_T_1 ? _GEN_3914 : valid_806; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4941 = _array_io_en_T_1 ? _GEN_3915 : valid_807; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4942 = _array_io_en_T_1 ? _GEN_3916 : valid_808; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4943 = _array_io_en_T_1 ? _GEN_3917 : valid_809; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4944 = _array_io_en_T_1 ? _GEN_3918 : valid_810; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4945 = _array_io_en_T_1 ? _GEN_3919 : valid_811; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4946 = _array_io_en_T_1 ? _GEN_3920 : valid_812; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4947 = _array_io_en_T_1 ? _GEN_3921 : valid_813; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4948 = _array_io_en_T_1 ? _GEN_3922 : valid_814; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4949 = _array_io_en_T_1 ? _GEN_3923 : valid_815; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4950 = _array_io_en_T_1 ? _GEN_3924 : valid_816; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4951 = _array_io_en_T_1 ? _GEN_3925 : valid_817; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4952 = _array_io_en_T_1 ? _GEN_3926 : valid_818; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4953 = _array_io_en_T_1 ? _GEN_3927 : valid_819; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4954 = _array_io_en_T_1 ? _GEN_3928 : valid_820; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4955 = _array_io_en_T_1 ? _GEN_3929 : valid_821; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4956 = _array_io_en_T_1 ? _GEN_3930 : valid_822; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4957 = _array_io_en_T_1 ? _GEN_3931 : valid_823; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4958 = _array_io_en_T_1 ? _GEN_3932 : valid_824; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4959 = _array_io_en_T_1 ? _GEN_3933 : valid_825; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4960 = _array_io_en_T_1 ? _GEN_3934 : valid_826; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4961 = _array_io_en_T_1 ? _GEN_3935 : valid_827; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4962 = _array_io_en_T_1 ? _GEN_3936 : valid_828; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4963 = _array_io_en_T_1 ? _GEN_3937 : valid_829; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4964 = _array_io_en_T_1 ? _GEN_3938 : valid_830; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4965 = _array_io_en_T_1 ? _GEN_3939 : valid_831; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4966 = _array_io_en_T_1 ? _GEN_3940 : valid_832; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4967 = _array_io_en_T_1 ? _GEN_3941 : valid_833; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4968 = _array_io_en_T_1 ? _GEN_3942 : valid_834; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4969 = _array_io_en_T_1 ? _GEN_3943 : valid_835; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4970 = _array_io_en_T_1 ? _GEN_3944 : valid_836; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4971 = _array_io_en_T_1 ? _GEN_3945 : valid_837; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4972 = _array_io_en_T_1 ? _GEN_3946 : valid_838; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4973 = _array_io_en_T_1 ? _GEN_3947 : valid_839; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4974 = _array_io_en_T_1 ? _GEN_3948 : valid_840; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4975 = _array_io_en_T_1 ? _GEN_3949 : valid_841; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4976 = _array_io_en_T_1 ? _GEN_3950 : valid_842; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4977 = _array_io_en_T_1 ? _GEN_3951 : valid_843; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4978 = _array_io_en_T_1 ? _GEN_3952 : valid_844; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4979 = _array_io_en_T_1 ? _GEN_3953 : valid_845; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4980 = _array_io_en_T_1 ? _GEN_3954 : valid_846; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4981 = _array_io_en_T_1 ? _GEN_3955 : valid_847; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4982 = _array_io_en_T_1 ? _GEN_3956 : valid_848; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4983 = _array_io_en_T_1 ? _GEN_3957 : valid_849; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4984 = _array_io_en_T_1 ? _GEN_3958 : valid_850; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4985 = _array_io_en_T_1 ? _GEN_3959 : valid_851; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4986 = _array_io_en_T_1 ? _GEN_3960 : valid_852; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4987 = _array_io_en_T_1 ? _GEN_3961 : valid_853; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4988 = _array_io_en_T_1 ? _GEN_3962 : valid_854; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4989 = _array_io_en_T_1 ? _GEN_3963 : valid_855; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4990 = _array_io_en_T_1 ? _GEN_3964 : valid_856; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4991 = _array_io_en_T_1 ? _GEN_3965 : valid_857; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4992 = _array_io_en_T_1 ? _GEN_3966 : valid_858; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4993 = _array_io_en_T_1 ? _GEN_3967 : valid_859; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4994 = _array_io_en_T_1 ? _GEN_3968 : valid_860; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4995 = _array_io_en_T_1 ? _GEN_3969 : valid_861; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4996 = _array_io_en_T_1 ? _GEN_3970 : valid_862; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4997 = _array_io_en_T_1 ? _GEN_3971 : valid_863; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4998 = _array_io_en_T_1 ? _GEN_3972 : valid_864; // @[DCache.scala 164:19 56:22]
  wire  _GEN_4999 = _array_io_en_T_1 ? _GEN_3973 : valid_865; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5000 = _array_io_en_T_1 ? _GEN_3974 : valid_866; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5001 = _array_io_en_T_1 ? _GEN_3975 : valid_867; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5002 = _array_io_en_T_1 ? _GEN_3976 : valid_868; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5003 = _array_io_en_T_1 ? _GEN_3977 : valid_869; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5004 = _array_io_en_T_1 ? _GEN_3978 : valid_870; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5005 = _array_io_en_T_1 ? _GEN_3979 : valid_871; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5006 = _array_io_en_T_1 ? _GEN_3980 : valid_872; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5007 = _array_io_en_T_1 ? _GEN_3981 : valid_873; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5008 = _array_io_en_T_1 ? _GEN_3982 : valid_874; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5009 = _array_io_en_T_1 ? _GEN_3983 : valid_875; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5010 = _array_io_en_T_1 ? _GEN_3984 : valid_876; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5011 = _array_io_en_T_1 ? _GEN_3985 : valid_877; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5012 = _array_io_en_T_1 ? _GEN_3986 : valid_878; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5013 = _array_io_en_T_1 ? _GEN_3987 : valid_879; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5014 = _array_io_en_T_1 ? _GEN_3988 : valid_880; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5015 = _array_io_en_T_1 ? _GEN_3989 : valid_881; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5016 = _array_io_en_T_1 ? _GEN_3990 : valid_882; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5017 = _array_io_en_T_1 ? _GEN_3991 : valid_883; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5018 = _array_io_en_T_1 ? _GEN_3992 : valid_884; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5019 = _array_io_en_T_1 ? _GEN_3993 : valid_885; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5020 = _array_io_en_T_1 ? _GEN_3994 : valid_886; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5021 = _array_io_en_T_1 ? _GEN_3995 : valid_887; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5022 = _array_io_en_T_1 ? _GEN_3996 : valid_888; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5023 = _array_io_en_T_1 ? _GEN_3997 : valid_889; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5024 = _array_io_en_T_1 ? _GEN_3998 : valid_890; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5025 = _array_io_en_T_1 ? _GEN_3999 : valid_891; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5026 = _array_io_en_T_1 ? _GEN_4000 : valid_892; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5027 = _array_io_en_T_1 ? _GEN_4001 : valid_893; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5028 = _array_io_en_T_1 ? _GEN_4002 : valid_894; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5029 = _array_io_en_T_1 ? _GEN_4003 : valid_895; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5030 = _array_io_en_T_1 ? _GEN_4004 : valid_896; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5031 = _array_io_en_T_1 ? _GEN_4005 : valid_897; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5032 = _array_io_en_T_1 ? _GEN_4006 : valid_898; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5033 = _array_io_en_T_1 ? _GEN_4007 : valid_899; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5034 = _array_io_en_T_1 ? _GEN_4008 : valid_900; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5035 = _array_io_en_T_1 ? _GEN_4009 : valid_901; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5036 = _array_io_en_T_1 ? _GEN_4010 : valid_902; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5037 = _array_io_en_T_1 ? _GEN_4011 : valid_903; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5038 = _array_io_en_T_1 ? _GEN_4012 : valid_904; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5039 = _array_io_en_T_1 ? _GEN_4013 : valid_905; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5040 = _array_io_en_T_1 ? _GEN_4014 : valid_906; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5041 = _array_io_en_T_1 ? _GEN_4015 : valid_907; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5042 = _array_io_en_T_1 ? _GEN_4016 : valid_908; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5043 = _array_io_en_T_1 ? _GEN_4017 : valid_909; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5044 = _array_io_en_T_1 ? _GEN_4018 : valid_910; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5045 = _array_io_en_T_1 ? _GEN_4019 : valid_911; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5046 = _array_io_en_T_1 ? _GEN_4020 : valid_912; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5047 = _array_io_en_T_1 ? _GEN_4021 : valid_913; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5048 = _array_io_en_T_1 ? _GEN_4022 : valid_914; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5049 = _array_io_en_T_1 ? _GEN_4023 : valid_915; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5050 = _array_io_en_T_1 ? _GEN_4024 : valid_916; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5051 = _array_io_en_T_1 ? _GEN_4025 : valid_917; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5052 = _array_io_en_T_1 ? _GEN_4026 : valid_918; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5053 = _array_io_en_T_1 ? _GEN_4027 : valid_919; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5054 = _array_io_en_T_1 ? _GEN_4028 : valid_920; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5055 = _array_io_en_T_1 ? _GEN_4029 : valid_921; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5056 = _array_io_en_T_1 ? _GEN_4030 : valid_922; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5057 = _array_io_en_T_1 ? _GEN_4031 : valid_923; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5058 = _array_io_en_T_1 ? _GEN_4032 : valid_924; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5059 = _array_io_en_T_1 ? _GEN_4033 : valid_925; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5060 = _array_io_en_T_1 ? _GEN_4034 : valid_926; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5061 = _array_io_en_T_1 ? _GEN_4035 : valid_927; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5062 = _array_io_en_T_1 ? _GEN_4036 : valid_928; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5063 = _array_io_en_T_1 ? _GEN_4037 : valid_929; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5064 = _array_io_en_T_1 ? _GEN_4038 : valid_930; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5065 = _array_io_en_T_1 ? _GEN_4039 : valid_931; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5066 = _array_io_en_T_1 ? _GEN_4040 : valid_932; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5067 = _array_io_en_T_1 ? _GEN_4041 : valid_933; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5068 = _array_io_en_T_1 ? _GEN_4042 : valid_934; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5069 = _array_io_en_T_1 ? _GEN_4043 : valid_935; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5070 = _array_io_en_T_1 ? _GEN_4044 : valid_936; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5071 = _array_io_en_T_1 ? _GEN_4045 : valid_937; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5072 = _array_io_en_T_1 ? _GEN_4046 : valid_938; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5073 = _array_io_en_T_1 ? _GEN_4047 : valid_939; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5074 = _array_io_en_T_1 ? _GEN_4048 : valid_940; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5075 = _array_io_en_T_1 ? _GEN_4049 : valid_941; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5076 = _array_io_en_T_1 ? _GEN_4050 : valid_942; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5077 = _array_io_en_T_1 ? _GEN_4051 : valid_943; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5078 = _array_io_en_T_1 ? _GEN_4052 : valid_944; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5079 = _array_io_en_T_1 ? _GEN_4053 : valid_945; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5080 = _array_io_en_T_1 ? _GEN_4054 : valid_946; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5081 = _array_io_en_T_1 ? _GEN_4055 : valid_947; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5082 = _array_io_en_T_1 ? _GEN_4056 : valid_948; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5083 = _array_io_en_T_1 ? _GEN_4057 : valid_949; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5084 = _array_io_en_T_1 ? _GEN_4058 : valid_950; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5085 = _array_io_en_T_1 ? _GEN_4059 : valid_951; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5086 = _array_io_en_T_1 ? _GEN_4060 : valid_952; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5087 = _array_io_en_T_1 ? _GEN_4061 : valid_953; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5088 = _array_io_en_T_1 ? _GEN_4062 : valid_954; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5089 = _array_io_en_T_1 ? _GEN_4063 : valid_955; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5090 = _array_io_en_T_1 ? _GEN_4064 : valid_956; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5091 = _array_io_en_T_1 ? _GEN_4065 : valid_957; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5092 = _array_io_en_T_1 ? _GEN_4066 : valid_958; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5093 = _array_io_en_T_1 ? _GEN_4067 : valid_959; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5094 = _array_io_en_T_1 ? _GEN_4068 : valid_960; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5095 = _array_io_en_T_1 ? _GEN_4069 : valid_961; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5096 = _array_io_en_T_1 ? _GEN_4070 : valid_962; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5097 = _array_io_en_T_1 ? _GEN_4071 : valid_963; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5098 = _array_io_en_T_1 ? _GEN_4072 : valid_964; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5099 = _array_io_en_T_1 ? _GEN_4073 : valid_965; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5100 = _array_io_en_T_1 ? _GEN_4074 : valid_966; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5101 = _array_io_en_T_1 ? _GEN_4075 : valid_967; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5102 = _array_io_en_T_1 ? _GEN_4076 : valid_968; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5103 = _array_io_en_T_1 ? _GEN_4077 : valid_969; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5104 = _array_io_en_T_1 ? _GEN_4078 : valid_970; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5105 = _array_io_en_T_1 ? _GEN_4079 : valid_971; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5106 = _array_io_en_T_1 ? _GEN_4080 : valid_972; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5107 = _array_io_en_T_1 ? _GEN_4081 : valid_973; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5108 = _array_io_en_T_1 ? _GEN_4082 : valid_974; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5109 = _array_io_en_T_1 ? _GEN_4083 : valid_975; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5110 = _array_io_en_T_1 ? _GEN_4084 : valid_976; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5111 = _array_io_en_T_1 ? _GEN_4085 : valid_977; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5112 = _array_io_en_T_1 ? _GEN_4086 : valid_978; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5113 = _array_io_en_T_1 ? _GEN_4087 : valid_979; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5114 = _array_io_en_T_1 ? _GEN_4088 : valid_980; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5115 = _array_io_en_T_1 ? _GEN_4089 : valid_981; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5116 = _array_io_en_T_1 ? _GEN_4090 : valid_982; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5117 = _array_io_en_T_1 ? _GEN_4091 : valid_983; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5118 = _array_io_en_T_1 ? _GEN_4092 : valid_984; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5119 = _array_io_en_T_1 ? _GEN_4093 : valid_985; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5120 = _array_io_en_T_1 ? _GEN_4094 : valid_986; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5121 = _array_io_en_T_1 ? _GEN_4095 : valid_987; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5122 = _array_io_en_T_1 ? _GEN_4096 : valid_988; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5123 = _array_io_en_T_1 ? _GEN_4097 : valid_989; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5124 = _array_io_en_T_1 ? _GEN_4098 : valid_990; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5125 = _array_io_en_T_1 ? _GEN_4099 : valid_991; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5126 = _array_io_en_T_1 ? _GEN_4100 : valid_992; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5127 = _array_io_en_T_1 ? _GEN_4101 : valid_993; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5128 = _array_io_en_T_1 ? _GEN_4102 : valid_994; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5129 = _array_io_en_T_1 ? _GEN_4103 : valid_995; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5130 = _array_io_en_T_1 ? _GEN_4104 : valid_996; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5131 = _array_io_en_T_1 ? _GEN_4105 : valid_997; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5132 = _array_io_en_T_1 ? _GEN_4106 : valid_998; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5133 = _array_io_en_T_1 ? _GEN_4107 : valid_999; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5134 = _array_io_en_T_1 ? _GEN_4108 : valid_1000; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5135 = _array_io_en_T_1 ? _GEN_4109 : valid_1001; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5136 = _array_io_en_T_1 ? _GEN_4110 : valid_1002; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5137 = _array_io_en_T_1 ? _GEN_4111 : valid_1003; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5138 = _array_io_en_T_1 ? _GEN_4112 : valid_1004; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5139 = _array_io_en_T_1 ? _GEN_4113 : valid_1005; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5140 = _array_io_en_T_1 ? _GEN_4114 : valid_1006; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5141 = _array_io_en_T_1 ? _GEN_4115 : valid_1007; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5142 = _array_io_en_T_1 ? _GEN_4116 : valid_1008; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5143 = _array_io_en_T_1 ? _GEN_4117 : valid_1009; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5144 = _array_io_en_T_1 ? _GEN_4118 : valid_1010; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5145 = _array_io_en_T_1 ? _GEN_4119 : valid_1011; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5146 = _array_io_en_T_1 ? _GEN_4120 : valid_1012; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5147 = _array_io_en_T_1 ? _GEN_4121 : valid_1013; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5148 = _array_io_en_T_1 ? _GEN_4122 : valid_1014; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5149 = _array_io_en_T_1 ? _GEN_4123 : valid_1015; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5150 = _array_io_en_T_1 ? _GEN_4124 : valid_1016; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5151 = _array_io_en_T_1 ? _GEN_4125 : valid_1017; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5152 = _array_io_en_T_1 ? _GEN_4126 : valid_1018; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5153 = _array_io_en_T_1 ? _GEN_4127 : valid_1019; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5154 = _array_io_en_T_1 ? _GEN_4128 : valid_1020; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5155 = _array_io_en_T_1 ? _GEN_4129 : valid_1021; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5156 = _array_io_en_T_1 ? _GEN_4130 : valid_1022; // @[DCache.scala 164:19 56:22]
  wire  _GEN_5157 = _array_io_en_T_1 ? _GEN_4131 : valid_1023; // @[DCache.scala 164:19 56:22]
  wire  tl_c_valid = probing | state == 3'h2 & _GEN_1047; // @[DCache.scala 260:25]
  wire  _probing_T_1 = auto_out_c_ready & tl_c_valid; // @[Decoupled.scala 51:35]
  wire  _GEN_5158 = _probing_T_1 ? 1'h0 : probing; // @[Utils.scala 38:18 36:20 38:22]
  wire  _GEN_5159 = _tl_b_bits_r_T | _GEN_5158; // @[Utils.scala 39:{19,23}]
  wire [2:0] _state_T_1 = _GEN_1047 ? 3'h2 : 3'h4; // @[DCache.scala 194:21]
  wire [2:0] _GEN_5161 = ~array_hit ? _state_T_1 : state; // @[DCache.scala 193:30 194:15 60:118]
  wire [2:0] _GEN_5163 = _probing_T_1 & _x1_b_ready_T ? 3'h3 : state; // @[DCache.scala 200:41 201:15 60:118]
  wire [2:0] _GEN_5164 = ~_GEN_1047 ? 3'h4 : _GEN_5163; // @[DCache.scala 198:26 199:15]
  wire [2:0] _GEN_5165 = _tl_d_bits_r_T ? 3'h4 : state; // @[DCache.scala 205:23 206:15 60:118]
  wire  tl_a_valid = state == 3'h4; // @[DCache.scala 257:24]
  wire  _T_27 = auto_out_a_ready & tl_a_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_5166 = _T_27 ? 3'h5 : state; // @[DCache.scala 210:23 211:15 60:118]
  wire [2:0] _GEN_5167 = _tl_d_bits_r_T ? 3'h6 : state; // @[DCache.scala 215:23 216:15 60:118]
  wire  tl_e_valid = state == 3'h6; // @[DCache.scala 263:24]
  wire  _T_31 = auto_out_e_ready & tl_e_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_5168 = _T_31 ? 3'h7 : state; // @[DCache.scala 220:23 221:15 60:118]
  wire [2:0] _GEN_5169 = _array_io_en_T_1 ? 3'h0 : state; // @[DCache.scala 225:23 226:15 60:118]
  wire [2:0] _GEN_5170 = 3'h7 == state ? _GEN_5169 : state; // @[DCache.scala 184:17 60:118]
  wire [2:0] _GEN_5171 = 3'h6 == state ? _GEN_5168 : _GEN_5170; // @[DCache.scala 184:17]
  wire [2:0] _GEN_5172 = 3'h5 == state ? _GEN_5167 : _GEN_5171; // @[DCache.scala 184:17]
  wire [2:0] _GEN_5173 = 3'h4 == state ? _GEN_5166 : _GEN_5172; // @[DCache.scala 184:17]
  wire [2:0] _GEN_5174 = 3'h3 == state ? _GEN_5165 : _GEN_5173; // @[DCache.scala 184:17]
  reg  probe_out_REG; // @[DCache.scala 233:54]
  reg [272:0] probe_out_r; // @[Reg.scala 35:20]
  wire [272:0] _GEN_5178 = probe_out_REG ? array_io_rdata : probe_out_r; // @[Reg.scala 36:18 35:20 36:22]
  wire [255:0] probe_out_data = _GEN_5178[255:0]; // @[DCache.scala 233:75]
  wire [16:0] probe_out_tag = _GEN_5178[272:256]; // @[DCache.scala 233:75]
  wire  _GEN_5180 = 10'h1 == _GEN_4[14:5] ? valid_1 : valid_0; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5181 = 10'h2 == _GEN_4[14:5] ? valid_2 : _GEN_5180; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5182 = 10'h3 == _GEN_4[14:5] ? valid_3 : _GEN_5181; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5183 = 10'h4 == _GEN_4[14:5] ? valid_4 : _GEN_5182; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5184 = 10'h5 == _GEN_4[14:5] ? valid_5 : _GEN_5183; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5185 = 10'h6 == _GEN_4[14:5] ? valid_6 : _GEN_5184; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5186 = 10'h7 == _GEN_4[14:5] ? valid_7 : _GEN_5185; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5187 = 10'h8 == _GEN_4[14:5] ? valid_8 : _GEN_5186; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5188 = 10'h9 == _GEN_4[14:5] ? valid_9 : _GEN_5187; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5189 = 10'ha == _GEN_4[14:5] ? valid_10 : _GEN_5188; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5190 = 10'hb == _GEN_4[14:5] ? valid_11 : _GEN_5189; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5191 = 10'hc == _GEN_4[14:5] ? valid_12 : _GEN_5190; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5192 = 10'hd == _GEN_4[14:5] ? valid_13 : _GEN_5191; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5193 = 10'he == _GEN_4[14:5] ? valid_14 : _GEN_5192; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5194 = 10'hf == _GEN_4[14:5] ? valid_15 : _GEN_5193; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5195 = 10'h10 == _GEN_4[14:5] ? valid_16 : _GEN_5194; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5196 = 10'h11 == _GEN_4[14:5] ? valid_17 : _GEN_5195; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5197 = 10'h12 == _GEN_4[14:5] ? valid_18 : _GEN_5196; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5198 = 10'h13 == _GEN_4[14:5] ? valid_19 : _GEN_5197; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5199 = 10'h14 == _GEN_4[14:5] ? valid_20 : _GEN_5198; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5200 = 10'h15 == _GEN_4[14:5] ? valid_21 : _GEN_5199; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5201 = 10'h16 == _GEN_4[14:5] ? valid_22 : _GEN_5200; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5202 = 10'h17 == _GEN_4[14:5] ? valid_23 : _GEN_5201; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5203 = 10'h18 == _GEN_4[14:5] ? valid_24 : _GEN_5202; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5204 = 10'h19 == _GEN_4[14:5] ? valid_25 : _GEN_5203; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5205 = 10'h1a == _GEN_4[14:5] ? valid_26 : _GEN_5204; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5206 = 10'h1b == _GEN_4[14:5] ? valid_27 : _GEN_5205; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5207 = 10'h1c == _GEN_4[14:5] ? valid_28 : _GEN_5206; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5208 = 10'h1d == _GEN_4[14:5] ? valid_29 : _GEN_5207; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5209 = 10'h1e == _GEN_4[14:5] ? valid_30 : _GEN_5208; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5210 = 10'h1f == _GEN_4[14:5] ? valid_31 : _GEN_5209; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5211 = 10'h20 == _GEN_4[14:5] ? valid_32 : _GEN_5210; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5212 = 10'h21 == _GEN_4[14:5] ? valid_33 : _GEN_5211; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5213 = 10'h22 == _GEN_4[14:5] ? valid_34 : _GEN_5212; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5214 = 10'h23 == _GEN_4[14:5] ? valid_35 : _GEN_5213; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5215 = 10'h24 == _GEN_4[14:5] ? valid_36 : _GEN_5214; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5216 = 10'h25 == _GEN_4[14:5] ? valid_37 : _GEN_5215; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5217 = 10'h26 == _GEN_4[14:5] ? valid_38 : _GEN_5216; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5218 = 10'h27 == _GEN_4[14:5] ? valid_39 : _GEN_5217; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5219 = 10'h28 == _GEN_4[14:5] ? valid_40 : _GEN_5218; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5220 = 10'h29 == _GEN_4[14:5] ? valid_41 : _GEN_5219; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5221 = 10'h2a == _GEN_4[14:5] ? valid_42 : _GEN_5220; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5222 = 10'h2b == _GEN_4[14:5] ? valid_43 : _GEN_5221; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5223 = 10'h2c == _GEN_4[14:5] ? valid_44 : _GEN_5222; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5224 = 10'h2d == _GEN_4[14:5] ? valid_45 : _GEN_5223; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5225 = 10'h2e == _GEN_4[14:5] ? valid_46 : _GEN_5224; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5226 = 10'h2f == _GEN_4[14:5] ? valid_47 : _GEN_5225; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5227 = 10'h30 == _GEN_4[14:5] ? valid_48 : _GEN_5226; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5228 = 10'h31 == _GEN_4[14:5] ? valid_49 : _GEN_5227; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5229 = 10'h32 == _GEN_4[14:5] ? valid_50 : _GEN_5228; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5230 = 10'h33 == _GEN_4[14:5] ? valid_51 : _GEN_5229; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5231 = 10'h34 == _GEN_4[14:5] ? valid_52 : _GEN_5230; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5232 = 10'h35 == _GEN_4[14:5] ? valid_53 : _GEN_5231; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5233 = 10'h36 == _GEN_4[14:5] ? valid_54 : _GEN_5232; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5234 = 10'h37 == _GEN_4[14:5] ? valid_55 : _GEN_5233; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5235 = 10'h38 == _GEN_4[14:5] ? valid_56 : _GEN_5234; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5236 = 10'h39 == _GEN_4[14:5] ? valid_57 : _GEN_5235; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5237 = 10'h3a == _GEN_4[14:5] ? valid_58 : _GEN_5236; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5238 = 10'h3b == _GEN_4[14:5] ? valid_59 : _GEN_5237; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5239 = 10'h3c == _GEN_4[14:5] ? valid_60 : _GEN_5238; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5240 = 10'h3d == _GEN_4[14:5] ? valid_61 : _GEN_5239; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5241 = 10'h3e == _GEN_4[14:5] ? valid_62 : _GEN_5240; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5242 = 10'h3f == _GEN_4[14:5] ? valid_63 : _GEN_5241; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5243 = 10'h40 == _GEN_4[14:5] ? valid_64 : _GEN_5242; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5244 = 10'h41 == _GEN_4[14:5] ? valid_65 : _GEN_5243; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5245 = 10'h42 == _GEN_4[14:5] ? valid_66 : _GEN_5244; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5246 = 10'h43 == _GEN_4[14:5] ? valid_67 : _GEN_5245; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5247 = 10'h44 == _GEN_4[14:5] ? valid_68 : _GEN_5246; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5248 = 10'h45 == _GEN_4[14:5] ? valid_69 : _GEN_5247; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5249 = 10'h46 == _GEN_4[14:5] ? valid_70 : _GEN_5248; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5250 = 10'h47 == _GEN_4[14:5] ? valid_71 : _GEN_5249; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5251 = 10'h48 == _GEN_4[14:5] ? valid_72 : _GEN_5250; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5252 = 10'h49 == _GEN_4[14:5] ? valid_73 : _GEN_5251; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5253 = 10'h4a == _GEN_4[14:5] ? valid_74 : _GEN_5252; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5254 = 10'h4b == _GEN_4[14:5] ? valid_75 : _GEN_5253; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5255 = 10'h4c == _GEN_4[14:5] ? valid_76 : _GEN_5254; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5256 = 10'h4d == _GEN_4[14:5] ? valid_77 : _GEN_5255; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5257 = 10'h4e == _GEN_4[14:5] ? valid_78 : _GEN_5256; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5258 = 10'h4f == _GEN_4[14:5] ? valid_79 : _GEN_5257; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5259 = 10'h50 == _GEN_4[14:5] ? valid_80 : _GEN_5258; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5260 = 10'h51 == _GEN_4[14:5] ? valid_81 : _GEN_5259; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5261 = 10'h52 == _GEN_4[14:5] ? valid_82 : _GEN_5260; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5262 = 10'h53 == _GEN_4[14:5] ? valid_83 : _GEN_5261; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5263 = 10'h54 == _GEN_4[14:5] ? valid_84 : _GEN_5262; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5264 = 10'h55 == _GEN_4[14:5] ? valid_85 : _GEN_5263; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5265 = 10'h56 == _GEN_4[14:5] ? valid_86 : _GEN_5264; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5266 = 10'h57 == _GEN_4[14:5] ? valid_87 : _GEN_5265; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5267 = 10'h58 == _GEN_4[14:5] ? valid_88 : _GEN_5266; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5268 = 10'h59 == _GEN_4[14:5] ? valid_89 : _GEN_5267; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5269 = 10'h5a == _GEN_4[14:5] ? valid_90 : _GEN_5268; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5270 = 10'h5b == _GEN_4[14:5] ? valid_91 : _GEN_5269; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5271 = 10'h5c == _GEN_4[14:5] ? valid_92 : _GEN_5270; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5272 = 10'h5d == _GEN_4[14:5] ? valid_93 : _GEN_5271; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5273 = 10'h5e == _GEN_4[14:5] ? valid_94 : _GEN_5272; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5274 = 10'h5f == _GEN_4[14:5] ? valid_95 : _GEN_5273; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5275 = 10'h60 == _GEN_4[14:5] ? valid_96 : _GEN_5274; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5276 = 10'h61 == _GEN_4[14:5] ? valid_97 : _GEN_5275; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5277 = 10'h62 == _GEN_4[14:5] ? valid_98 : _GEN_5276; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5278 = 10'h63 == _GEN_4[14:5] ? valid_99 : _GEN_5277; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5279 = 10'h64 == _GEN_4[14:5] ? valid_100 : _GEN_5278; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5280 = 10'h65 == _GEN_4[14:5] ? valid_101 : _GEN_5279; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5281 = 10'h66 == _GEN_4[14:5] ? valid_102 : _GEN_5280; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5282 = 10'h67 == _GEN_4[14:5] ? valid_103 : _GEN_5281; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5283 = 10'h68 == _GEN_4[14:5] ? valid_104 : _GEN_5282; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5284 = 10'h69 == _GEN_4[14:5] ? valid_105 : _GEN_5283; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5285 = 10'h6a == _GEN_4[14:5] ? valid_106 : _GEN_5284; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5286 = 10'h6b == _GEN_4[14:5] ? valid_107 : _GEN_5285; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5287 = 10'h6c == _GEN_4[14:5] ? valid_108 : _GEN_5286; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5288 = 10'h6d == _GEN_4[14:5] ? valid_109 : _GEN_5287; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5289 = 10'h6e == _GEN_4[14:5] ? valid_110 : _GEN_5288; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5290 = 10'h6f == _GEN_4[14:5] ? valid_111 : _GEN_5289; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5291 = 10'h70 == _GEN_4[14:5] ? valid_112 : _GEN_5290; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5292 = 10'h71 == _GEN_4[14:5] ? valid_113 : _GEN_5291; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5293 = 10'h72 == _GEN_4[14:5] ? valid_114 : _GEN_5292; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5294 = 10'h73 == _GEN_4[14:5] ? valid_115 : _GEN_5293; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5295 = 10'h74 == _GEN_4[14:5] ? valid_116 : _GEN_5294; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5296 = 10'h75 == _GEN_4[14:5] ? valid_117 : _GEN_5295; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5297 = 10'h76 == _GEN_4[14:5] ? valid_118 : _GEN_5296; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5298 = 10'h77 == _GEN_4[14:5] ? valid_119 : _GEN_5297; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5299 = 10'h78 == _GEN_4[14:5] ? valid_120 : _GEN_5298; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5300 = 10'h79 == _GEN_4[14:5] ? valid_121 : _GEN_5299; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5301 = 10'h7a == _GEN_4[14:5] ? valid_122 : _GEN_5300; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5302 = 10'h7b == _GEN_4[14:5] ? valid_123 : _GEN_5301; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5303 = 10'h7c == _GEN_4[14:5] ? valid_124 : _GEN_5302; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5304 = 10'h7d == _GEN_4[14:5] ? valid_125 : _GEN_5303; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5305 = 10'h7e == _GEN_4[14:5] ? valid_126 : _GEN_5304; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5306 = 10'h7f == _GEN_4[14:5] ? valid_127 : _GEN_5305; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5307 = 10'h80 == _GEN_4[14:5] ? valid_128 : _GEN_5306; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5308 = 10'h81 == _GEN_4[14:5] ? valid_129 : _GEN_5307; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5309 = 10'h82 == _GEN_4[14:5] ? valid_130 : _GEN_5308; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5310 = 10'h83 == _GEN_4[14:5] ? valid_131 : _GEN_5309; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5311 = 10'h84 == _GEN_4[14:5] ? valid_132 : _GEN_5310; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5312 = 10'h85 == _GEN_4[14:5] ? valid_133 : _GEN_5311; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5313 = 10'h86 == _GEN_4[14:5] ? valid_134 : _GEN_5312; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5314 = 10'h87 == _GEN_4[14:5] ? valid_135 : _GEN_5313; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5315 = 10'h88 == _GEN_4[14:5] ? valid_136 : _GEN_5314; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5316 = 10'h89 == _GEN_4[14:5] ? valid_137 : _GEN_5315; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5317 = 10'h8a == _GEN_4[14:5] ? valid_138 : _GEN_5316; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5318 = 10'h8b == _GEN_4[14:5] ? valid_139 : _GEN_5317; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5319 = 10'h8c == _GEN_4[14:5] ? valid_140 : _GEN_5318; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5320 = 10'h8d == _GEN_4[14:5] ? valid_141 : _GEN_5319; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5321 = 10'h8e == _GEN_4[14:5] ? valid_142 : _GEN_5320; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5322 = 10'h8f == _GEN_4[14:5] ? valid_143 : _GEN_5321; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5323 = 10'h90 == _GEN_4[14:5] ? valid_144 : _GEN_5322; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5324 = 10'h91 == _GEN_4[14:5] ? valid_145 : _GEN_5323; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5325 = 10'h92 == _GEN_4[14:5] ? valid_146 : _GEN_5324; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5326 = 10'h93 == _GEN_4[14:5] ? valid_147 : _GEN_5325; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5327 = 10'h94 == _GEN_4[14:5] ? valid_148 : _GEN_5326; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5328 = 10'h95 == _GEN_4[14:5] ? valid_149 : _GEN_5327; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5329 = 10'h96 == _GEN_4[14:5] ? valid_150 : _GEN_5328; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5330 = 10'h97 == _GEN_4[14:5] ? valid_151 : _GEN_5329; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5331 = 10'h98 == _GEN_4[14:5] ? valid_152 : _GEN_5330; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5332 = 10'h99 == _GEN_4[14:5] ? valid_153 : _GEN_5331; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5333 = 10'h9a == _GEN_4[14:5] ? valid_154 : _GEN_5332; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5334 = 10'h9b == _GEN_4[14:5] ? valid_155 : _GEN_5333; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5335 = 10'h9c == _GEN_4[14:5] ? valid_156 : _GEN_5334; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5336 = 10'h9d == _GEN_4[14:5] ? valid_157 : _GEN_5335; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5337 = 10'h9e == _GEN_4[14:5] ? valid_158 : _GEN_5336; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5338 = 10'h9f == _GEN_4[14:5] ? valid_159 : _GEN_5337; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5339 = 10'ha0 == _GEN_4[14:5] ? valid_160 : _GEN_5338; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5340 = 10'ha1 == _GEN_4[14:5] ? valid_161 : _GEN_5339; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5341 = 10'ha2 == _GEN_4[14:5] ? valid_162 : _GEN_5340; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5342 = 10'ha3 == _GEN_4[14:5] ? valid_163 : _GEN_5341; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5343 = 10'ha4 == _GEN_4[14:5] ? valid_164 : _GEN_5342; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5344 = 10'ha5 == _GEN_4[14:5] ? valid_165 : _GEN_5343; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5345 = 10'ha6 == _GEN_4[14:5] ? valid_166 : _GEN_5344; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5346 = 10'ha7 == _GEN_4[14:5] ? valid_167 : _GEN_5345; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5347 = 10'ha8 == _GEN_4[14:5] ? valid_168 : _GEN_5346; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5348 = 10'ha9 == _GEN_4[14:5] ? valid_169 : _GEN_5347; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5349 = 10'haa == _GEN_4[14:5] ? valid_170 : _GEN_5348; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5350 = 10'hab == _GEN_4[14:5] ? valid_171 : _GEN_5349; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5351 = 10'hac == _GEN_4[14:5] ? valid_172 : _GEN_5350; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5352 = 10'had == _GEN_4[14:5] ? valid_173 : _GEN_5351; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5353 = 10'hae == _GEN_4[14:5] ? valid_174 : _GEN_5352; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5354 = 10'haf == _GEN_4[14:5] ? valid_175 : _GEN_5353; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5355 = 10'hb0 == _GEN_4[14:5] ? valid_176 : _GEN_5354; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5356 = 10'hb1 == _GEN_4[14:5] ? valid_177 : _GEN_5355; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5357 = 10'hb2 == _GEN_4[14:5] ? valid_178 : _GEN_5356; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5358 = 10'hb3 == _GEN_4[14:5] ? valid_179 : _GEN_5357; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5359 = 10'hb4 == _GEN_4[14:5] ? valid_180 : _GEN_5358; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5360 = 10'hb5 == _GEN_4[14:5] ? valid_181 : _GEN_5359; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5361 = 10'hb6 == _GEN_4[14:5] ? valid_182 : _GEN_5360; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5362 = 10'hb7 == _GEN_4[14:5] ? valid_183 : _GEN_5361; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5363 = 10'hb8 == _GEN_4[14:5] ? valid_184 : _GEN_5362; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5364 = 10'hb9 == _GEN_4[14:5] ? valid_185 : _GEN_5363; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5365 = 10'hba == _GEN_4[14:5] ? valid_186 : _GEN_5364; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5366 = 10'hbb == _GEN_4[14:5] ? valid_187 : _GEN_5365; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5367 = 10'hbc == _GEN_4[14:5] ? valid_188 : _GEN_5366; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5368 = 10'hbd == _GEN_4[14:5] ? valid_189 : _GEN_5367; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5369 = 10'hbe == _GEN_4[14:5] ? valid_190 : _GEN_5368; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5370 = 10'hbf == _GEN_4[14:5] ? valid_191 : _GEN_5369; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5371 = 10'hc0 == _GEN_4[14:5] ? valid_192 : _GEN_5370; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5372 = 10'hc1 == _GEN_4[14:5] ? valid_193 : _GEN_5371; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5373 = 10'hc2 == _GEN_4[14:5] ? valid_194 : _GEN_5372; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5374 = 10'hc3 == _GEN_4[14:5] ? valid_195 : _GEN_5373; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5375 = 10'hc4 == _GEN_4[14:5] ? valid_196 : _GEN_5374; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5376 = 10'hc5 == _GEN_4[14:5] ? valid_197 : _GEN_5375; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5377 = 10'hc6 == _GEN_4[14:5] ? valid_198 : _GEN_5376; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5378 = 10'hc7 == _GEN_4[14:5] ? valid_199 : _GEN_5377; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5379 = 10'hc8 == _GEN_4[14:5] ? valid_200 : _GEN_5378; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5380 = 10'hc9 == _GEN_4[14:5] ? valid_201 : _GEN_5379; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5381 = 10'hca == _GEN_4[14:5] ? valid_202 : _GEN_5380; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5382 = 10'hcb == _GEN_4[14:5] ? valid_203 : _GEN_5381; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5383 = 10'hcc == _GEN_4[14:5] ? valid_204 : _GEN_5382; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5384 = 10'hcd == _GEN_4[14:5] ? valid_205 : _GEN_5383; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5385 = 10'hce == _GEN_4[14:5] ? valid_206 : _GEN_5384; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5386 = 10'hcf == _GEN_4[14:5] ? valid_207 : _GEN_5385; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5387 = 10'hd0 == _GEN_4[14:5] ? valid_208 : _GEN_5386; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5388 = 10'hd1 == _GEN_4[14:5] ? valid_209 : _GEN_5387; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5389 = 10'hd2 == _GEN_4[14:5] ? valid_210 : _GEN_5388; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5390 = 10'hd3 == _GEN_4[14:5] ? valid_211 : _GEN_5389; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5391 = 10'hd4 == _GEN_4[14:5] ? valid_212 : _GEN_5390; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5392 = 10'hd5 == _GEN_4[14:5] ? valid_213 : _GEN_5391; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5393 = 10'hd6 == _GEN_4[14:5] ? valid_214 : _GEN_5392; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5394 = 10'hd7 == _GEN_4[14:5] ? valid_215 : _GEN_5393; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5395 = 10'hd8 == _GEN_4[14:5] ? valid_216 : _GEN_5394; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5396 = 10'hd9 == _GEN_4[14:5] ? valid_217 : _GEN_5395; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5397 = 10'hda == _GEN_4[14:5] ? valid_218 : _GEN_5396; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5398 = 10'hdb == _GEN_4[14:5] ? valid_219 : _GEN_5397; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5399 = 10'hdc == _GEN_4[14:5] ? valid_220 : _GEN_5398; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5400 = 10'hdd == _GEN_4[14:5] ? valid_221 : _GEN_5399; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5401 = 10'hde == _GEN_4[14:5] ? valid_222 : _GEN_5400; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5402 = 10'hdf == _GEN_4[14:5] ? valid_223 : _GEN_5401; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5403 = 10'he0 == _GEN_4[14:5] ? valid_224 : _GEN_5402; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5404 = 10'he1 == _GEN_4[14:5] ? valid_225 : _GEN_5403; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5405 = 10'he2 == _GEN_4[14:5] ? valid_226 : _GEN_5404; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5406 = 10'he3 == _GEN_4[14:5] ? valid_227 : _GEN_5405; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5407 = 10'he4 == _GEN_4[14:5] ? valid_228 : _GEN_5406; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5408 = 10'he5 == _GEN_4[14:5] ? valid_229 : _GEN_5407; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5409 = 10'he6 == _GEN_4[14:5] ? valid_230 : _GEN_5408; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5410 = 10'he7 == _GEN_4[14:5] ? valid_231 : _GEN_5409; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5411 = 10'he8 == _GEN_4[14:5] ? valid_232 : _GEN_5410; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5412 = 10'he9 == _GEN_4[14:5] ? valid_233 : _GEN_5411; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5413 = 10'hea == _GEN_4[14:5] ? valid_234 : _GEN_5412; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5414 = 10'heb == _GEN_4[14:5] ? valid_235 : _GEN_5413; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5415 = 10'hec == _GEN_4[14:5] ? valid_236 : _GEN_5414; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5416 = 10'hed == _GEN_4[14:5] ? valid_237 : _GEN_5415; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5417 = 10'hee == _GEN_4[14:5] ? valid_238 : _GEN_5416; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5418 = 10'hef == _GEN_4[14:5] ? valid_239 : _GEN_5417; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5419 = 10'hf0 == _GEN_4[14:5] ? valid_240 : _GEN_5418; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5420 = 10'hf1 == _GEN_4[14:5] ? valid_241 : _GEN_5419; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5421 = 10'hf2 == _GEN_4[14:5] ? valid_242 : _GEN_5420; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5422 = 10'hf3 == _GEN_4[14:5] ? valid_243 : _GEN_5421; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5423 = 10'hf4 == _GEN_4[14:5] ? valid_244 : _GEN_5422; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5424 = 10'hf5 == _GEN_4[14:5] ? valid_245 : _GEN_5423; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5425 = 10'hf6 == _GEN_4[14:5] ? valid_246 : _GEN_5424; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5426 = 10'hf7 == _GEN_4[14:5] ? valid_247 : _GEN_5425; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5427 = 10'hf8 == _GEN_4[14:5] ? valid_248 : _GEN_5426; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5428 = 10'hf9 == _GEN_4[14:5] ? valid_249 : _GEN_5427; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5429 = 10'hfa == _GEN_4[14:5] ? valid_250 : _GEN_5428; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5430 = 10'hfb == _GEN_4[14:5] ? valid_251 : _GEN_5429; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5431 = 10'hfc == _GEN_4[14:5] ? valid_252 : _GEN_5430; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5432 = 10'hfd == _GEN_4[14:5] ? valid_253 : _GEN_5431; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5433 = 10'hfe == _GEN_4[14:5] ? valid_254 : _GEN_5432; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5434 = 10'hff == _GEN_4[14:5] ? valid_255 : _GEN_5433; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5435 = 10'h100 == _GEN_4[14:5] ? valid_256 : _GEN_5434; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5436 = 10'h101 == _GEN_4[14:5] ? valid_257 : _GEN_5435; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5437 = 10'h102 == _GEN_4[14:5] ? valid_258 : _GEN_5436; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5438 = 10'h103 == _GEN_4[14:5] ? valid_259 : _GEN_5437; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5439 = 10'h104 == _GEN_4[14:5] ? valid_260 : _GEN_5438; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5440 = 10'h105 == _GEN_4[14:5] ? valid_261 : _GEN_5439; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5441 = 10'h106 == _GEN_4[14:5] ? valid_262 : _GEN_5440; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5442 = 10'h107 == _GEN_4[14:5] ? valid_263 : _GEN_5441; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5443 = 10'h108 == _GEN_4[14:5] ? valid_264 : _GEN_5442; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5444 = 10'h109 == _GEN_4[14:5] ? valid_265 : _GEN_5443; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5445 = 10'h10a == _GEN_4[14:5] ? valid_266 : _GEN_5444; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5446 = 10'h10b == _GEN_4[14:5] ? valid_267 : _GEN_5445; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5447 = 10'h10c == _GEN_4[14:5] ? valid_268 : _GEN_5446; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5448 = 10'h10d == _GEN_4[14:5] ? valid_269 : _GEN_5447; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5449 = 10'h10e == _GEN_4[14:5] ? valid_270 : _GEN_5448; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5450 = 10'h10f == _GEN_4[14:5] ? valid_271 : _GEN_5449; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5451 = 10'h110 == _GEN_4[14:5] ? valid_272 : _GEN_5450; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5452 = 10'h111 == _GEN_4[14:5] ? valid_273 : _GEN_5451; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5453 = 10'h112 == _GEN_4[14:5] ? valid_274 : _GEN_5452; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5454 = 10'h113 == _GEN_4[14:5] ? valid_275 : _GEN_5453; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5455 = 10'h114 == _GEN_4[14:5] ? valid_276 : _GEN_5454; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5456 = 10'h115 == _GEN_4[14:5] ? valid_277 : _GEN_5455; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5457 = 10'h116 == _GEN_4[14:5] ? valid_278 : _GEN_5456; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5458 = 10'h117 == _GEN_4[14:5] ? valid_279 : _GEN_5457; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5459 = 10'h118 == _GEN_4[14:5] ? valid_280 : _GEN_5458; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5460 = 10'h119 == _GEN_4[14:5] ? valid_281 : _GEN_5459; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5461 = 10'h11a == _GEN_4[14:5] ? valid_282 : _GEN_5460; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5462 = 10'h11b == _GEN_4[14:5] ? valid_283 : _GEN_5461; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5463 = 10'h11c == _GEN_4[14:5] ? valid_284 : _GEN_5462; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5464 = 10'h11d == _GEN_4[14:5] ? valid_285 : _GEN_5463; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5465 = 10'h11e == _GEN_4[14:5] ? valid_286 : _GEN_5464; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5466 = 10'h11f == _GEN_4[14:5] ? valid_287 : _GEN_5465; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5467 = 10'h120 == _GEN_4[14:5] ? valid_288 : _GEN_5466; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5468 = 10'h121 == _GEN_4[14:5] ? valid_289 : _GEN_5467; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5469 = 10'h122 == _GEN_4[14:5] ? valid_290 : _GEN_5468; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5470 = 10'h123 == _GEN_4[14:5] ? valid_291 : _GEN_5469; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5471 = 10'h124 == _GEN_4[14:5] ? valid_292 : _GEN_5470; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5472 = 10'h125 == _GEN_4[14:5] ? valid_293 : _GEN_5471; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5473 = 10'h126 == _GEN_4[14:5] ? valid_294 : _GEN_5472; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5474 = 10'h127 == _GEN_4[14:5] ? valid_295 : _GEN_5473; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5475 = 10'h128 == _GEN_4[14:5] ? valid_296 : _GEN_5474; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5476 = 10'h129 == _GEN_4[14:5] ? valid_297 : _GEN_5475; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5477 = 10'h12a == _GEN_4[14:5] ? valid_298 : _GEN_5476; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5478 = 10'h12b == _GEN_4[14:5] ? valid_299 : _GEN_5477; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5479 = 10'h12c == _GEN_4[14:5] ? valid_300 : _GEN_5478; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5480 = 10'h12d == _GEN_4[14:5] ? valid_301 : _GEN_5479; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5481 = 10'h12e == _GEN_4[14:5] ? valid_302 : _GEN_5480; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5482 = 10'h12f == _GEN_4[14:5] ? valid_303 : _GEN_5481; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5483 = 10'h130 == _GEN_4[14:5] ? valid_304 : _GEN_5482; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5484 = 10'h131 == _GEN_4[14:5] ? valid_305 : _GEN_5483; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5485 = 10'h132 == _GEN_4[14:5] ? valid_306 : _GEN_5484; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5486 = 10'h133 == _GEN_4[14:5] ? valid_307 : _GEN_5485; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5487 = 10'h134 == _GEN_4[14:5] ? valid_308 : _GEN_5486; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5488 = 10'h135 == _GEN_4[14:5] ? valid_309 : _GEN_5487; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5489 = 10'h136 == _GEN_4[14:5] ? valid_310 : _GEN_5488; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5490 = 10'h137 == _GEN_4[14:5] ? valid_311 : _GEN_5489; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5491 = 10'h138 == _GEN_4[14:5] ? valid_312 : _GEN_5490; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5492 = 10'h139 == _GEN_4[14:5] ? valid_313 : _GEN_5491; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5493 = 10'h13a == _GEN_4[14:5] ? valid_314 : _GEN_5492; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5494 = 10'h13b == _GEN_4[14:5] ? valid_315 : _GEN_5493; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5495 = 10'h13c == _GEN_4[14:5] ? valid_316 : _GEN_5494; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5496 = 10'h13d == _GEN_4[14:5] ? valid_317 : _GEN_5495; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5497 = 10'h13e == _GEN_4[14:5] ? valid_318 : _GEN_5496; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5498 = 10'h13f == _GEN_4[14:5] ? valid_319 : _GEN_5497; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5499 = 10'h140 == _GEN_4[14:5] ? valid_320 : _GEN_5498; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5500 = 10'h141 == _GEN_4[14:5] ? valid_321 : _GEN_5499; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5501 = 10'h142 == _GEN_4[14:5] ? valid_322 : _GEN_5500; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5502 = 10'h143 == _GEN_4[14:5] ? valid_323 : _GEN_5501; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5503 = 10'h144 == _GEN_4[14:5] ? valid_324 : _GEN_5502; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5504 = 10'h145 == _GEN_4[14:5] ? valid_325 : _GEN_5503; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5505 = 10'h146 == _GEN_4[14:5] ? valid_326 : _GEN_5504; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5506 = 10'h147 == _GEN_4[14:5] ? valid_327 : _GEN_5505; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5507 = 10'h148 == _GEN_4[14:5] ? valid_328 : _GEN_5506; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5508 = 10'h149 == _GEN_4[14:5] ? valid_329 : _GEN_5507; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5509 = 10'h14a == _GEN_4[14:5] ? valid_330 : _GEN_5508; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5510 = 10'h14b == _GEN_4[14:5] ? valid_331 : _GEN_5509; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5511 = 10'h14c == _GEN_4[14:5] ? valid_332 : _GEN_5510; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5512 = 10'h14d == _GEN_4[14:5] ? valid_333 : _GEN_5511; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5513 = 10'h14e == _GEN_4[14:5] ? valid_334 : _GEN_5512; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5514 = 10'h14f == _GEN_4[14:5] ? valid_335 : _GEN_5513; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5515 = 10'h150 == _GEN_4[14:5] ? valid_336 : _GEN_5514; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5516 = 10'h151 == _GEN_4[14:5] ? valid_337 : _GEN_5515; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5517 = 10'h152 == _GEN_4[14:5] ? valid_338 : _GEN_5516; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5518 = 10'h153 == _GEN_4[14:5] ? valid_339 : _GEN_5517; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5519 = 10'h154 == _GEN_4[14:5] ? valid_340 : _GEN_5518; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5520 = 10'h155 == _GEN_4[14:5] ? valid_341 : _GEN_5519; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5521 = 10'h156 == _GEN_4[14:5] ? valid_342 : _GEN_5520; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5522 = 10'h157 == _GEN_4[14:5] ? valid_343 : _GEN_5521; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5523 = 10'h158 == _GEN_4[14:5] ? valid_344 : _GEN_5522; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5524 = 10'h159 == _GEN_4[14:5] ? valid_345 : _GEN_5523; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5525 = 10'h15a == _GEN_4[14:5] ? valid_346 : _GEN_5524; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5526 = 10'h15b == _GEN_4[14:5] ? valid_347 : _GEN_5525; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5527 = 10'h15c == _GEN_4[14:5] ? valid_348 : _GEN_5526; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5528 = 10'h15d == _GEN_4[14:5] ? valid_349 : _GEN_5527; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5529 = 10'h15e == _GEN_4[14:5] ? valid_350 : _GEN_5528; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5530 = 10'h15f == _GEN_4[14:5] ? valid_351 : _GEN_5529; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5531 = 10'h160 == _GEN_4[14:5] ? valid_352 : _GEN_5530; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5532 = 10'h161 == _GEN_4[14:5] ? valid_353 : _GEN_5531; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5533 = 10'h162 == _GEN_4[14:5] ? valid_354 : _GEN_5532; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5534 = 10'h163 == _GEN_4[14:5] ? valid_355 : _GEN_5533; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5535 = 10'h164 == _GEN_4[14:5] ? valid_356 : _GEN_5534; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5536 = 10'h165 == _GEN_4[14:5] ? valid_357 : _GEN_5535; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5537 = 10'h166 == _GEN_4[14:5] ? valid_358 : _GEN_5536; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5538 = 10'h167 == _GEN_4[14:5] ? valid_359 : _GEN_5537; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5539 = 10'h168 == _GEN_4[14:5] ? valid_360 : _GEN_5538; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5540 = 10'h169 == _GEN_4[14:5] ? valid_361 : _GEN_5539; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5541 = 10'h16a == _GEN_4[14:5] ? valid_362 : _GEN_5540; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5542 = 10'h16b == _GEN_4[14:5] ? valid_363 : _GEN_5541; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5543 = 10'h16c == _GEN_4[14:5] ? valid_364 : _GEN_5542; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5544 = 10'h16d == _GEN_4[14:5] ? valid_365 : _GEN_5543; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5545 = 10'h16e == _GEN_4[14:5] ? valid_366 : _GEN_5544; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5546 = 10'h16f == _GEN_4[14:5] ? valid_367 : _GEN_5545; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5547 = 10'h170 == _GEN_4[14:5] ? valid_368 : _GEN_5546; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5548 = 10'h171 == _GEN_4[14:5] ? valid_369 : _GEN_5547; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5549 = 10'h172 == _GEN_4[14:5] ? valid_370 : _GEN_5548; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5550 = 10'h173 == _GEN_4[14:5] ? valid_371 : _GEN_5549; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5551 = 10'h174 == _GEN_4[14:5] ? valid_372 : _GEN_5550; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5552 = 10'h175 == _GEN_4[14:5] ? valid_373 : _GEN_5551; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5553 = 10'h176 == _GEN_4[14:5] ? valid_374 : _GEN_5552; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5554 = 10'h177 == _GEN_4[14:5] ? valid_375 : _GEN_5553; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5555 = 10'h178 == _GEN_4[14:5] ? valid_376 : _GEN_5554; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5556 = 10'h179 == _GEN_4[14:5] ? valid_377 : _GEN_5555; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5557 = 10'h17a == _GEN_4[14:5] ? valid_378 : _GEN_5556; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5558 = 10'h17b == _GEN_4[14:5] ? valid_379 : _GEN_5557; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5559 = 10'h17c == _GEN_4[14:5] ? valid_380 : _GEN_5558; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5560 = 10'h17d == _GEN_4[14:5] ? valid_381 : _GEN_5559; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5561 = 10'h17e == _GEN_4[14:5] ? valid_382 : _GEN_5560; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5562 = 10'h17f == _GEN_4[14:5] ? valid_383 : _GEN_5561; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5563 = 10'h180 == _GEN_4[14:5] ? valid_384 : _GEN_5562; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5564 = 10'h181 == _GEN_4[14:5] ? valid_385 : _GEN_5563; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5565 = 10'h182 == _GEN_4[14:5] ? valid_386 : _GEN_5564; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5566 = 10'h183 == _GEN_4[14:5] ? valid_387 : _GEN_5565; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5567 = 10'h184 == _GEN_4[14:5] ? valid_388 : _GEN_5566; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5568 = 10'h185 == _GEN_4[14:5] ? valid_389 : _GEN_5567; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5569 = 10'h186 == _GEN_4[14:5] ? valid_390 : _GEN_5568; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5570 = 10'h187 == _GEN_4[14:5] ? valid_391 : _GEN_5569; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5571 = 10'h188 == _GEN_4[14:5] ? valid_392 : _GEN_5570; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5572 = 10'h189 == _GEN_4[14:5] ? valid_393 : _GEN_5571; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5573 = 10'h18a == _GEN_4[14:5] ? valid_394 : _GEN_5572; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5574 = 10'h18b == _GEN_4[14:5] ? valid_395 : _GEN_5573; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5575 = 10'h18c == _GEN_4[14:5] ? valid_396 : _GEN_5574; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5576 = 10'h18d == _GEN_4[14:5] ? valid_397 : _GEN_5575; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5577 = 10'h18e == _GEN_4[14:5] ? valid_398 : _GEN_5576; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5578 = 10'h18f == _GEN_4[14:5] ? valid_399 : _GEN_5577; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5579 = 10'h190 == _GEN_4[14:5] ? valid_400 : _GEN_5578; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5580 = 10'h191 == _GEN_4[14:5] ? valid_401 : _GEN_5579; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5581 = 10'h192 == _GEN_4[14:5] ? valid_402 : _GEN_5580; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5582 = 10'h193 == _GEN_4[14:5] ? valid_403 : _GEN_5581; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5583 = 10'h194 == _GEN_4[14:5] ? valid_404 : _GEN_5582; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5584 = 10'h195 == _GEN_4[14:5] ? valid_405 : _GEN_5583; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5585 = 10'h196 == _GEN_4[14:5] ? valid_406 : _GEN_5584; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5586 = 10'h197 == _GEN_4[14:5] ? valid_407 : _GEN_5585; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5587 = 10'h198 == _GEN_4[14:5] ? valid_408 : _GEN_5586; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5588 = 10'h199 == _GEN_4[14:5] ? valid_409 : _GEN_5587; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5589 = 10'h19a == _GEN_4[14:5] ? valid_410 : _GEN_5588; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5590 = 10'h19b == _GEN_4[14:5] ? valid_411 : _GEN_5589; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5591 = 10'h19c == _GEN_4[14:5] ? valid_412 : _GEN_5590; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5592 = 10'h19d == _GEN_4[14:5] ? valid_413 : _GEN_5591; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5593 = 10'h19e == _GEN_4[14:5] ? valid_414 : _GEN_5592; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5594 = 10'h19f == _GEN_4[14:5] ? valid_415 : _GEN_5593; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5595 = 10'h1a0 == _GEN_4[14:5] ? valid_416 : _GEN_5594; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5596 = 10'h1a1 == _GEN_4[14:5] ? valid_417 : _GEN_5595; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5597 = 10'h1a2 == _GEN_4[14:5] ? valid_418 : _GEN_5596; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5598 = 10'h1a3 == _GEN_4[14:5] ? valid_419 : _GEN_5597; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5599 = 10'h1a4 == _GEN_4[14:5] ? valid_420 : _GEN_5598; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5600 = 10'h1a5 == _GEN_4[14:5] ? valid_421 : _GEN_5599; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5601 = 10'h1a6 == _GEN_4[14:5] ? valid_422 : _GEN_5600; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5602 = 10'h1a7 == _GEN_4[14:5] ? valid_423 : _GEN_5601; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5603 = 10'h1a8 == _GEN_4[14:5] ? valid_424 : _GEN_5602; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5604 = 10'h1a9 == _GEN_4[14:5] ? valid_425 : _GEN_5603; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5605 = 10'h1aa == _GEN_4[14:5] ? valid_426 : _GEN_5604; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5606 = 10'h1ab == _GEN_4[14:5] ? valid_427 : _GEN_5605; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5607 = 10'h1ac == _GEN_4[14:5] ? valid_428 : _GEN_5606; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5608 = 10'h1ad == _GEN_4[14:5] ? valid_429 : _GEN_5607; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5609 = 10'h1ae == _GEN_4[14:5] ? valid_430 : _GEN_5608; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5610 = 10'h1af == _GEN_4[14:5] ? valid_431 : _GEN_5609; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5611 = 10'h1b0 == _GEN_4[14:5] ? valid_432 : _GEN_5610; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5612 = 10'h1b1 == _GEN_4[14:5] ? valid_433 : _GEN_5611; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5613 = 10'h1b2 == _GEN_4[14:5] ? valid_434 : _GEN_5612; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5614 = 10'h1b3 == _GEN_4[14:5] ? valid_435 : _GEN_5613; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5615 = 10'h1b4 == _GEN_4[14:5] ? valid_436 : _GEN_5614; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5616 = 10'h1b5 == _GEN_4[14:5] ? valid_437 : _GEN_5615; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5617 = 10'h1b6 == _GEN_4[14:5] ? valid_438 : _GEN_5616; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5618 = 10'h1b7 == _GEN_4[14:5] ? valid_439 : _GEN_5617; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5619 = 10'h1b8 == _GEN_4[14:5] ? valid_440 : _GEN_5618; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5620 = 10'h1b9 == _GEN_4[14:5] ? valid_441 : _GEN_5619; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5621 = 10'h1ba == _GEN_4[14:5] ? valid_442 : _GEN_5620; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5622 = 10'h1bb == _GEN_4[14:5] ? valid_443 : _GEN_5621; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5623 = 10'h1bc == _GEN_4[14:5] ? valid_444 : _GEN_5622; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5624 = 10'h1bd == _GEN_4[14:5] ? valid_445 : _GEN_5623; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5625 = 10'h1be == _GEN_4[14:5] ? valid_446 : _GEN_5624; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5626 = 10'h1bf == _GEN_4[14:5] ? valid_447 : _GEN_5625; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5627 = 10'h1c0 == _GEN_4[14:5] ? valid_448 : _GEN_5626; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5628 = 10'h1c1 == _GEN_4[14:5] ? valid_449 : _GEN_5627; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5629 = 10'h1c2 == _GEN_4[14:5] ? valid_450 : _GEN_5628; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5630 = 10'h1c3 == _GEN_4[14:5] ? valid_451 : _GEN_5629; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5631 = 10'h1c4 == _GEN_4[14:5] ? valid_452 : _GEN_5630; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5632 = 10'h1c5 == _GEN_4[14:5] ? valid_453 : _GEN_5631; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5633 = 10'h1c6 == _GEN_4[14:5] ? valid_454 : _GEN_5632; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5634 = 10'h1c7 == _GEN_4[14:5] ? valid_455 : _GEN_5633; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5635 = 10'h1c8 == _GEN_4[14:5] ? valid_456 : _GEN_5634; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5636 = 10'h1c9 == _GEN_4[14:5] ? valid_457 : _GEN_5635; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5637 = 10'h1ca == _GEN_4[14:5] ? valid_458 : _GEN_5636; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5638 = 10'h1cb == _GEN_4[14:5] ? valid_459 : _GEN_5637; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5639 = 10'h1cc == _GEN_4[14:5] ? valid_460 : _GEN_5638; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5640 = 10'h1cd == _GEN_4[14:5] ? valid_461 : _GEN_5639; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5641 = 10'h1ce == _GEN_4[14:5] ? valid_462 : _GEN_5640; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5642 = 10'h1cf == _GEN_4[14:5] ? valid_463 : _GEN_5641; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5643 = 10'h1d0 == _GEN_4[14:5] ? valid_464 : _GEN_5642; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5644 = 10'h1d1 == _GEN_4[14:5] ? valid_465 : _GEN_5643; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5645 = 10'h1d2 == _GEN_4[14:5] ? valid_466 : _GEN_5644; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5646 = 10'h1d3 == _GEN_4[14:5] ? valid_467 : _GEN_5645; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5647 = 10'h1d4 == _GEN_4[14:5] ? valid_468 : _GEN_5646; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5648 = 10'h1d5 == _GEN_4[14:5] ? valid_469 : _GEN_5647; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5649 = 10'h1d6 == _GEN_4[14:5] ? valid_470 : _GEN_5648; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5650 = 10'h1d7 == _GEN_4[14:5] ? valid_471 : _GEN_5649; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5651 = 10'h1d8 == _GEN_4[14:5] ? valid_472 : _GEN_5650; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5652 = 10'h1d9 == _GEN_4[14:5] ? valid_473 : _GEN_5651; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5653 = 10'h1da == _GEN_4[14:5] ? valid_474 : _GEN_5652; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5654 = 10'h1db == _GEN_4[14:5] ? valid_475 : _GEN_5653; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5655 = 10'h1dc == _GEN_4[14:5] ? valid_476 : _GEN_5654; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5656 = 10'h1dd == _GEN_4[14:5] ? valid_477 : _GEN_5655; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5657 = 10'h1de == _GEN_4[14:5] ? valid_478 : _GEN_5656; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5658 = 10'h1df == _GEN_4[14:5] ? valid_479 : _GEN_5657; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5659 = 10'h1e0 == _GEN_4[14:5] ? valid_480 : _GEN_5658; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5660 = 10'h1e1 == _GEN_4[14:5] ? valid_481 : _GEN_5659; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5661 = 10'h1e2 == _GEN_4[14:5] ? valid_482 : _GEN_5660; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5662 = 10'h1e3 == _GEN_4[14:5] ? valid_483 : _GEN_5661; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5663 = 10'h1e4 == _GEN_4[14:5] ? valid_484 : _GEN_5662; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5664 = 10'h1e5 == _GEN_4[14:5] ? valid_485 : _GEN_5663; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5665 = 10'h1e6 == _GEN_4[14:5] ? valid_486 : _GEN_5664; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5666 = 10'h1e7 == _GEN_4[14:5] ? valid_487 : _GEN_5665; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5667 = 10'h1e8 == _GEN_4[14:5] ? valid_488 : _GEN_5666; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5668 = 10'h1e9 == _GEN_4[14:5] ? valid_489 : _GEN_5667; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5669 = 10'h1ea == _GEN_4[14:5] ? valid_490 : _GEN_5668; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5670 = 10'h1eb == _GEN_4[14:5] ? valid_491 : _GEN_5669; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5671 = 10'h1ec == _GEN_4[14:5] ? valid_492 : _GEN_5670; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5672 = 10'h1ed == _GEN_4[14:5] ? valid_493 : _GEN_5671; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5673 = 10'h1ee == _GEN_4[14:5] ? valid_494 : _GEN_5672; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5674 = 10'h1ef == _GEN_4[14:5] ? valid_495 : _GEN_5673; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5675 = 10'h1f0 == _GEN_4[14:5] ? valid_496 : _GEN_5674; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5676 = 10'h1f1 == _GEN_4[14:5] ? valid_497 : _GEN_5675; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5677 = 10'h1f2 == _GEN_4[14:5] ? valid_498 : _GEN_5676; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5678 = 10'h1f3 == _GEN_4[14:5] ? valid_499 : _GEN_5677; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5679 = 10'h1f4 == _GEN_4[14:5] ? valid_500 : _GEN_5678; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5680 = 10'h1f5 == _GEN_4[14:5] ? valid_501 : _GEN_5679; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5681 = 10'h1f6 == _GEN_4[14:5] ? valid_502 : _GEN_5680; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5682 = 10'h1f7 == _GEN_4[14:5] ? valid_503 : _GEN_5681; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5683 = 10'h1f8 == _GEN_4[14:5] ? valid_504 : _GEN_5682; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5684 = 10'h1f9 == _GEN_4[14:5] ? valid_505 : _GEN_5683; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5685 = 10'h1fa == _GEN_4[14:5] ? valid_506 : _GEN_5684; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5686 = 10'h1fb == _GEN_4[14:5] ? valid_507 : _GEN_5685; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5687 = 10'h1fc == _GEN_4[14:5] ? valid_508 : _GEN_5686; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5688 = 10'h1fd == _GEN_4[14:5] ? valid_509 : _GEN_5687; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5689 = 10'h1fe == _GEN_4[14:5] ? valid_510 : _GEN_5688; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5690 = 10'h1ff == _GEN_4[14:5] ? valid_511 : _GEN_5689; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5691 = 10'h200 == _GEN_4[14:5] ? valid_512 : _GEN_5690; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5692 = 10'h201 == _GEN_4[14:5] ? valid_513 : _GEN_5691; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5693 = 10'h202 == _GEN_4[14:5] ? valid_514 : _GEN_5692; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5694 = 10'h203 == _GEN_4[14:5] ? valid_515 : _GEN_5693; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5695 = 10'h204 == _GEN_4[14:5] ? valid_516 : _GEN_5694; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5696 = 10'h205 == _GEN_4[14:5] ? valid_517 : _GEN_5695; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5697 = 10'h206 == _GEN_4[14:5] ? valid_518 : _GEN_5696; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5698 = 10'h207 == _GEN_4[14:5] ? valid_519 : _GEN_5697; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5699 = 10'h208 == _GEN_4[14:5] ? valid_520 : _GEN_5698; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5700 = 10'h209 == _GEN_4[14:5] ? valid_521 : _GEN_5699; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5701 = 10'h20a == _GEN_4[14:5] ? valid_522 : _GEN_5700; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5702 = 10'h20b == _GEN_4[14:5] ? valid_523 : _GEN_5701; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5703 = 10'h20c == _GEN_4[14:5] ? valid_524 : _GEN_5702; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5704 = 10'h20d == _GEN_4[14:5] ? valid_525 : _GEN_5703; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5705 = 10'h20e == _GEN_4[14:5] ? valid_526 : _GEN_5704; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5706 = 10'h20f == _GEN_4[14:5] ? valid_527 : _GEN_5705; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5707 = 10'h210 == _GEN_4[14:5] ? valid_528 : _GEN_5706; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5708 = 10'h211 == _GEN_4[14:5] ? valid_529 : _GEN_5707; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5709 = 10'h212 == _GEN_4[14:5] ? valid_530 : _GEN_5708; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5710 = 10'h213 == _GEN_4[14:5] ? valid_531 : _GEN_5709; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5711 = 10'h214 == _GEN_4[14:5] ? valid_532 : _GEN_5710; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5712 = 10'h215 == _GEN_4[14:5] ? valid_533 : _GEN_5711; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5713 = 10'h216 == _GEN_4[14:5] ? valid_534 : _GEN_5712; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5714 = 10'h217 == _GEN_4[14:5] ? valid_535 : _GEN_5713; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5715 = 10'h218 == _GEN_4[14:5] ? valid_536 : _GEN_5714; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5716 = 10'h219 == _GEN_4[14:5] ? valid_537 : _GEN_5715; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5717 = 10'h21a == _GEN_4[14:5] ? valid_538 : _GEN_5716; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5718 = 10'h21b == _GEN_4[14:5] ? valid_539 : _GEN_5717; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5719 = 10'h21c == _GEN_4[14:5] ? valid_540 : _GEN_5718; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5720 = 10'h21d == _GEN_4[14:5] ? valid_541 : _GEN_5719; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5721 = 10'h21e == _GEN_4[14:5] ? valid_542 : _GEN_5720; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5722 = 10'h21f == _GEN_4[14:5] ? valid_543 : _GEN_5721; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5723 = 10'h220 == _GEN_4[14:5] ? valid_544 : _GEN_5722; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5724 = 10'h221 == _GEN_4[14:5] ? valid_545 : _GEN_5723; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5725 = 10'h222 == _GEN_4[14:5] ? valid_546 : _GEN_5724; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5726 = 10'h223 == _GEN_4[14:5] ? valid_547 : _GEN_5725; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5727 = 10'h224 == _GEN_4[14:5] ? valid_548 : _GEN_5726; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5728 = 10'h225 == _GEN_4[14:5] ? valid_549 : _GEN_5727; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5729 = 10'h226 == _GEN_4[14:5] ? valid_550 : _GEN_5728; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5730 = 10'h227 == _GEN_4[14:5] ? valid_551 : _GEN_5729; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5731 = 10'h228 == _GEN_4[14:5] ? valid_552 : _GEN_5730; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5732 = 10'h229 == _GEN_4[14:5] ? valid_553 : _GEN_5731; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5733 = 10'h22a == _GEN_4[14:5] ? valid_554 : _GEN_5732; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5734 = 10'h22b == _GEN_4[14:5] ? valid_555 : _GEN_5733; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5735 = 10'h22c == _GEN_4[14:5] ? valid_556 : _GEN_5734; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5736 = 10'h22d == _GEN_4[14:5] ? valid_557 : _GEN_5735; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5737 = 10'h22e == _GEN_4[14:5] ? valid_558 : _GEN_5736; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5738 = 10'h22f == _GEN_4[14:5] ? valid_559 : _GEN_5737; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5739 = 10'h230 == _GEN_4[14:5] ? valid_560 : _GEN_5738; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5740 = 10'h231 == _GEN_4[14:5] ? valid_561 : _GEN_5739; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5741 = 10'h232 == _GEN_4[14:5] ? valid_562 : _GEN_5740; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5742 = 10'h233 == _GEN_4[14:5] ? valid_563 : _GEN_5741; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5743 = 10'h234 == _GEN_4[14:5] ? valid_564 : _GEN_5742; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5744 = 10'h235 == _GEN_4[14:5] ? valid_565 : _GEN_5743; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5745 = 10'h236 == _GEN_4[14:5] ? valid_566 : _GEN_5744; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5746 = 10'h237 == _GEN_4[14:5] ? valid_567 : _GEN_5745; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5747 = 10'h238 == _GEN_4[14:5] ? valid_568 : _GEN_5746; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5748 = 10'h239 == _GEN_4[14:5] ? valid_569 : _GEN_5747; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5749 = 10'h23a == _GEN_4[14:5] ? valid_570 : _GEN_5748; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5750 = 10'h23b == _GEN_4[14:5] ? valid_571 : _GEN_5749; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5751 = 10'h23c == _GEN_4[14:5] ? valid_572 : _GEN_5750; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5752 = 10'h23d == _GEN_4[14:5] ? valid_573 : _GEN_5751; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5753 = 10'h23e == _GEN_4[14:5] ? valid_574 : _GEN_5752; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5754 = 10'h23f == _GEN_4[14:5] ? valid_575 : _GEN_5753; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5755 = 10'h240 == _GEN_4[14:5] ? valid_576 : _GEN_5754; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5756 = 10'h241 == _GEN_4[14:5] ? valid_577 : _GEN_5755; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5757 = 10'h242 == _GEN_4[14:5] ? valid_578 : _GEN_5756; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5758 = 10'h243 == _GEN_4[14:5] ? valid_579 : _GEN_5757; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5759 = 10'h244 == _GEN_4[14:5] ? valid_580 : _GEN_5758; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5760 = 10'h245 == _GEN_4[14:5] ? valid_581 : _GEN_5759; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5761 = 10'h246 == _GEN_4[14:5] ? valid_582 : _GEN_5760; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5762 = 10'h247 == _GEN_4[14:5] ? valid_583 : _GEN_5761; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5763 = 10'h248 == _GEN_4[14:5] ? valid_584 : _GEN_5762; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5764 = 10'h249 == _GEN_4[14:5] ? valid_585 : _GEN_5763; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5765 = 10'h24a == _GEN_4[14:5] ? valid_586 : _GEN_5764; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5766 = 10'h24b == _GEN_4[14:5] ? valid_587 : _GEN_5765; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5767 = 10'h24c == _GEN_4[14:5] ? valid_588 : _GEN_5766; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5768 = 10'h24d == _GEN_4[14:5] ? valid_589 : _GEN_5767; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5769 = 10'h24e == _GEN_4[14:5] ? valid_590 : _GEN_5768; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5770 = 10'h24f == _GEN_4[14:5] ? valid_591 : _GEN_5769; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5771 = 10'h250 == _GEN_4[14:5] ? valid_592 : _GEN_5770; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5772 = 10'h251 == _GEN_4[14:5] ? valid_593 : _GEN_5771; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5773 = 10'h252 == _GEN_4[14:5] ? valid_594 : _GEN_5772; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5774 = 10'h253 == _GEN_4[14:5] ? valid_595 : _GEN_5773; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5775 = 10'h254 == _GEN_4[14:5] ? valid_596 : _GEN_5774; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5776 = 10'h255 == _GEN_4[14:5] ? valid_597 : _GEN_5775; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5777 = 10'h256 == _GEN_4[14:5] ? valid_598 : _GEN_5776; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5778 = 10'h257 == _GEN_4[14:5] ? valid_599 : _GEN_5777; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5779 = 10'h258 == _GEN_4[14:5] ? valid_600 : _GEN_5778; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5780 = 10'h259 == _GEN_4[14:5] ? valid_601 : _GEN_5779; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5781 = 10'h25a == _GEN_4[14:5] ? valid_602 : _GEN_5780; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5782 = 10'h25b == _GEN_4[14:5] ? valid_603 : _GEN_5781; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5783 = 10'h25c == _GEN_4[14:5] ? valid_604 : _GEN_5782; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5784 = 10'h25d == _GEN_4[14:5] ? valid_605 : _GEN_5783; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5785 = 10'h25e == _GEN_4[14:5] ? valid_606 : _GEN_5784; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5786 = 10'h25f == _GEN_4[14:5] ? valid_607 : _GEN_5785; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5787 = 10'h260 == _GEN_4[14:5] ? valid_608 : _GEN_5786; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5788 = 10'h261 == _GEN_4[14:5] ? valid_609 : _GEN_5787; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5789 = 10'h262 == _GEN_4[14:5] ? valid_610 : _GEN_5788; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5790 = 10'h263 == _GEN_4[14:5] ? valid_611 : _GEN_5789; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5791 = 10'h264 == _GEN_4[14:5] ? valid_612 : _GEN_5790; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5792 = 10'h265 == _GEN_4[14:5] ? valid_613 : _GEN_5791; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5793 = 10'h266 == _GEN_4[14:5] ? valid_614 : _GEN_5792; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5794 = 10'h267 == _GEN_4[14:5] ? valid_615 : _GEN_5793; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5795 = 10'h268 == _GEN_4[14:5] ? valid_616 : _GEN_5794; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5796 = 10'h269 == _GEN_4[14:5] ? valid_617 : _GEN_5795; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5797 = 10'h26a == _GEN_4[14:5] ? valid_618 : _GEN_5796; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5798 = 10'h26b == _GEN_4[14:5] ? valid_619 : _GEN_5797; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5799 = 10'h26c == _GEN_4[14:5] ? valid_620 : _GEN_5798; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5800 = 10'h26d == _GEN_4[14:5] ? valid_621 : _GEN_5799; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5801 = 10'h26e == _GEN_4[14:5] ? valid_622 : _GEN_5800; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5802 = 10'h26f == _GEN_4[14:5] ? valid_623 : _GEN_5801; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5803 = 10'h270 == _GEN_4[14:5] ? valid_624 : _GEN_5802; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5804 = 10'h271 == _GEN_4[14:5] ? valid_625 : _GEN_5803; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5805 = 10'h272 == _GEN_4[14:5] ? valid_626 : _GEN_5804; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5806 = 10'h273 == _GEN_4[14:5] ? valid_627 : _GEN_5805; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5807 = 10'h274 == _GEN_4[14:5] ? valid_628 : _GEN_5806; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5808 = 10'h275 == _GEN_4[14:5] ? valid_629 : _GEN_5807; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5809 = 10'h276 == _GEN_4[14:5] ? valid_630 : _GEN_5808; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5810 = 10'h277 == _GEN_4[14:5] ? valid_631 : _GEN_5809; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5811 = 10'h278 == _GEN_4[14:5] ? valid_632 : _GEN_5810; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5812 = 10'h279 == _GEN_4[14:5] ? valid_633 : _GEN_5811; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5813 = 10'h27a == _GEN_4[14:5] ? valid_634 : _GEN_5812; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5814 = 10'h27b == _GEN_4[14:5] ? valid_635 : _GEN_5813; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5815 = 10'h27c == _GEN_4[14:5] ? valid_636 : _GEN_5814; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5816 = 10'h27d == _GEN_4[14:5] ? valid_637 : _GEN_5815; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5817 = 10'h27e == _GEN_4[14:5] ? valid_638 : _GEN_5816; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5818 = 10'h27f == _GEN_4[14:5] ? valid_639 : _GEN_5817; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5819 = 10'h280 == _GEN_4[14:5] ? valid_640 : _GEN_5818; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5820 = 10'h281 == _GEN_4[14:5] ? valid_641 : _GEN_5819; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5821 = 10'h282 == _GEN_4[14:5] ? valid_642 : _GEN_5820; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5822 = 10'h283 == _GEN_4[14:5] ? valid_643 : _GEN_5821; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5823 = 10'h284 == _GEN_4[14:5] ? valid_644 : _GEN_5822; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5824 = 10'h285 == _GEN_4[14:5] ? valid_645 : _GEN_5823; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5825 = 10'h286 == _GEN_4[14:5] ? valid_646 : _GEN_5824; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5826 = 10'h287 == _GEN_4[14:5] ? valid_647 : _GEN_5825; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5827 = 10'h288 == _GEN_4[14:5] ? valid_648 : _GEN_5826; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5828 = 10'h289 == _GEN_4[14:5] ? valid_649 : _GEN_5827; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5829 = 10'h28a == _GEN_4[14:5] ? valid_650 : _GEN_5828; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5830 = 10'h28b == _GEN_4[14:5] ? valid_651 : _GEN_5829; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5831 = 10'h28c == _GEN_4[14:5] ? valid_652 : _GEN_5830; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5832 = 10'h28d == _GEN_4[14:5] ? valid_653 : _GEN_5831; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5833 = 10'h28e == _GEN_4[14:5] ? valid_654 : _GEN_5832; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5834 = 10'h28f == _GEN_4[14:5] ? valid_655 : _GEN_5833; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5835 = 10'h290 == _GEN_4[14:5] ? valid_656 : _GEN_5834; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5836 = 10'h291 == _GEN_4[14:5] ? valid_657 : _GEN_5835; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5837 = 10'h292 == _GEN_4[14:5] ? valid_658 : _GEN_5836; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5838 = 10'h293 == _GEN_4[14:5] ? valid_659 : _GEN_5837; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5839 = 10'h294 == _GEN_4[14:5] ? valid_660 : _GEN_5838; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5840 = 10'h295 == _GEN_4[14:5] ? valid_661 : _GEN_5839; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5841 = 10'h296 == _GEN_4[14:5] ? valid_662 : _GEN_5840; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5842 = 10'h297 == _GEN_4[14:5] ? valid_663 : _GEN_5841; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5843 = 10'h298 == _GEN_4[14:5] ? valid_664 : _GEN_5842; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5844 = 10'h299 == _GEN_4[14:5] ? valid_665 : _GEN_5843; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5845 = 10'h29a == _GEN_4[14:5] ? valid_666 : _GEN_5844; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5846 = 10'h29b == _GEN_4[14:5] ? valid_667 : _GEN_5845; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5847 = 10'h29c == _GEN_4[14:5] ? valid_668 : _GEN_5846; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5848 = 10'h29d == _GEN_4[14:5] ? valid_669 : _GEN_5847; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5849 = 10'h29e == _GEN_4[14:5] ? valid_670 : _GEN_5848; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5850 = 10'h29f == _GEN_4[14:5] ? valid_671 : _GEN_5849; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5851 = 10'h2a0 == _GEN_4[14:5] ? valid_672 : _GEN_5850; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5852 = 10'h2a1 == _GEN_4[14:5] ? valid_673 : _GEN_5851; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5853 = 10'h2a2 == _GEN_4[14:5] ? valid_674 : _GEN_5852; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5854 = 10'h2a3 == _GEN_4[14:5] ? valid_675 : _GEN_5853; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5855 = 10'h2a4 == _GEN_4[14:5] ? valid_676 : _GEN_5854; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5856 = 10'h2a5 == _GEN_4[14:5] ? valid_677 : _GEN_5855; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5857 = 10'h2a6 == _GEN_4[14:5] ? valid_678 : _GEN_5856; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5858 = 10'h2a7 == _GEN_4[14:5] ? valid_679 : _GEN_5857; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5859 = 10'h2a8 == _GEN_4[14:5] ? valid_680 : _GEN_5858; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5860 = 10'h2a9 == _GEN_4[14:5] ? valid_681 : _GEN_5859; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5861 = 10'h2aa == _GEN_4[14:5] ? valid_682 : _GEN_5860; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5862 = 10'h2ab == _GEN_4[14:5] ? valid_683 : _GEN_5861; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5863 = 10'h2ac == _GEN_4[14:5] ? valid_684 : _GEN_5862; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5864 = 10'h2ad == _GEN_4[14:5] ? valid_685 : _GEN_5863; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5865 = 10'h2ae == _GEN_4[14:5] ? valid_686 : _GEN_5864; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5866 = 10'h2af == _GEN_4[14:5] ? valid_687 : _GEN_5865; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5867 = 10'h2b0 == _GEN_4[14:5] ? valid_688 : _GEN_5866; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5868 = 10'h2b1 == _GEN_4[14:5] ? valid_689 : _GEN_5867; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5869 = 10'h2b2 == _GEN_4[14:5] ? valid_690 : _GEN_5868; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5870 = 10'h2b3 == _GEN_4[14:5] ? valid_691 : _GEN_5869; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5871 = 10'h2b4 == _GEN_4[14:5] ? valid_692 : _GEN_5870; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5872 = 10'h2b5 == _GEN_4[14:5] ? valid_693 : _GEN_5871; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5873 = 10'h2b6 == _GEN_4[14:5] ? valid_694 : _GEN_5872; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5874 = 10'h2b7 == _GEN_4[14:5] ? valid_695 : _GEN_5873; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5875 = 10'h2b8 == _GEN_4[14:5] ? valid_696 : _GEN_5874; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5876 = 10'h2b9 == _GEN_4[14:5] ? valid_697 : _GEN_5875; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5877 = 10'h2ba == _GEN_4[14:5] ? valid_698 : _GEN_5876; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5878 = 10'h2bb == _GEN_4[14:5] ? valid_699 : _GEN_5877; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5879 = 10'h2bc == _GEN_4[14:5] ? valid_700 : _GEN_5878; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5880 = 10'h2bd == _GEN_4[14:5] ? valid_701 : _GEN_5879; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5881 = 10'h2be == _GEN_4[14:5] ? valid_702 : _GEN_5880; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5882 = 10'h2bf == _GEN_4[14:5] ? valid_703 : _GEN_5881; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5883 = 10'h2c0 == _GEN_4[14:5] ? valid_704 : _GEN_5882; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5884 = 10'h2c1 == _GEN_4[14:5] ? valid_705 : _GEN_5883; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5885 = 10'h2c2 == _GEN_4[14:5] ? valid_706 : _GEN_5884; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5886 = 10'h2c3 == _GEN_4[14:5] ? valid_707 : _GEN_5885; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5887 = 10'h2c4 == _GEN_4[14:5] ? valid_708 : _GEN_5886; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5888 = 10'h2c5 == _GEN_4[14:5] ? valid_709 : _GEN_5887; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5889 = 10'h2c6 == _GEN_4[14:5] ? valid_710 : _GEN_5888; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5890 = 10'h2c7 == _GEN_4[14:5] ? valid_711 : _GEN_5889; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5891 = 10'h2c8 == _GEN_4[14:5] ? valid_712 : _GEN_5890; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5892 = 10'h2c9 == _GEN_4[14:5] ? valid_713 : _GEN_5891; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5893 = 10'h2ca == _GEN_4[14:5] ? valid_714 : _GEN_5892; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5894 = 10'h2cb == _GEN_4[14:5] ? valid_715 : _GEN_5893; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5895 = 10'h2cc == _GEN_4[14:5] ? valid_716 : _GEN_5894; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5896 = 10'h2cd == _GEN_4[14:5] ? valid_717 : _GEN_5895; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5897 = 10'h2ce == _GEN_4[14:5] ? valid_718 : _GEN_5896; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5898 = 10'h2cf == _GEN_4[14:5] ? valid_719 : _GEN_5897; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5899 = 10'h2d0 == _GEN_4[14:5] ? valid_720 : _GEN_5898; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5900 = 10'h2d1 == _GEN_4[14:5] ? valid_721 : _GEN_5899; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5901 = 10'h2d2 == _GEN_4[14:5] ? valid_722 : _GEN_5900; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5902 = 10'h2d3 == _GEN_4[14:5] ? valid_723 : _GEN_5901; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5903 = 10'h2d4 == _GEN_4[14:5] ? valid_724 : _GEN_5902; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5904 = 10'h2d5 == _GEN_4[14:5] ? valid_725 : _GEN_5903; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5905 = 10'h2d6 == _GEN_4[14:5] ? valid_726 : _GEN_5904; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5906 = 10'h2d7 == _GEN_4[14:5] ? valid_727 : _GEN_5905; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5907 = 10'h2d8 == _GEN_4[14:5] ? valid_728 : _GEN_5906; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5908 = 10'h2d9 == _GEN_4[14:5] ? valid_729 : _GEN_5907; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5909 = 10'h2da == _GEN_4[14:5] ? valid_730 : _GEN_5908; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5910 = 10'h2db == _GEN_4[14:5] ? valid_731 : _GEN_5909; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5911 = 10'h2dc == _GEN_4[14:5] ? valid_732 : _GEN_5910; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5912 = 10'h2dd == _GEN_4[14:5] ? valid_733 : _GEN_5911; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5913 = 10'h2de == _GEN_4[14:5] ? valid_734 : _GEN_5912; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5914 = 10'h2df == _GEN_4[14:5] ? valid_735 : _GEN_5913; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5915 = 10'h2e0 == _GEN_4[14:5] ? valid_736 : _GEN_5914; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5916 = 10'h2e1 == _GEN_4[14:5] ? valid_737 : _GEN_5915; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5917 = 10'h2e2 == _GEN_4[14:5] ? valid_738 : _GEN_5916; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5918 = 10'h2e3 == _GEN_4[14:5] ? valid_739 : _GEN_5917; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5919 = 10'h2e4 == _GEN_4[14:5] ? valid_740 : _GEN_5918; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5920 = 10'h2e5 == _GEN_4[14:5] ? valid_741 : _GEN_5919; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5921 = 10'h2e6 == _GEN_4[14:5] ? valid_742 : _GEN_5920; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5922 = 10'h2e7 == _GEN_4[14:5] ? valid_743 : _GEN_5921; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5923 = 10'h2e8 == _GEN_4[14:5] ? valid_744 : _GEN_5922; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5924 = 10'h2e9 == _GEN_4[14:5] ? valid_745 : _GEN_5923; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5925 = 10'h2ea == _GEN_4[14:5] ? valid_746 : _GEN_5924; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5926 = 10'h2eb == _GEN_4[14:5] ? valid_747 : _GEN_5925; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5927 = 10'h2ec == _GEN_4[14:5] ? valid_748 : _GEN_5926; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5928 = 10'h2ed == _GEN_4[14:5] ? valid_749 : _GEN_5927; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5929 = 10'h2ee == _GEN_4[14:5] ? valid_750 : _GEN_5928; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5930 = 10'h2ef == _GEN_4[14:5] ? valid_751 : _GEN_5929; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5931 = 10'h2f0 == _GEN_4[14:5] ? valid_752 : _GEN_5930; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5932 = 10'h2f1 == _GEN_4[14:5] ? valid_753 : _GEN_5931; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5933 = 10'h2f2 == _GEN_4[14:5] ? valid_754 : _GEN_5932; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5934 = 10'h2f3 == _GEN_4[14:5] ? valid_755 : _GEN_5933; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5935 = 10'h2f4 == _GEN_4[14:5] ? valid_756 : _GEN_5934; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5936 = 10'h2f5 == _GEN_4[14:5] ? valid_757 : _GEN_5935; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5937 = 10'h2f6 == _GEN_4[14:5] ? valid_758 : _GEN_5936; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5938 = 10'h2f7 == _GEN_4[14:5] ? valid_759 : _GEN_5937; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5939 = 10'h2f8 == _GEN_4[14:5] ? valid_760 : _GEN_5938; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5940 = 10'h2f9 == _GEN_4[14:5] ? valid_761 : _GEN_5939; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5941 = 10'h2fa == _GEN_4[14:5] ? valid_762 : _GEN_5940; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5942 = 10'h2fb == _GEN_4[14:5] ? valid_763 : _GEN_5941; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5943 = 10'h2fc == _GEN_4[14:5] ? valid_764 : _GEN_5942; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5944 = 10'h2fd == _GEN_4[14:5] ? valid_765 : _GEN_5943; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5945 = 10'h2fe == _GEN_4[14:5] ? valid_766 : _GEN_5944; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5946 = 10'h2ff == _GEN_4[14:5] ? valid_767 : _GEN_5945; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5947 = 10'h300 == _GEN_4[14:5] ? valid_768 : _GEN_5946; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5948 = 10'h301 == _GEN_4[14:5] ? valid_769 : _GEN_5947; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5949 = 10'h302 == _GEN_4[14:5] ? valid_770 : _GEN_5948; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5950 = 10'h303 == _GEN_4[14:5] ? valid_771 : _GEN_5949; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5951 = 10'h304 == _GEN_4[14:5] ? valid_772 : _GEN_5950; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5952 = 10'h305 == _GEN_4[14:5] ? valid_773 : _GEN_5951; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5953 = 10'h306 == _GEN_4[14:5] ? valid_774 : _GEN_5952; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5954 = 10'h307 == _GEN_4[14:5] ? valid_775 : _GEN_5953; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5955 = 10'h308 == _GEN_4[14:5] ? valid_776 : _GEN_5954; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5956 = 10'h309 == _GEN_4[14:5] ? valid_777 : _GEN_5955; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5957 = 10'h30a == _GEN_4[14:5] ? valid_778 : _GEN_5956; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5958 = 10'h30b == _GEN_4[14:5] ? valid_779 : _GEN_5957; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5959 = 10'h30c == _GEN_4[14:5] ? valid_780 : _GEN_5958; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5960 = 10'h30d == _GEN_4[14:5] ? valid_781 : _GEN_5959; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5961 = 10'h30e == _GEN_4[14:5] ? valid_782 : _GEN_5960; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5962 = 10'h30f == _GEN_4[14:5] ? valid_783 : _GEN_5961; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5963 = 10'h310 == _GEN_4[14:5] ? valid_784 : _GEN_5962; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5964 = 10'h311 == _GEN_4[14:5] ? valid_785 : _GEN_5963; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5965 = 10'h312 == _GEN_4[14:5] ? valid_786 : _GEN_5964; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5966 = 10'h313 == _GEN_4[14:5] ? valid_787 : _GEN_5965; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5967 = 10'h314 == _GEN_4[14:5] ? valid_788 : _GEN_5966; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5968 = 10'h315 == _GEN_4[14:5] ? valid_789 : _GEN_5967; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5969 = 10'h316 == _GEN_4[14:5] ? valid_790 : _GEN_5968; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5970 = 10'h317 == _GEN_4[14:5] ? valid_791 : _GEN_5969; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5971 = 10'h318 == _GEN_4[14:5] ? valid_792 : _GEN_5970; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5972 = 10'h319 == _GEN_4[14:5] ? valid_793 : _GEN_5971; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5973 = 10'h31a == _GEN_4[14:5] ? valid_794 : _GEN_5972; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5974 = 10'h31b == _GEN_4[14:5] ? valid_795 : _GEN_5973; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5975 = 10'h31c == _GEN_4[14:5] ? valid_796 : _GEN_5974; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5976 = 10'h31d == _GEN_4[14:5] ? valid_797 : _GEN_5975; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5977 = 10'h31e == _GEN_4[14:5] ? valid_798 : _GEN_5976; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5978 = 10'h31f == _GEN_4[14:5] ? valid_799 : _GEN_5977; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5979 = 10'h320 == _GEN_4[14:5] ? valid_800 : _GEN_5978; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5980 = 10'h321 == _GEN_4[14:5] ? valid_801 : _GEN_5979; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5981 = 10'h322 == _GEN_4[14:5] ? valid_802 : _GEN_5980; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5982 = 10'h323 == _GEN_4[14:5] ? valid_803 : _GEN_5981; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5983 = 10'h324 == _GEN_4[14:5] ? valid_804 : _GEN_5982; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5984 = 10'h325 == _GEN_4[14:5] ? valid_805 : _GEN_5983; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5985 = 10'h326 == _GEN_4[14:5] ? valid_806 : _GEN_5984; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5986 = 10'h327 == _GEN_4[14:5] ? valid_807 : _GEN_5985; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5987 = 10'h328 == _GEN_4[14:5] ? valid_808 : _GEN_5986; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5988 = 10'h329 == _GEN_4[14:5] ? valid_809 : _GEN_5987; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5989 = 10'h32a == _GEN_4[14:5] ? valid_810 : _GEN_5988; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5990 = 10'h32b == _GEN_4[14:5] ? valid_811 : _GEN_5989; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5991 = 10'h32c == _GEN_4[14:5] ? valid_812 : _GEN_5990; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5992 = 10'h32d == _GEN_4[14:5] ? valid_813 : _GEN_5991; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5993 = 10'h32e == _GEN_4[14:5] ? valid_814 : _GEN_5992; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5994 = 10'h32f == _GEN_4[14:5] ? valid_815 : _GEN_5993; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5995 = 10'h330 == _GEN_4[14:5] ? valid_816 : _GEN_5994; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5996 = 10'h331 == _GEN_4[14:5] ? valid_817 : _GEN_5995; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5997 = 10'h332 == _GEN_4[14:5] ? valid_818 : _GEN_5996; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5998 = 10'h333 == _GEN_4[14:5] ? valid_819 : _GEN_5997; // @[DCache.scala 234:{48,48}]
  wire  _GEN_5999 = 10'h334 == _GEN_4[14:5] ? valid_820 : _GEN_5998; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6000 = 10'h335 == _GEN_4[14:5] ? valid_821 : _GEN_5999; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6001 = 10'h336 == _GEN_4[14:5] ? valid_822 : _GEN_6000; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6002 = 10'h337 == _GEN_4[14:5] ? valid_823 : _GEN_6001; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6003 = 10'h338 == _GEN_4[14:5] ? valid_824 : _GEN_6002; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6004 = 10'h339 == _GEN_4[14:5] ? valid_825 : _GEN_6003; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6005 = 10'h33a == _GEN_4[14:5] ? valid_826 : _GEN_6004; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6006 = 10'h33b == _GEN_4[14:5] ? valid_827 : _GEN_6005; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6007 = 10'h33c == _GEN_4[14:5] ? valid_828 : _GEN_6006; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6008 = 10'h33d == _GEN_4[14:5] ? valid_829 : _GEN_6007; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6009 = 10'h33e == _GEN_4[14:5] ? valid_830 : _GEN_6008; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6010 = 10'h33f == _GEN_4[14:5] ? valid_831 : _GEN_6009; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6011 = 10'h340 == _GEN_4[14:5] ? valid_832 : _GEN_6010; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6012 = 10'h341 == _GEN_4[14:5] ? valid_833 : _GEN_6011; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6013 = 10'h342 == _GEN_4[14:5] ? valid_834 : _GEN_6012; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6014 = 10'h343 == _GEN_4[14:5] ? valid_835 : _GEN_6013; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6015 = 10'h344 == _GEN_4[14:5] ? valid_836 : _GEN_6014; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6016 = 10'h345 == _GEN_4[14:5] ? valid_837 : _GEN_6015; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6017 = 10'h346 == _GEN_4[14:5] ? valid_838 : _GEN_6016; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6018 = 10'h347 == _GEN_4[14:5] ? valid_839 : _GEN_6017; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6019 = 10'h348 == _GEN_4[14:5] ? valid_840 : _GEN_6018; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6020 = 10'h349 == _GEN_4[14:5] ? valid_841 : _GEN_6019; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6021 = 10'h34a == _GEN_4[14:5] ? valid_842 : _GEN_6020; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6022 = 10'h34b == _GEN_4[14:5] ? valid_843 : _GEN_6021; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6023 = 10'h34c == _GEN_4[14:5] ? valid_844 : _GEN_6022; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6024 = 10'h34d == _GEN_4[14:5] ? valid_845 : _GEN_6023; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6025 = 10'h34e == _GEN_4[14:5] ? valid_846 : _GEN_6024; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6026 = 10'h34f == _GEN_4[14:5] ? valid_847 : _GEN_6025; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6027 = 10'h350 == _GEN_4[14:5] ? valid_848 : _GEN_6026; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6028 = 10'h351 == _GEN_4[14:5] ? valid_849 : _GEN_6027; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6029 = 10'h352 == _GEN_4[14:5] ? valid_850 : _GEN_6028; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6030 = 10'h353 == _GEN_4[14:5] ? valid_851 : _GEN_6029; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6031 = 10'h354 == _GEN_4[14:5] ? valid_852 : _GEN_6030; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6032 = 10'h355 == _GEN_4[14:5] ? valid_853 : _GEN_6031; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6033 = 10'h356 == _GEN_4[14:5] ? valid_854 : _GEN_6032; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6034 = 10'h357 == _GEN_4[14:5] ? valid_855 : _GEN_6033; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6035 = 10'h358 == _GEN_4[14:5] ? valid_856 : _GEN_6034; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6036 = 10'h359 == _GEN_4[14:5] ? valid_857 : _GEN_6035; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6037 = 10'h35a == _GEN_4[14:5] ? valid_858 : _GEN_6036; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6038 = 10'h35b == _GEN_4[14:5] ? valid_859 : _GEN_6037; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6039 = 10'h35c == _GEN_4[14:5] ? valid_860 : _GEN_6038; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6040 = 10'h35d == _GEN_4[14:5] ? valid_861 : _GEN_6039; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6041 = 10'h35e == _GEN_4[14:5] ? valid_862 : _GEN_6040; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6042 = 10'h35f == _GEN_4[14:5] ? valid_863 : _GEN_6041; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6043 = 10'h360 == _GEN_4[14:5] ? valid_864 : _GEN_6042; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6044 = 10'h361 == _GEN_4[14:5] ? valid_865 : _GEN_6043; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6045 = 10'h362 == _GEN_4[14:5] ? valid_866 : _GEN_6044; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6046 = 10'h363 == _GEN_4[14:5] ? valid_867 : _GEN_6045; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6047 = 10'h364 == _GEN_4[14:5] ? valid_868 : _GEN_6046; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6048 = 10'h365 == _GEN_4[14:5] ? valid_869 : _GEN_6047; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6049 = 10'h366 == _GEN_4[14:5] ? valid_870 : _GEN_6048; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6050 = 10'h367 == _GEN_4[14:5] ? valid_871 : _GEN_6049; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6051 = 10'h368 == _GEN_4[14:5] ? valid_872 : _GEN_6050; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6052 = 10'h369 == _GEN_4[14:5] ? valid_873 : _GEN_6051; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6053 = 10'h36a == _GEN_4[14:5] ? valid_874 : _GEN_6052; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6054 = 10'h36b == _GEN_4[14:5] ? valid_875 : _GEN_6053; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6055 = 10'h36c == _GEN_4[14:5] ? valid_876 : _GEN_6054; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6056 = 10'h36d == _GEN_4[14:5] ? valid_877 : _GEN_6055; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6057 = 10'h36e == _GEN_4[14:5] ? valid_878 : _GEN_6056; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6058 = 10'h36f == _GEN_4[14:5] ? valid_879 : _GEN_6057; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6059 = 10'h370 == _GEN_4[14:5] ? valid_880 : _GEN_6058; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6060 = 10'h371 == _GEN_4[14:5] ? valid_881 : _GEN_6059; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6061 = 10'h372 == _GEN_4[14:5] ? valid_882 : _GEN_6060; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6062 = 10'h373 == _GEN_4[14:5] ? valid_883 : _GEN_6061; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6063 = 10'h374 == _GEN_4[14:5] ? valid_884 : _GEN_6062; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6064 = 10'h375 == _GEN_4[14:5] ? valid_885 : _GEN_6063; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6065 = 10'h376 == _GEN_4[14:5] ? valid_886 : _GEN_6064; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6066 = 10'h377 == _GEN_4[14:5] ? valid_887 : _GEN_6065; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6067 = 10'h378 == _GEN_4[14:5] ? valid_888 : _GEN_6066; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6068 = 10'h379 == _GEN_4[14:5] ? valid_889 : _GEN_6067; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6069 = 10'h37a == _GEN_4[14:5] ? valid_890 : _GEN_6068; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6070 = 10'h37b == _GEN_4[14:5] ? valid_891 : _GEN_6069; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6071 = 10'h37c == _GEN_4[14:5] ? valid_892 : _GEN_6070; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6072 = 10'h37d == _GEN_4[14:5] ? valid_893 : _GEN_6071; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6073 = 10'h37e == _GEN_4[14:5] ? valid_894 : _GEN_6072; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6074 = 10'h37f == _GEN_4[14:5] ? valid_895 : _GEN_6073; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6075 = 10'h380 == _GEN_4[14:5] ? valid_896 : _GEN_6074; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6076 = 10'h381 == _GEN_4[14:5] ? valid_897 : _GEN_6075; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6077 = 10'h382 == _GEN_4[14:5] ? valid_898 : _GEN_6076; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6078 = 10'h383 == _GEN_4[14:5] ? valid_899 : _GEN_6077; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6079 = 10'h384 == _GEN_4[14:5] ? valid_900 : _GEN_6078; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6080 = 10'h385 == _GEN_4[14:5] ? valid_901 : _GEN_6079; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6081 = 10'h386 == _GEN_4[14:5] ? valid_902 : _GEN_6080; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6082 = 10'h387 == _GEN_4[14:5] ? valid_903 : _GEN_6081; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6083 = 10'h388 == _GEN_4[14:5] ? valid_904 : _GEN_6082; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6084 = 10'h389 == _GEN_4[14:5] ? valid_905 : _GEN_6083; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6085 = 10'h38a == _GEN_4[14:5] ? valid_906 : _GEN_6084; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6086 = 10'h38b == _GEN_4[14:5] ? valid_907 : _GEN_6085; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6087 = 10'h38c == _GEN_4[14:5] ? valid_908 : _GEN_6086; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6088 = 10'h38d == _GEN_4[14:5] ? valid_909 : _GEN_6087; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6089 = 10'h38e == _GEN_4[14:5] ? valid_910 : _GEN_6088; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6090 = 10'h38f == _GEN_4[14:5] ? valid_911 : _GEN_6089; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6091 = 10'h390 == _GEN_4[14:5] ? valid_912 : _GEN_6090; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6092 = 10'h391 == _GEN_4[14:5] ? valid_913 : _GEN_6091; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6093 = 10'h392 == _GEN_4[14:5] ? valid_914 : _GEN_6092; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6094 = 10'h393 == _GEN_4[14:5] ? valid_915 : _GEN_6093; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6095 = 10'h394 == _GEN_4[14:5] ? valid_916 : _GEN_6094; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6096 = 10'h395 == _GEN_4[14:5] ? valid_917 : _GEN_6095; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6097 = 10'h396 == _GEN_4[14:5] ? valid_918 : _GEN_6096; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6098 = 10'h397 == _GEN_4[14:5] ? valid_919 : _GEN_6097; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6099 = 10'h398 == _GEN_4[14:5] ? valid_920 : _GEN_6098; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6100 = 10'h399 == _GEN_4[14:5] ? valid_921 : _GEN_6099; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6101 = 10'h39a == _GEN_4[14:5] ? valid_922 : _GEN_6100; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6102 = 10'h39b == _GEN_4[14:5] ? valid_923 : _GEN_6101; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6103 = 10'h39c == _GEN_4[14:5] ? valid_924 : _GEN_6102; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6104 = 10'h39d == _GEN_4[14:5] ? valid_925 : _GEN_6103; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6105 = 10'h39e == _GEN_4[14:5] ? valid_926 : _GEN_6104; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6106 = 10'h39f == _GEN_4[14:5] ? valid_927 : _GEN_6105; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6107 = 10'h3a0 == _GEN_4[14:5] ? valid_928 : _GEN_6106; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6108 = 10'h3a1 == _GEN_4[14:5] ? valid_929 : _GEN_6107; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6109 = 10'h3a2 == _GEN_4[14:5] ? valid_930 : _GEN_6108; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6110 = 10'h3a3 == _GEN_4[14:5] ? valid_931 : _GEN_6109; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6111 = 10'h3a4 == _GEN_4[14:5] ? valid_932 : _GEN_6110; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6112 = 10'h3a5 == _GEN_4[14:5] ? valid_933 : _GEN_6111; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6113 = 10'h3a6 == _GEN_4[14:5] ? valid_934 : _GEN_6112; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6114 = 10'h3a7 == _GEN_4[14:5] ? valid_935 : _GEN_6113; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6115 = 10'h3a8 == _GEN_4[14:5] ? valid_936 : _GEN_6114; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6116 = 10'h3a9 == _GEN_4[14:5] ? valid_937 : _GEN_6115; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6117 = 10'h3aa == _GEN_4[14:5] ? valid_938 : _GEN_6116; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6118 = 10'h3ab == _GEN_4[14:5] ? valid_939 : _GEN_6117; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6119 = 10'h3ac == _GEN_4[14:5] ? valid_940 : _GEN_6118; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6120 = 10'h3ad == _GEN_4[14:5] ? valid_941 : _GEN_6119; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6121 = 10'h3ae == _GEN_4[14:5] ? valid_942 : _GEN_6120; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6122 = 10'h3af == _GEN_4[14:5] ? valid_943 : _GEN_6121; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6123 = 10'h3b0 == _GEN_4[14:5] ? valid_944 : _GEN_6122; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6124 = 10'h3b1 == _GEN_4[14:5] ? valid_945 : _GEN_6123; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6125 = 10'h3b2 == _GEN_4[14:5] ? valid_946 : _GEN_6124; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6126 = 10'h3b3 == _GEN_4[14:5] ? valid_947 : _GEN_6125; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6127 = 10'h3b4 == _GEN_4[14:5] ? valid_948 : _GEN_6126; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6128 = 10'h3b5 == _GEN_4[14:5] ? valid_949 : _GEN_6127; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6129 = 10'h3b6 == _GEN_4[14:5] ? valid_950 : _GEN_6128; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6130 = 10'h3b7 == _GEN_4[14:5] ? valid_951 : _GEN_6129; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6131 = 10'h3b8 == _GEN_4[14:5] ? valid_952 : _GEN_6130; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6132 = 10'h3b9 == _GEN_4[14:5] ? valid_953 : _GEN_6131; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6133 = 10'h3ba == _GEN_4[14:5] ? valid_954 : _GEN_6132; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6134 = 10'h3bb == _GEN_4[14:5] ? valid_955 : _GEN_6133; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6135 = 10'h3bc == _GEN_4[14:5] ? valid_956 : _GEN_6134; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6136 = 10'h3bd == _GEN_4[14:5] ? valid_957 : _GEN_6135; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6137 = 10'h3be == _GEN_4[14:5] ? valid_958 : _GEN_6136; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6138 = 10'h3bf == _GEN_4[14:5] ? valid_959 : _GEN_6137; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6139 = 10'h3c0 == _GEN_4[14:5] ? valid_960 : _GEN_6138; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6140 = 10'h3c1 == _GEN_4[14:5] ? valid_961 : _GEN_6139; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6141 = 10'h3c2 == _GEN_4[14:5] ? valid_962 : _GEN_6140; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6142 = 10'h3c3 == _GEN_4[14:5] ? valid_963 : _GEN_6141; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6143 = 10'h3c4 == _GEN_4[14:5] ? valid_964 : _GEN_6142; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6144 = 10'h3c5 == _GEN_4[14:5] ? valid_965 : _GEN_6143; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6145 = 10'h3c6 == _GEN_4[14:5] ? valid_966 : _GEN_6144; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6146 = 10'h3c7 == _GEN_4[14:5] ? valid_967 : _GEN_6145; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6147 = 10'h3c8 == _GEN_4[14:5] ? valid_968 : _GEN_6146; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6148 = 10'h3c9 == _GEN_4[14:5] ? valid_969 : _GEN_6147; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6149 = 10'h3ca == _GEN_4[14:5] ? valid_970 : _GEN_6148; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6150 = 10'h3cb == _GEN_4[14:5] ? valid_971 : _GEN_6149; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6151 = 10'h3cc == _GEN_4[14:5] ? valid_972 : _GEN_6150; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6152 = 10'h3cd == _GEN_4[14:5] ? valid_973 : _GEN_6151; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6153 = 10'h3ce == _GEN_4[14:5] ? valid_974 : _GEN_6152; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6154 = 10'h3cf == _GEN_4[14:5] ? valid_975 : _GEN_6153; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6155 = 10'h3d0 == _GEN_4[14:5] ? valid_976 : _GEN_6154; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6156 = 10'h3d1 == _GEN_4[14:5] ? valid_977 : _GEN_6155; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6157 = 10'h3d2 == _GEN_4[14:5] ? valid_978 : _GEN_6156; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6158 = 10'h3d3 == _GEN_4[14:5] ? valid_979 : _GEN_6157; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6159 = 10'h3d4 == _GEN_4[14:5] ? valid_980 : _GEN_6158; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6160 = 10'h3d5 == _GEN_4[14:5] ? valid_981 : _GEN_6159; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6161 = 10'h3d6 == _GEN_4[14:5] ? valid_982 : _GEN_6160; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6162 = 10'h3d7 == _GEN_4[14:5] ? valid_983 : _GEN_6161; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6163 = 10'h3d8 == _GEN_4[14:5] ? valid_984 : _GEN_6162; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6164 = 10'h3d9 == _GEN_4[14:5] ? valid_985 : _GEN_6163; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6165 = 10'h3da == _GEN_4[14:5] ? valid_986 : _GEN_6164; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6166 = 10'h3db == _GEN_4[14:5] ? valid_987 : _GEN_6165; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6167 = 10'h3dc == _GEN_4[14:5] ? valid_988 : _GEN_6166; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6168 = 10'h3dd == _GEN_4[14:5] ? valid_989 : _GEN_6167; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6169 = 10'h3de == _GEN_4[14:5] ? valid_990 : _GEN_6168; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6170 = 10'h3df == _GEN_4[14:5] ? valid_991 : _GEN_6169; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6171 = 10'h3e0 == _GEN_4[14:5] ? valid_992 : _GEN_6170; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6172 = 10'h3e1 == _GEN_4[14:5] ? valid_993 : _GEN_6171; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6173 = 10'h3e2 == _GEN_4[14:5] ? valid_994 : _GEN_6172; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6174 = 10'h3e3 == _GEN_4[14:5] ? valid_995 : _GEN_6173; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6175 = 10'h3e4 == _GEN_4[14:5] ? valid_996 : _GEN_6174; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6176 = 10'h3e5 == _GEN_4[14:5] ? valid_997 : _GEN_6175; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6177 = 10'h3e6 == _GEN_4[14:5] ? valid_998 : _GEN_6176; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6178 = 10'h3e7 == _GEN_4[14:5] ? valid_999 : _GEN_6177; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6179 = 10'h3e8 == _GEN_4[14:5] ? valid_1000 : _GEN_6178; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6180 = 10'h3e9 == _GEN_4[14:5] ? valid_1001 : _GEN_6179; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6181 = 10'h3ea == _GEN_4[14:5] ? valid_1002 : _GEN_6180; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6182 = 10'h3eb == _GEN_4[14:5] ? valid_1003 : _GEN_6181; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6183 = 10'h3ec == _GEN_4[14:5] ? valid_1004 : _GEN_6182; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6184 = 10'h3ed == _GEN_4[14:5] ? valid_1005 : _GEN_6183; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6185 = 10'h3ee == _GEN_4[14:5] ? valid_1006 : _GEN_6184; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6186 = 10'h3ef == _GEN_4[14:5] ? valid_1007 : _GEN_6185; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6187 = 10'h3f0 == _GEN_4[14:5] ? valid_1008 : _GEN_6186; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6188 = 10'h3f1 == _GEN_4[14:5] ? valid_1009 : _GEN_6187; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6189 = 10'h3f2 == _GEN_4[14:5] ? valid_1010 : _GEN_6188; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6190 = 10'h3f3 == _GEN_4[14:5] ? valid_1011 : _GEN_6189; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6191 = 10'h3f4 == _GEN_4[14:5] ? valid_1012 : _GEN_6190; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6192 = 10'h3f5 == _GEN_4[14:5] ? valid_1013 : _GEN_6191; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6193 = 10'h3f6 == _GEN_4[14:5] ? valid_1014 : _GEN_6192; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6194 = 10'h3f7 == _GEN_4[14:5] ? valid_1015 : _GEN_6193; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6195 = 10'h3f8 == _GEN_4[14:5] ? valid_1016 : _GEN_6194; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6196 = 10'h3f9 == _GEN_4[14:5] ? valid_1017 : _GEN_6195; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6197 = 10'h3fa == _GEN_4[14:5] ? valid_1018 : _GEN_6196; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6198 = 10'h3fb == _GEN_4[14:5] ? valid_1019 : _GEN_6197; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6199 = 10'h3fc == _GEN_4[14:5] ? valid_1020 : _GEN_6198; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6200 = 10'h3fd == _GEN_4[14:5] ? valid_1021 : _GEN_6199; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6201 = 10'h3fe == _GEN_4[14:5] ? valid_1022 : _GEN_6200; // @[DCache.scala 234:{48,48}]
  wire  _GEN_6202 = 10'h3ff == _GEN_4[14:5] ? valid_1023 : _GEN_6201; // @[DCache.scala 234:{48,48}]
  wire  probe_hit = _GEN_6202 & _GEN_4[31:15] == probe_out_tag; // @[DCache.scala 234:48]
  reg [9:0] release_addr_aligned_REG; // @[DCache.scala 245:56]
  wire [31:0] release_addr_aligned = {array_out_tag,release_addr_aligned_REG,5'h0}; // @[Cat.scala 33:92]
  wire  _source_T_2 = _T_27 | _probing_T_1; // @[DCache.scala 249:47]
  reg [1:0] source; // @[Counter.scala 61:40]
  wire [1:0] _source_wrap_value_T_1 = source + 2'h1; // @[Counter.scala 77:24]
  wire [2:0] _x1_c_bits_T_opcode = probe_hit ? 3'h5 : 3'h4; // @[DCache.scala 259:33]
  wire [2:0] _x1_c_bits_T_param = probe_hit ? 3'h1 : 3'h5; // @[DCache.scala 259:33]
  wire [255:0] _x1_c_bits_T_data = probe_hit ? probe_out_data : 256'h0; // @[DCache.scala 259:33]
  wire  _io_cache_req_ready_T_3 = ~(probing | _tl_b_bits_r_T); // @[DCache.scala 266:44]
  SRAM array ( // @[DCache.scala 55:21]
    .clock(array_clock),
    .io_en(array_io_en),
    .io_addr(array_io_addr),
    .io_wdata(array_io_wdata),
    .io_wen(array_io_wen),
    .io_rdata(array_io_rdata)
  );
  assign auto_out_a_valid = state == 3'h4; // @[DCache.scala 257:24]
  assign auto_out_a_bits_source = source; // @[Edges.scala 345:17 349:15]
  assign auto_out_a_bits_address = {req_r_addr[31:5],5'h0}; // @[Cat.scala 33:92]
  assign auto_out_b_ready = ~probing & (~lrsc_reserved | lrsc_backoff); // @[DCache.scala 258:26]
  assign auto_out_c_valid = probing | state == 3'h2 & _GEN_1047; // @[DCache.scala 260:25]
  assign auto_out_c_bits_opcode = probing ? _x1_c_bits_T_opcode : 3'h7; // @[DCache.scala 259:20]
  assign auto_out_c_bits_param = probing ? _x1_c_bits_T_param : 3'h1; // @[DCache.scala 259:20]
  assign auto_out_c_bits_size = probing ? tl_b_bits_r_size : 3'h5; // @[DCache.scala 259:20]
  assign auto_out_c_bits_source = probing ? tl_b_bits_r_source : source; // @[DCache.scala 259:20]
  assign auto_out_c_bits_address = probing ? tl_b_bits_r_address : release_addr_aligned; // @[DCache.scala 259:20]
  assign auto_out_c_bits_data = probing ? _x1_c_bits_T_data : array_out_data; // @[DCache.scala 259:20]
  assign auto_out_d_ready = state == 3'h3 | state == 3'h5; // @[DCache.scala 261:43]
  assign auto_out_e_valid = state == 3'h6; // @[DCache.scala 263:24]
  assign auto_out_e_bits_sink = tl_d_bits_r_sink; // @[Edges.scala 438:17 439:12]
  assign io_cache_req_ready = state == 3'h0 & ~(probing | _tl_b_bits_r_T); // @[DCache.scala 266:41]
  assign io_cache_resp_valid = (state == 3'h1 & array_hit | _T_11) & _io_cache_req_ready_T_3; // @[DCache.scala 267:77]
  assign io_cache_resp_bits_rdata = is_sc_r ? sc_rdata_64 : rdata_64; // @[DCache.scala 269:25]
  assign array_clock = clock;
  assign array_io_en = _req_r_T | _array_io_en_T_1 | _tl_b_bits_r_T; // @[DCache.scala 70:45]
  assign array_io_addr = _tl_b_bits_r_T ? _GEN_4[14:5] : array_addr[14:5]; // @[DCache.scala 235:19 236:19 71:20]
  assign array_io_wdata = {array_wdata_tag,array_wdata_data}; // @[DCache.scala 72:35]
  assign array_io_wen = _array_io_en_T_1 & _GEN_3107; // @[DCache.scala 164:19 73:20]
  always @(posedge clock) begin
    if (reset) begin // @[Utils.scala 36:20]
      probing <= 1'h0; // @[Utils.scala 36:20]
    end else begin
      probing <= _GEN_5159;
    end
    if (reset) begin // @[DCache.scala 127:30]
      lrsc_reserved <= 1'h0; // @[DCache.scala 127:30]
    end else if (_array_io_en_T_1 & req_r_wen) begin // @[DCache.scala 147:32]
      lrsc_reserved <= 1'h0; // @[DCache.scala 148:19]
    end else if (_tl_b_bits_r_T & auto_out_b_bits_address[31:5] == lrsc_addr) begin // @[DCache.scala 139:73]
      lrsc_reserved <= 1'h0; // @[DCache.scala 140:19]
    end else begin
      lrsc_reserved <= _GEN_1048;
    end
    if (reset) begin // @[DCache.scala 129:30]
      lrsc_counter <= 5'h0; // @[DCache.scala 129:30]
    end else if (_array_io_en_T_1 & req_r_wen) begin // @[DCache.scala 147:32]
      lrsc_counter <= 5'h0; // @[DCache.scala 149:19]
    end else if (_tl_b_bits_r_T & auto_out_b_bits_address[31:5] == lrsc_addr) begin // @[DCache.scala 139:73]
      lrsc_counter <= 5'h0; // @[DCache.scala 141:19]
    end else if (lrsc_reserved & ~lrsc_backoff) begin // @[DCache.scala 136:40]
      lrsc_counter <= _lrsc_counter_T_1; // @[DCache.scala 137:18]
    end
    if (reset) begin // @[Reg.scala 35:20]
      tl_b_bits_r_size <= 3'h0; // @[Reg.scala 35:20]
    end else if (_tl_b_bits_r_T) begin // @[Reg.scala 36:18]
      tl_b_bits_r_size <= auto_out_b_bits_size; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      tl_b_bits_r_source <= 2'h0; // @[Reg.scala 35:20]
    end else if (_tl_b_bits_r_T) begin // @[Reg.scala 36:18]
      tl_b_bits_r_source <= auto_out_b_bits_source; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      tl_b_bits_r_address <= 32'h0; // @[Reg.scala 35:20]
    end else if (_tl_b_bits_r_T) begin // @[Reg.scala 36:18]
      tl_b_bits_r_address <= auto_out_b_bits_address; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[DCache.scala 60:118]
      state <= 3'h0; // @[DCache.scala 60:118]
    end else if (3'h0 == state) begin // @[DCache.scala 184:17]
      if (_req_r_T) begin // @[DCache.scala 186:22]
        if (sc_fail) begin // @[DCache.scala 187:21]
          state <= 3'h7;
        end else begin
          state <= 3'h1;
        end
      end
    end else if (3'h1 == state) begin // @[DCache.scala 184:17]
      if (_array_io_en_T_1) begin // @[DCache.scala 191:23]
        state <= 3'h0; // @[DCache.scala 192:15]
      end else begin
        state <= _GEN_5161;
      end
    end else if (3'h2 == state) begin // @[DCache.scala 184:17]
      state <= _GEN_5164;
    end else begin
      state <= _GEN_5174;
    end
    if (reset) begin // @[Reg.scala 35:20]
      tl_d_bits_r_sink <= 6'h0; // @[Reg.scala 35:20]
    end else if (_tl_d_bits_r_T) begin // @[Reg.scala 36:18]
      tl_d_bits_r_sink <= auto_out_d_bits_sink; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      tl_d_bits_r_data <= 256'h0; // @[Reg.scala 35:20]
    end else if (_tl_d_bits_r_T) begin // @[Reg.scala 36:18]
      tl_d_bits_r_data <= auto_out_d_bits_data; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      req_r_addr <= 39'h0; // @[Reg.scala 35:20]
    end else if (_req_r_T) begin // @[Reg.scala 36:18]
      req_r_addr <= io_cache_req_bits_addr; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      req_r_wdata <= 64'h0; // @[Reg.scala 35:20]
    end else if (_req_r_T) begin // @[Reg.scala 36:18]
      req_r_wdata <= io_cache_req_bits_wdata; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      req_r_wmask <= 8'h0; // @[Reg.scala 35:20]
    end else if (_req_r_T) begin // @[Reg.scala 36:18]
      req_r_wmask <= io_cache_req_bits_wmask; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      req_r_wen <= 1'h0; // @[Reg.scala 35:20]
    end else if (_req_r_T) begin // @[Reg.scala 36:18]
      req_r_wen <= io_cache_req_bits_wen; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      req_r_len <= 2'h0; // @[Reg.scala 35:20]
    end else if (_req_r_T) begin // @[Reg.scala 36:18]
      req_r_len <= io_cache_req_bits_len; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      req_r_lrsc <= 1'h0; // @[Reg.scala 35:20]
    end else if (_req_r_T) begin // @[Reg.scala 36:18]
      req_r_lrsc <= io_cache_req_bits_lrsc; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      req_r_amo <= 5'h0; // @[Reg.scala 35:20]
    end else if (_req_r_T) begin // @[Reg.scala 36:18]
      req_r_amo <= io_cache_req_bits_amo; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_0 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h0 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_0 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_0 <= _GEN_4134;
      end
    end else begin
      valid_0 <= _GEN_4134;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_1 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_1 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_1 <= _GEN_4135;
      end
    end else begin
      valid_1 <= _GEN_4135;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_2 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_2 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_2 <= _GEN_4136;
      end
    end else begin
      valid_2 <= _GEN_4136;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_3 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_3 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_3 <= _GEN_4137;
      end
    end else begin
      valid_3 <= _GEN_4137;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_4 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h4 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_4 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_4 <= _GEN_4138;
      end
    end else begin
      valid_4 <= _GEN_4138;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_5 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h5 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_5 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_5 <= _GEN_4139;
      end
    end else begin
      valid_5 <= _GEN_4139;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_6 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h6 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_6 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_6 <= _GEN_4140;
      end
    end else begin
      valid_6 <= _GEN_4140;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_7 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h7 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_7 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_7 <= _GEN_4141;
      end
    end else begin
      valid_7 <= _GEN_4141;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_8 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h8 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_8 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_8 <= _GEN_4142;
      end
    end else begin
      valid_8 <= _GEN_4142;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_9 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h9 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_9 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_9 <= _GEN_4143;
      end
    end else begin
      valid_9 <= _GEN_4143;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_10 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'ha == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_10 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_10 <= _GEN_4144;
      end
    end else begin
      valid_10 <= _GEN_4144;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_11 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hb == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_11 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_11 <= _GEN_4145;
      end
    end else begin
      valid_11 <= _GEN_4145;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_12 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hc == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_12 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_12 <= _GEN_4146;
      end
    end else begin
      valid_12 <= _GEN_4146;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_13 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hd == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_13 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_13 <= _GEN_4147;
      end
    end else begin
      valid_13 <= _GEN_4147;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_14 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'he == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_14 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_14 <= _GEN_4148;
      end
    end else begin
      valid_14 <= _GEN_4148;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_15 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hf == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_15 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_15 <= _GEN_4149;
      end
    end else begin
      valid_15 <= _GEN_4149;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_16 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h10 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_16 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_16 <= _GEN_4150;
      end
    end else begin
      valid_16 <= _GEN_4150;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_17 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h11 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_17 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_17 <= _GEN_4151;
      end
    end else begin
      valid_17 <= _GEN_4151;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_18 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h12 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_18 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_18 <= _GEN_4152;
      end
    end else begin
      valid_18 <= _GEN_4152;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_19 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h13 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_19 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_19 <= _GEN_4153;
      end
    end else begin
      valid_19 <= _GEN_4153;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_20 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h14 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_20 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_20 <= _GEN_4154;
      end
    end else begin
      valid_20 <= _GEN_4154;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_21 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h15 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_21 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_21 <= _GEN_4155;
      end
    end else begin
      valid_21 <= _GEN_4155;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_22 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h16 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_22 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_22 <= _GEN_4156;
      end
    end else begin
      valid_22 <= _GEN_4156;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_23 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h17 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_23 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_23 <= _GEN_4157;
      end
    end else begin
      valid_23 <= _GEN_4157;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_24 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h18 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_24 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_24 <= _GEN_4158;
      end
    end else begin
      valid_24 <= _GEN_4158;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_25 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h19 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_25 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_25 <= _GEN_4159;
      end
    end else begin
      valid_25 <= _GEN_4159;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_26 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1a == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_26 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_26 <= _GEN_4160;
      end
    end else begin
      valid_26 <= _GEN_4160;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_27 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1b == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_27 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_27 <= _GEN_4161;
      end
    end else begin
      valid_27 <= _GEN_4161;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_28 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1c == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_28 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_28 <= _GEN_4162;
      end
    end else begin
      valid_28 <= _GEN_4162;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_29 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1d == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_29 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_29 <= _GEN_4163;
      end
    end else begin
      valid_29 <= _GEN_4163;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_30 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1e == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_30 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_30 <= _GEN_4164;
      end
    end else begin
      valid_30 <= _GEN_4164;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_31 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1f == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_31 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_31 <= _GEN_4165;
      end
    end else begin
      valid_31 <= _GEN_4165;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_32 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h20 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_32 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_32 <= _GEN_4166;
      end
    end else begin
      valid_32 <= _GEN_4166;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_33 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h21 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_33 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_33 <= _GEN_4167;
      end
    end else begin
      valid_33 <= _GEN_4167;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_34 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h22 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_34 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_34 <= _GEN_4168;
      end
    end else begin
      valid_34 <= _GEN_4168;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_35 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h23 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_35 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_35 <= _GEN_4169;
      end
    end else begin
      valid_35 <= _GEN_4169;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_36 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h24 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_36 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_36 <= _GEN_4170;
      end
    end else begin
      valid_36 <= _GEN_4170;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_37 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h25 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_37 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_37 <= _GEN_4171;
      end
    end else begin
      valid_37 <= _GEN_4171;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_38 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h26 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_38 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_38 <= _GEN_4172;
      end
    end else begin
      valid_38 <= _GEN_4172;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_39 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h27 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_39 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_39 <= _GEN_4173;
      end
    end else begin
      valid_39 <= _GEN_4173;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_40 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h28 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_40 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_40 <= _GEN_4174;
      end
    end else begin
      valid_40 <= _GEN_4174;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_41 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h29 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_41 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_41 <= _GEN_4175;
      end
    end else begin
      valid_41 <= _GEN_4175;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_42 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2a == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_42 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_42 <= _GEN_4176;
      end
    end else begin
      valid_42 <= _GEN_4176;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_43 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2b == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_43 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_43 <= _GEN_4177;
      end
    end else begin
      valid_43 <= _GEN_4177;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_44 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2c == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_44 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_44 <= _GEN_4178;
      end
    end else begin
      valid_44 <= _GEN_4178;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_45 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2d == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_45 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_45 <= _GEN_4179;
      end
    end else begin
      valid_45 <= _GEN_4179;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_46 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2e == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_46 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_46 <= _GEN_4180;
      end
    end else begin
      valid_46 <= _GEN_4180;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_47 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2f == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_47 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_47 <= _GEN_4181;
      end
    end else begin
      valid_47 <= _GEN_4181;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_48 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h30 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_48 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_48 <= _GEN_4182;
      end
    end else begin
      valid_48 <= _GEN_4182;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_49 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h31 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_49 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_49 <= _GEN_4183;
      end
    end else begin
      valid_49 <= _GEN_4183;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_50 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h32 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_50 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_50 <= _GEN_4184;
      end
    end else begin
      valid_50 <= _GEN_4184;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_51 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h33 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_51 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_51 <= _GEN_4185;
      end
    end else begin
      valid_51 <= _GEN_4185;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_52 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h34 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_52 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_52 <= _GEN_4186;
      end
    end else begin
      valid_52 <= _GEN_4186;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_53 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h35 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_53 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_53 <= _GEN_4187;
      end
    end else begin
      valid_53 <= _GEN_4187;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_54 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h36 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_54 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_54 <= _GEN_4188;
      end
    end else begin
      valid_54 <= _GEN_4188;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_55 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h37 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_55 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_55 <= _GEN_4189;
      end
    end else begin
      valid_55 <= _GEN_4189;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_56 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h38 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_56 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_56 <= _GEN_4190;
      end
    end else begin
      valid_56 <= _GEN_4190;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_57 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h39 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_57 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_57 <= _GEN_4191;
      end
    end else begin
      valid_57 <= _GEN_4191;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_58 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3a == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_58 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_58 <= _GEN_4192;
      end
    end else begin
      valid_58 <= _GEN_4192;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_59 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3b == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_59 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_59 <= _GEN_4193;
      end
    end else begin
      valid_59 <= _GEN_4193;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_60 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3c == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_60 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_60 <= _GEN_4194;
      end
    end else begin
      valid_60 <= _GEN_4194;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_61 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3d == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_61 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_61 <= _GEN_4195;
      end
    end else begin
      valid_61 <= _GEN_4195;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_62 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3e == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_62 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_62 <= _GEN_4196;
      end
    end else begin
      valid_62 <= _GEN_4196;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_63 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3f == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_63 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_63 <= _GEN_4197;
      end
    end else begin
      valid_63 <= _GEN_4197;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_64 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h40 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_64 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_64 <= _GEN_4198;
      end
    end else begin
      valid_64 <= _GEN_4198;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_65 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h41 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_65 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_65 <= _GEN_4199;
      end
    end else begin
      valid_65 <= _GEN_4199;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_66 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h42 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_66 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_66 <= _GEN_4200;
      end
    end else begin
      valid_66 <= _GEN_4200;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_67 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h43 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_67 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_67 <= _GEN_4201;
      end
    end else begin
      valid_67 <= _GEN_4201;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_68 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h44 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_68 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_68 <= _GEN_4202;
      end
    end else begin
      valid_68 <= _GEN_4202;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_69 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h45 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_69 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_69 <= _GEN_4203;
      end
    end else begin
      valid_69 <= _GEN_4203;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_70 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h46 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_70 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_70 <= _GEN_4204;
      end
    end else begin
      valid_70 <= _GEN_4204;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_71 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h47 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_71 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_71 <= _GEN_4205;
      end
    end else begin
      valid_71 <= _GEN_4205;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_72 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h48 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_72 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_72 <= _GEN_4206;
      end
    end else begin
      valid_72 <= _GEN_4206;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_73 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h49 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_73 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_73 <= _GEN_4207;
      end
    end else begin
      valid_73 <= _GEN_4207;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_74 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h4a == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_74 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_74 <= _GEN_4208;
      end
    end else begin
      valid_74 <= _GEN_4208;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_75 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h4b == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_75 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_75 <= _GEN_4209;
      end
    end else begin
      valid_75 <= _GEN_4209;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_76 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h4c == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_76 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_76 <= _GEN_4210;
      end
    end else begin
      valid_76 <= _GEN_4210;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_77 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h4d == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_77 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_77 <= _GEN_4211;
      end
    end else begin
      valid_77 <= _GEN_4211;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_78 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h4e == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_78 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_78 <= _GEN_4212;
      end
    end else begin
      valid_78 <= _GEN_4212;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_79 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h4f == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_79 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_79 <= _GEN_4213;
      end
    end else begin
      valid_79 <= _GEN_4213;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_80 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h50 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_80 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_80 <= _GEN_4214;
      end
    end else begin
      valid_80 <= _GEN_4214;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_81 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h51 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_81 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_81 <= _GEN_4215;
      end
    end else begin
      valid_81 <= _GEN_4215;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_82 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h52 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_82 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_82 <= _GEN_4216;
      end
    end else begin
      valid_82 <= _GEN_4216;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_83 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h53 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_83 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_83 <= _GEN_4217;
      end
    end else begin
      valid_83 <= _GEN_4217;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_84 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h54 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_84 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_84 <= _GEN_4218;
      end
    end else begin
      valid_84 <= _GEN_4218;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_85 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h55 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_85 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_85 <= _GEN_4219;
      end
    end else begin
      valid_85 <= _GEN_4219;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_86 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h56 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_86 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_86 <= _GEN_4220;
      end
    end else begin
      valid_86 <= _GEN_4220;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_87 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h57 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_87 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_87 <= _GEN_4221;
      end
    end else begin
      valid_87 <= _GEN_4221;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_88 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h58 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_88 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_88 <= _GEN_4222;
      end
    end else begin
      valid_88 <= _GEN_4222;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_89 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h59 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_89 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_89 <= _GEN_4223;
      end
    end else begin
      valid_89 <= _GEN_4223;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_90 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h5a == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_90 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_90 <= _GEN_4224;
      end
    end else begin
      valid_90 <= _GEN_4224;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_91 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h5b == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_91 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_91 <= _GEN_4225;
      end
    end else begin
      valid_91 <= _GEN_4225;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_92 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h5c == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_92 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_92 <= _GEN_4226;
      end
    end else begin
      valid_92 <= _GEN_4226;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_93 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h5d == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_93 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_93 <= _GEN_4227;
      end
    end else begin
      valid_93 <= _GEN_4227;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_94 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h5e == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_94 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_94 <= _GEN_4228;
      end
    end else begin
      valid_94 <= _GEN_4228;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_95 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h5f == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_95 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_95 <= _GEN_4229;
      end
    end else begin
      valid_95 <= _GEN_4229;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_96 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h60 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_96 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_96 <= _GEN_4230;
      end
    end else begin
      valid_96 <= _GEN_4230;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_97 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h61 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_97 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_97 <= _GEN_4231;
      end
    end else begin
      valid_97 <= _GEN_4231;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_98 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h62 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_98 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_98 <= _GEN_4232;
      end
    end else begin
      valid_98 <= _GEN_4232;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_99 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h63 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_99 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_99 <= _GEN_4233;
      end
    end else begin
      valid_99 <= _GEN_4233;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_100 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h64 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_100 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_100 <= _GEN_4234;
      end
    end else begin
      valid_100 <= _GEN_4234;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_101 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h65 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_101 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_101 <= _GEN_4235;
      end
    end else begin
      valid_101 <= _GEN_4235;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_102 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h66 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_102 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_102 <= _GEN_4236;
      end
    end else begin
      valid_102 <= _GEN_4236;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_103 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h67 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_103 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_103 <= _GEN_4237;
      end
    end else begin
      valid_103 <= _GEN_4237;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_104 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h68 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_104 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_104 <= _GEN_4238;
      end
    end else begin
      valid_104 <= _GEN_4238;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_105 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h69 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_105 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_105 <= _GEN_4239;
      end
    end else begin
      valid_105 <= _GEN_4239;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_106 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h6a == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_106 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_106 <= _GEN_4240;
      end
    end else begin
      valid_106 <= _GEN_4240;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_107 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h6b == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_107 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_107 <= _GEN_4241;
      end
    end else begin
      valid_107 <= _GEN_4241;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_108 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h6c == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_108 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_108 <= _GEN_4242;
      end
    end else begin
      valid_108 <= _GEN_4242;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_109 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h6d == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_109 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_109 <= _GEN_4243;
      end
    end else begin
      valid_109 <= _GEN_4243;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_110 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h6e == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_110 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_110 <= _GEN_4244;
      end
    end else begin
      valid_110 <= _GEN_4244;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_111 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h6f == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_111 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_111 <= _GEN_4245;
      end
    end else begin
      valid_111 <= _GEN_4245;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_112 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h70 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_112 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_112 <= _GEN_4246;
      end
    end else begin
      valid_112 <= _GEN_4246;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_113 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h71 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_113 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_113 <= _GEN_4247;
      end
    end else begin
      valid_113 <= _GEN_4247;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_114 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h72 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_114 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_114 <= _GEN_4248;
      end
    end else begin
      valid_114 <= _GEN_4248;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_115 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h73 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_115 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_115 <= _GEN_4249;
      end
    end else begin
      valid_115 <= _GEN_4249;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_116 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h74 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_116 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_116 <= _GEN_4250;
      end
    end else begin
      valid_116 <= _GEN_4250;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_117 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h75 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_117 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_117 <= _GEN_4251;
      end
    end else begin
      valid_117 <= _GEN_4251;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_118 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h76 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_118 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_118 <= _GEN_4252;
      end
    end else begin
      valid_118 <= _GEN_4252;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_119 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h77 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_119 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_119 <= _GEN_4253;
      end
    end else begin
      valid_119 <= _GEN_4253;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_120 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h78 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_120 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_120 <= _GEN_4254;
      end
    end else begin
      valid_120 <= _GEN_4254;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_121 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h79 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_121 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_121 <= _GEN_4255;
      end
    end else begin
      valid_121 <= _GEN_4255;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_122 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h7a == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_122 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_122 <= _GEN_4256;
      end
    end else begin
      valid_122 <= _GEN_4256;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_123 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h7b == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_123 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_123 <= _GEN_4257;
      end
    end else begin
      valid_123 <= _GEN_4257;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_124 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h7c == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_124 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_124 <= _GEN_4258;
      end
    end else begin
      valid_124 <= _GEN_4258;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_125 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h7d == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_125 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_125 <= _GEN_4259;
      end
    end else begin
      valid_125 <= _GEN_4259;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_126 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h7e == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_126 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_126 <= _GEN_4260;
      end
    end else begin
      valid_126 <= _GEN_4260;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_127 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h7f == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_127 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_127 <= _GEN_4261;
      end
    end else begin
      valid_127 <= _GEN_4261;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_128 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h80 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_128 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_128 <= _GEN_4262;
      end
    end else begin
      valid_128 <= _GEN_4262;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_129 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h81 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_129 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_129 <= _GEN_4263;
      end
    end else begin
      valid_129 <= _GEN_4263;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_130 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h82 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_130 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_130 <= _GEN_4264;
      end
    end else begin
      valid_130 <= _GEN_4264;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_131 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h83 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_131 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_131 <= _GEN_4265;
      end
    end else begin
      valid_131 <= _GEN_4265;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_132 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h84 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_132 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_132 <= _GEN_4266;
      end
    end else begin
      valid_132 <= _GEN_4266;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_133 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h85 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_133 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_133 <= _GEN_4267;
      end
    end else begin
      valid_133 <= _GEN_4267;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_134 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h86 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_134 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_134 <= _GEN_4268;
      end
    end else begin
      valid_134 <= _GEN_4268;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_135 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h87 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_135 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_135 <= _GEN_4269;
      end
    end else begin
      valid_135 <= _GEN_4269;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_136 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h88 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_136 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_136 <= _GEN_4270;
      end
    end else begin
      valid_136 <= _GEN_4270;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_137 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h89 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_137 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_137 <= _GEN_4271;
      end
    end else begin
      valid_137 <= _GEN_4271;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_138 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h8a == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_138 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_138 <= _GEN_4272;
      end
    end else begin
      valid_138 <= _GEN_4272;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_139 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h8b == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_139 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_139 <= _GEN_4273;
      end
    end else begin
      valid_139 <= _GEN_4273;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_140 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h8c == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_140 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_140 <= _GEN_4274;
      end
    end else begin
      valid_140 <= _GEN_4274;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_141 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h8d == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_141 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_141 <= _GEN_4275;
      end
    end else begin
      valid_141 <= _GEN_4275;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_142 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h8e == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_142 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_142 <= _GEN_4276;
      end
    end else begin
      valid_142 <= _GEN_4276;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_143 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h8f == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_143 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_143 <= _GEN_4277;
      end
    end else begin
      valid_143 <= _GEN_4277;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_144 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h90 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_144 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_144 <= _GEN_4278;
      end
    end else begin
      valid_144 <= _GEN_4278;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_145 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h91 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_145 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_145 <= _GEN_4279;
      end
    end else begin
      valid_145 <= _GEN_4279;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_146 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h92 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_146 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_146 <= _GEN_4280;
      end
    end else begin
      valid_146 <= _GEN_4280;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_147 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h93 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_147 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_147 <= _GEN_4281;
      end
    end else begin
      valid_147 <= _GEN_4281;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_148 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h94 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_148 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_148 <= _GEN_4282;
      end
    end else begin
      valid_148 <= _GEN_4282;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_149 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h95 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_149 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_149 <= _GEN_4283;
      end
    end else begin
      valid_149 <= _GEN_4283;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_150 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h96 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_150 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_150 <= _GEN_4284;
      end
    end else begin
      valid_150 <= _GEN_4284;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_151 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h97 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_151 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_151 <= _GEN_4285;
      end
    end else begin
      valid_151 <= _GEN_4285;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_152 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h98 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_152 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_152 <= _GEN_4286;
      end
    end else begin
      valid_152 <= _GEN_4286;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_153 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h99 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_153 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_153 <= _GEN_4287;
      end
    end else begin
      valid_153 <= _GEN_4287;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_154 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h9a == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_154 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_154 <= _GEN_4288;
      end
    end else begin
      valid_154 <= _GEN_4288;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_155 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h9b == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_155 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_155 <= _GEN_4289;
      end
    end else begin
      valid_155 <= _GEN_4289;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_156 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h9c == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_156 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_156 <= _GEN_4290;
      end
    end else begin
      valid_156 <= _GEN_4290;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_157 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h9d == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_157 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_157 <= _GEN_4291;
      end
    end else begin
      valid_157 <= _GEN_4291;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_158 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h9e == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_158 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_158 <= _GEN_4292;
      end
    end else begin
      valid_158 <= _GEN_4292;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_159 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h9f == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_159 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_159 <= _GEN_4293;
      end
    end else begin
      valid_159 <= _GEN_4293;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_160 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'ha0 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_160 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_160 <= _GEN_4294;
      end
    end else begin
      valid_160 <= _GEN_4294;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_161 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'ha1 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_161 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_161 <= _GEN_4295;
      end
    end else begin
      valid_161 <= _GEN_4295;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_162 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'ha2 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_162 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_162 <= _GEN_4296;
      end
    end else begin
      valid_162 <= _GEN_4296;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_163 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'ha3 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_163 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_163 <= _GEN_4297;
      end
    end else begin
      valid_163 <= _GEN_4297;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_164 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'ha4 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_164 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_164 <= _GEN_4298;
      end
    end else begin
      valid_164 <= _GEN_4298;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_165 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'ha5 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_165 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_165 <= _GEN_4299;
      end
    end else begin
      valid_165 <= _GEN_4299;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_166 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'ha6 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_166 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_166 <= _GEN_4300;
      end
    end else begin
      valid_166 <= _GEN_4300;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_167 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'ha7 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_167 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_167 <= _GEN_4301;
      end
    end else begin
      valid_167 <= _GEN_4301;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_168 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'ha8 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_168 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_168 <= _GEN_4302;
      end
    end else begin
      valid_168 <= _GEN_4302;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_169 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'ha9 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_169 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_169 <= _GEN_4303;
      end
    end else begin
      valid_169 <= _GEN_4303;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_170 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'haa == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_170 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_170 <= _GEN_4304;
      end
    end else begin
      valid_170 <= _GEN_4304;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_171 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hab == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_171 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_171 <= _GEN_4305;
      end
    end else begin
      valid_171 <= _GEN_4305;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_172 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hac == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_172 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_172 <= _GEN_4306;
      end
    end else begin
      valid_172 <= _GEN_4306;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_173 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'had == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_173 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_173 <= _GEN_4307;
      end
    end else begin
      valid_173 <= _GEN_4307;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_174 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hae == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_174 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_174 <= _GEN_4308;
      end
    end else begin
      valid_174 <= _GEN_4308;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_175 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'haf == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_175 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_175 <= _GEN_4309;
      end
    end else begin
      valid_175 <= _GEN_4309;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_176 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hb0 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_176 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_176 <= _GEN_4310;
      end
    end else begin
      valid_176 <= _GEN_4310;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_177 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hb1 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_177 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_177 <= _GEN_4311;
      end
    end else begin
      valid_177 <= _GEN_4311;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_178 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hb2 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_178 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_178 <= _GEN_4312;
      end
    end else begin
      valid_178 <= _GEN_4312;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_179 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hb3 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_179 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_179 <= _GEN_4313;
      end
    end else begin
      valid_179 <= _GEN_4313;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_180 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hb4 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_180 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_180 <= _GEN_4314;
      end
    end else begin
      valid_180 <= _GEN_4314;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_181 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hb5 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_181 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_181 <= _GEN_4315;
      end
    end else begin
      valid_181 <= _GEN_4315;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_182 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hb6 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_182 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_182 <= _GEN_4316;
      end
    end else begin
      valid_182 <= _GEN_4316;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_183 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hb7 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_183 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_183 <= _GEN_4317;
      end
    end else begin
      valid_183 <= _GEN_4317;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_184 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hb8 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_184 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_184 <= _GEN_4318;
      end
    end else begin
      valid_184 <= _GEN_4318;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_185 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hb9 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_185 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_185 <= _GEN_4319;
      end
    end else begin
      valid_185 <= _GEN_4319;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_186 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hba == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_186 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_186 <= _GEN_4320;
      end
    end else begin
      valid_186 <= _GEN_4320;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_187 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hbb == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_187 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_187 <= _GEN_4321;
      end
    end else begin
      valid_187 <= _GEN_4321;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_188 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hbc == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_188 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_188 <= _GEN_4322;
      end
    end else begin
      valid_188 <= _GEN_4322;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_189 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hbd == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_189 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_189 <= _GEN_4323;
      end
    end else begin
      valid_189 <= _GEN_4323;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_190 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hbe == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_190 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_190 <= _GEN_4324;
      end
    end else begin
      valid_190 <= _GEN_4324;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_191 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hbf == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_191 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_191 <= _GEN_4325;
      end
    end else begin
      valid_191 <= _GEN_4325;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_192 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hc0 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_192 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_192 <= _GEN_4326;
      end
    end else begin
      valid_192 <= _GEN_4326;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_193 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hc1 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_193 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_193 <= _GEN_4327;
      end
    end else begin
      valid_193 <= _GEN_4327;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_194 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hc2 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_194 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_194 <= _GEN_4328;
      end
    end else begin
      valid_194 <= _GEN_4328;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_195 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hc3 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_195 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_195 <= _GEN_4329;
      end
    end else begin
      valid_195 <= _GEN_4329;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_196 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hc4 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_196 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_196 <= _GEN_4330;
      end
    end else begin
      valid_196 <= _GEN_4330;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_197 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hc5 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_197 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_197 <= _GEN_4331;
      end
    end else begin
      valid_197 <= _GEN_4331;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_198 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hc6 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_198 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_198 <= _GEN_4332;
      end
    end else begin
      valid_198 <= _GEN_4332;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_199 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hc7 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_199 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_199 <= _GEN_4333;
      end
    end else begin
      valid_199 <= _GEN_4333;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_200 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hc8 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_200 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_200 <= _GEN_4334;
      end
    end else begin
      valid_200 <= _GEN_4334;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_201 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hc9 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_201 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_201 <= _GEN_4335;
      end
    end else begin
      valid_201 <= _GEN_4335;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_202 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hca == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_202 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_202 <= _GEN_4336;
      end
    end else begin
      valid_202 <= _GEN_4336;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_203 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hcb == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_203 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_203 <= _GEN_4337;
      end
    end else begin
      valid_203 <= _GEN_4337;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_204 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hcc == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_204 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_204 <= _GEN_4338;
      end
    end else begin
      valid_204 <= _GEN_4338;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_205 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hcd == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_205 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_205 <= _GEN_4339;
      end
    end else begin
      valid_205 <= _GEN_4339;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_206 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hce == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_206 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_206 <= _GEN_4340;
      end
    end else begin
      valid_206 <= _GEN_4340;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_207 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hcf == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_207 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_207 <= _GEN_4341;
      end
    end else begin
      valid_207 <= _GEN_4341;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_208 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hd0 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_208 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_208 <= _GEN_4342;
      end
    end else begin
      valid_208 <= _GEN_4342;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_209 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hd1 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_209 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_209 <= _GEN_4343;
      end
    end else begin
      valid_209 <= _GEN_4343;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_210 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hd2 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_210 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_210 <= _GEN_4344;
      end
    end else begin
      valid_210 <= _GEN_4344;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_211 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hd3 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_211 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_211 <= _GEN_4345;
      end
    end else begin
      valid_211 <= _GEN_4345;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_212 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hd4 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_212 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_212 <= _GEN_4346;
      end
    end else begin
      valid_212 <= _GEN_4346;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_213 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hd5 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_213 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_213 <= _GEN_4347;
      end
    end else begin
      valid_213 <= _GEN_4347;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_214 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hd6 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_214 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_214 <= _GEN_4348;
      end
    end else begin
      valid_214 <= _GEN_4348;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_215 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hd7 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_215 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_215 <= _GEN_4349;
      end
    end else begin
      valid_215 <= _GEN_4349;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_216 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hd8 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_216 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_216 <= _GEN_4350;
      end
    end else begin
      valid_216 <= _GEN_4350;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_217 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hd9 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_217 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_217 <= _GEN_4351;
      end
    end else begin
      valid_217 <= _GEN_4351;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_218 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hda == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_218 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_218 <= _GEN_4352;
      end
    end else begin
      valid_218 <= _GEN_4352;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_219 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hdb == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_219 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_219 <= _GEN_4353;
      end
    end else begin
      valid_219 <= _GEN_4353;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_220 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hdc == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_220 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_220 <= _GEN_4354;
      end
    end else begin
      valid_220 <= _GEN_4354;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_221 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hdd == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_221 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_221 <= _GEN_4355;
      end
    end else begin
      valid_221 <= _GEN_4355;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_222 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hde == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_222 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_222 <= _GEN_4356;
      end
    end else begin
      valid_222 <= _GEN_4356;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_223 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hdf == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_223 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_223 <= _GEN_4357;
      end
    end else begin
      valid_223 <= _GEN_4357;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_224 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'he0 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_224 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_224 <= _GEN_4358;
      end
    end else begin
      valid_224 <= _GEN_4358;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_225 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'he1 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_225 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_225 <= _GEN_4359;
      end
    end else begin
      valid_225 <= _GEN_4359;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_226 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'he2 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_226 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_226 <= _GEN_4360;
      end
    end else begin
      valid_226 <= _GEN_4360;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_227 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'he3 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_227 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_227 <= _GEN_4361;
      end
    end else begin
      valid_227 <= _GEN_4361;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_228 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'he4 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_228 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_228 <= _GEN_4362;
      end
    end else begin
      valid_228 <= _GEN_4362;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_229 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'he5 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_229 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_229 <= _GEN_4363;
      end
    end else begin
      valid_229 <= _GEN_4363;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_230 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'he6 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_230 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_230 <= _GEN_4364;
      end
    end else begin
      valid_230 <= _GEN_4364;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_231 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'he7 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_231 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_231 <= _GEN_4365;
      end
    end else begin
      valid_231 <= _GEN_4365;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_232 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'he8 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_232 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_232 <= _GEN_4366;
      end
    end else begin
      valid_232 <= _GEN_4366;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_233 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'he9 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_233 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_233 <= _GEN_4367;
      end
    end else begin
      valid_233 <= _GEN_4367;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_234 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hea == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_234 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_234 <= _GEN_4368;
      end
    end else begin
      valid_234 <= _GEN_4368;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_235 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'heb == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_235 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_235 <= _GEN_4369;
      end
    end else begin
      valid_235 <= _GEN_4369;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_236 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hec == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_236 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_236 <= _GEN_4370;
      end
    end else begin
      valid_236 <= _GEN_4370;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_237 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hed == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_237 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_237 <= _GEN_4371;
      end
    end else begin
      valid_237 <= _GEN_4371;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_238 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hee == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_238 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_238 <= _GEN_4372;
      end
    end else begin
      valid_238 <= _GEN_4372;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_239 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hef == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_239 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_239 <= _GEN_4373;
      end
    end else begin
      valid_239 <= _GEN_4373;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_240 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hf0 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_240 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_240 <= _GEN_4374;
      end
    end else begin
      valid_240 <= _GEN_4374;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_241 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hf1 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_241 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_241 <= _GEN_4375;
      end
    end else begin
      valid_241 <= _GEN_4375;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_242 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hf2 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_242 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_242 <= _GEN_4376;
      end
    end else begin
      valid_242 <= _GEN_4376;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_243 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hf3 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_243 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_243 <= _GEN_4377;
      end
    end else begin
      valid_243 <= _GEN_4377;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_244 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hf4 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_244 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_244 <= _GEN_4378;
      end
    end else begin
      valid_244 <= _GEN_4378;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_245 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hf5 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_245 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_245 <= _GEN_4379;
      end
    end else begin
      valid_245 <= _GEN_4379;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_246 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hf6 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_246 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_246 <= _GEN_4380;
      end
    end else begin
      valid_246 <= _GEN_4380;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_247 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hf7 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_247 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_247 <= _GEN_4381;
      end
    end else begin
      valid_247 <= _GEN_4381;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_248 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hf8 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_248 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_248 <= _GEN_4382;
      end
    end else begin
      valid_248 <= _GEN_4382;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_249 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hf9 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_249 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_249 <= _GEN_4383;
      end
    end else begin
      valid_249 <= _GEN_4383;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_250 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hfa == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_250 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_250 <= _GEN_4384;
      end
    end else begin
      valid_250 <= _GEN_4384;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_251 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hfb == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_251 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_251 <= _GEN_4385;
      end
    end else begin
      valid_251 <= _GEN_4385;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_252 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hfc == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_252 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_252 <= _GEN_4386;
      end
    end else begin
      valid_252 <= _GEN_4386;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_253 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hfd == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_253 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_253 <= _GEN_4387;
      end
    end else begin
      valid_253 <= _GEN_4387;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_254 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hfe == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_254 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_254 <= _GEN_4388;
      end
    end else begin
      valid_254 <= _GEN_4388;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_255 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'hff == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_255 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_255 <= _GEN_4389;
      end
    end else begin
      valid_255 <= _GEN_4389;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_256 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h100 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_256 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_256 <= _GEN_4390;
      end
    end else begin
      valid_256 <= _GEN_4390;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_257 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h101 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_257 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_257 <= _GEN_4391;
      end
    end else begin
      valid_257 <= _GEN_4391;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_258 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h102 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_258 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_258 <= _GEN_4392;
      end
    end else begin
      valid_258 <= _GEN_4392;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_259 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h103 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_259 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_259 <= _GEN_4393;
      end
    end else begin
      valid_259 <= _GEN_4393;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_260 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h104 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_260 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_260 <= _GEN_4394;
      end
    end else begin
      valid_260 <= _GEN_4394;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_261 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h105 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_261 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_261 <= _GEN_4395;
      end
    end else begin
      valid_261 <= _GEN_4395;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_262 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h106 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_262 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_262 <= _GEN_4396;
      end
    end else begin
      valid_262 <= _GEN_4396;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_263 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h107 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_263 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_263 <= _GEN_4397;
      end
    end else begin
      valid_263 <= _GEN_4397;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_264 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h108 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_264 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_264 <= _GEN_4398;
      end
    end else begin
      valid_264 <= _GEN_4398;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_265 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h109 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_265 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_265 <= _GEN_4399;
      end
    end else begin
      valid_265 <= _GEN_4399;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_266 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h10a == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_266 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_266 <= _GEN_4400;
      end
    end else begin
      valid_266 <= _GEN_4400;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_267 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h10b == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_267 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_267 <= _GEN_4401;
      end
    end else begin
      valid_267 <= _GEN_4401;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_268 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h10c == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_268 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_268 <= _GEN_4402;
      end
    end else begin
      valid_268 <= _GEN_4402;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_269 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h10d == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_269 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_269 <= _GEN_4403;
      end
    end else begin
      valid_269 <= _GEN_4403;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_270 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h10e == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_270 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_270 <= _GEN_4404;
      end
    end else begin
      valid_270 <= _GEN_4404;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_271 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h10f == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_271 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_271 <= _GEN_4405;
      end
    end else begin
      valid_271 <= _GEN_4405;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_272 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h110 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_272 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_272 <= _GEN_4406;
      end
    end else begin
      valid_272 <= _GEN_4406;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_273 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h111 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_273 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_273 <= _GEN_4407;
      end
    end else begin
      valid_273 <= _GEN_4407;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_274 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h112 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_274 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_274 <= _GEN_4408;
      end
    end else begin
      valid_274 <= _GEN_4408;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_275 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h113 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_275 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_275 <= _GEN_4409;
      end
    end else begin
      valid_275 <= _GEN_4409;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_276 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h114 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_276 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_276 <= _GEN_4410;
      end
    end else begin
      valid_276 <= _GEN_4410;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_277 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h115 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_277 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_277 <= _GEN_4411;
      end
    end else begin
      valid_277 <= _GEN_4411;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_278 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h116 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_278 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_278 <= _GEN_4412;
      end
    end else begin
      valid_278 <= _GEN_4412;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_279 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h117 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_279 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_279 <= _GEN_4413;
      end
    end else begin
      valid_279 <= _GEN_4413;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_280 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h118 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_280 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_280 <= _GEN_4414;
      end
    end else begin
      valid_280 <= _GEN_4414;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_281 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h119 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_281 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_281 <= _GEN_4415;
      end
    end else begin
      valid_281 <= _GEN_4415;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_282 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h11a == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_282 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_282 <= _GEN_4416;
      end
    end else begin
      valid_282 <= _GEN_4416;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_283 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h11b == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_283 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_283 <= _GEN_4417;
      end
    end else begin
      valid_283 <= _GEN_4417;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_284 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h11c == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_284 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_284 <= _GEN_4418;
      end
    end else begin
      valid_284 <= _GEN_4418;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_285 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h11d == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_285 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_285 <= _GEN_4419;
      end
    end else begin
      valid_285 <= _GEN_4419;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_286 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h11e == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_286 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_286 <= _GEN_4420;
      end
    end else begin
      valid_286 <= _GEN_4420;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_287 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h11f == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_287 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_287 <= _GEN_4421;
      end
    end else begin
      valid_287 <= _GEN_4421;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_288 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h120 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_288 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_288 <= _GEN_4422;
      end
    end else begin
      valid_288 <= _GEN_4422;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_289 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h121 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_289 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_289 <= _GEN_4423;
      end
    end else begin
      valid_289 <= _GEN_4423;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_290 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h122 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_290 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_290 <= _GEN_4424;
      end
    end else begin
      valid_290 <= _GEN_4424;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_291 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h123 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_291 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_291 <= _GEN_4425;
      end
    end else begin
      valid_291 <= _GEN_4425;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_292 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h124 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_292 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_292 <= _GEN_4426;
      end
    end else begin
      valid_292 <= _GEN_4426;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_293 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h125 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_293 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_293 <= _GEN_4427;
      end
    end else begin
      valid_293 <= _GEN_4427;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_294 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h126 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_294 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_294 <= _GEN_4428;
      end
    end else begin
      valid_294 <= _GEN_4428;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_295 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h127 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_295 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_295 <= _GEN_4429;
      end
    end else begin
      valid_295 <= _GEN_4429;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_296 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h128 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_296 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_296 <= _GEN_4430;
      end
    end else begin
      valid_296 <= _GEN_4430;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_297 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h129 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_297 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_297 <= _GEN_4431;
      end
    end else begin
      valid_297 <= _GEN_4431;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_298 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h12a == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_298 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_298 <= _GEN_4432;
      end
    end else begin
      valid_298 <= _GEN_4432;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_299 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h12b == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_299 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_299 <= _GEN_4433;
      end
    end else begin
      valid_299 <= _GEN_4433;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_300 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h12c == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_300 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_300 <= _GEN_4434;
      end
    end else begin
      valid_300 <= _GEN_4434;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_301 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h12d == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_301 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_301 <= _GEN_4435;
      end
    end else begin
      valid_301 <= _GEN_4435;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_302 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h12e == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_302 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_302 <= _GEN_4436;
      end
    end else begin
      valid_302 <= _GEN_4436;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_303 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h12f == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_303 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_303 <= _GEN_4437;
      end
    end else begin
      valid_303 <= _GEN_4437;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_304 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h130 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_304 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_304 <= _GEN_4438;
      end
    end else begin
      valid_304 <= _GEN_4438;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_305 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h131 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_305 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_305 <= _GEN_4439;
      end
    end else begin
      valid_305 <= _GEN_4439;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_306 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h132 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_306 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_306 <= _GEN_4440;
      end
    end else begin
      valid_306 <= _GEN_4440;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_307 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h133 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_307 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_307 <= _GEN_4441;
      end
    end else begin
      valid_307 <= _GEN_4441;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_308 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h134 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_308 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_308 <= _GEN_4442;
      end
    end else begin
      valid_308 <= _GEN_4442;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_309 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h135 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_309 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_309 <= _GEN_4443;
      end
    end else begin
      valid_309 <= _GEN_4443;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_310 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h136 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_310 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_310 <= _GEN_4444;
      end
    end else begin
      valid_310 <= _GEN_4444;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_311 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h137 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_311 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_311 <= _GEN_4445;
      end
    end else begin
      valid_311 <= _GEN_4445;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_312 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h138 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_312 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_312 <= _GEN_4446;
      end
    end else begin
      valid_312 <= _GEN_4446;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_313 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h139 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_313 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_313 <= _GEN_4447;
      end
    end else begin
      valid_313 <= _GEN_4447;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_314 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h13a == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_314 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_314 <= _GEN_4448;
      end
    end else begin
      valid_314 <= _GEN_4448;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_315 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h13b == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_315 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_315 <= _GEN_4449;
      end
    end else begin
      valid_315 <= _GEN_4449;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_316 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h13c == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_316 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_316 <= _GEN_4450;
      end
    end else begin
      valid_316 <= _GEN_4450;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_317 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h13d == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_317 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_317 <= _GEN_4451;
      end
    end else begin
      valid_317 <= _GEN_4451;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_318 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h13e == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_318 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_318 <= _GEN_4452;
      end
    end else begin
      valid_318 <= _GEN_4452;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_319 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h13f == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_319 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_319 <= _GEN_4453;
      end
    end else begin
      valid_319 <= _GEN_4453;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_320 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h140 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_320 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_320 <= _GEN_4454;
      end
    end else begin
      valid_320 <= _GEN_4454;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_321 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h141 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_321 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_321 <= _GEN_4455;
      end
    end else begin
      valid_321 <= _GEN_4455;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_322 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h142 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_322 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_322 <= _GEN_4456;
      end
    end else begin
      valid_322 <= _GEN_4456;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_323 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h143 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_323 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_323 <= _GEN_4457;
      end
    end else begin
      valid_323 <= _GEN_4457;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_324 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h144 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_324 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_324 <= _GEN_4458;
      end
    end else begin
      valid_324 <= _GEN_4458;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_325 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h145 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_325 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_325 <= _GEN_4459;
      end
    end else begin
      valid_325 <= _GEN_4459;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_326 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h146 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_326 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_326 <= _GEN_4460;
      end
    end else begin
      valid_326 <= _GEN_4460;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_327 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h147 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_327 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_327 <= _GEN_4461;
      end
    end else begin
      valid_327 <= _GEN_4461;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_328 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h148 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_328 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_328 <= _GEN_4462;
      end
    end else begin
      valid_328 <= _GEN_4462;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_329 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h149 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_329 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_329 <= _GEN_4463;
      end
    end else begin
      valid_329 <= _GEN_4463;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_330 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h14a == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_330 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_330 <= _GEN_4464;
      end
    end else begin
      valid_330 <= _GEN_4464;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_331 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h14b == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_331 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_331 <= _GEN_4465;
      end
    end else begin
      valid_331 <= _GEN_4465;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_332 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h14c == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_332 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_332 <= _GEN_4466;
      end
    end else begin
      valid_332 <= _GEN_4466;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_333 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h14d == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_333 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_333 <= _GEN_4467;
      end
    end else begin
      valid_333 <= _GEN_4467;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_334 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h14e == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_334 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_334 <= _GEN_4468;
      end
    end else begin
      valid_334 <= _GEN_4468;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_335 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h14f == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_335 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_335 <= _GEN_4469;
      end
    end else begin
      valid_335 <= _GEN_4469;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_336 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h150 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_336 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_336 <= _GEN_4470;
      end
    end else begin
      valid_336 <= _GEN_4470;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_337 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h151 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_337 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_337 <= _GEN_4471;
      end
    end else begin
      valid_337 <= _GEN_4471;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_338 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h152 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_338 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_338 <= _GEN_4472;
      end
    end else begin
      valid_338 <= _GEN_4472;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_339 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h153 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_339 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_339 <= _GEN_4473;
      end
    end else begin
      valid_339 <= _GEN_4473;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_340 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h154 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_340 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_340 <= _GEN_4474;
      end
    end else begin
      valid_340 <= _GEN_4474;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_341 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h155 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_341 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_341 <= _GEN_4475;
      end
    end else begin
      valid_341 <= _GEN_4475;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_342 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h156 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_342 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_342 <= _GEN_4476;
      end
    end else begin
      valid_342 <= _GEN_4476;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_343 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h157 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_343 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_343 <= _GEN_4477;
      end
    end else begin
      valid_343 <= _GEN_4477;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_344 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h158 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_344 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_344 <= _GEN_4478;
      end
    end else begin
      valid_344 <= _GEN_4478;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_345 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h159 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_345 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_345 <= _GEN_4479;
      end
    end else begin
      valid_345 <= _GEN_4479;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_346 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h15a == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_346 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_346 <= _GEN_4480;
      end
    end else begin
      valid_346 <= _GEN_4480;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_347 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h15b == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_347 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_347 <= _GEN_4481;
      end
    end else begin
      valid_347 <= _GEN_4481;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_348 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h15c == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_348 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_348 <= _GEN_4482;
      end
    end else begin
      valid_348 <= _GEN_4482;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_349 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h15d == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_349 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_349 <= _GEN_4483;
      end
    end else begin
      valid_349 <= _GEN_4483;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_350 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h15e == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_350 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_350 <= _GEN_4484;
      end
    end else begin
      valid_350 <= _GEN_4484;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_351 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h15f == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_351 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_351 <= _GEN_4485;
      end
    end else begin
      valid_351 <= _GEN_4485;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_352 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h160 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_352 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_352 <= _GEN_4486;
      end
    end else begin
      valid_352 <= _GEN_4486;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_353 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h161 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_353 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_353 <= _GEN_4487;
      end
    end else begin
      valid_353 <= _GEN_4487;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_354 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h162 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_354 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_354 <= _GEN_4488;
      end
    end else begin
      valid_354 <= _GEN_4488;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_355 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h163 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_355 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_355 <= _GEN_4489;
      end
    end else begin
      valid_355 <= _GEN_4489;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_356 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h164 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_356 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_356 <= _GEN_4490;
      end
    end else begin
      valid_356 <= _GEN_4490;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_357 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h165 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_357 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_357 <= _GEN_4491;
      end
    end else begin
      valid_357 <= _GEN_4491;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_358 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h166 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_358 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_358 <= _GEN_4492;
      end
    end else begin
      valid_358 <= _GEN_4492;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_359 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h167 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_359 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_359 <= _GEN_4493;
      end
    end else begin
      valid_359 <= _GEN_4493;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_360 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h168 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_360 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_360 <= _GEN_4494;
      end
    end else begin
      valid_360 <= _GEN_4494;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_361 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h169 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_361 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_361 <= _GEN_4495;
      end
    end else begin
      valid_361 <= _GEN_4495;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_362 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h16a == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_362 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_362 <= _GEN_4496;
      end
    end else begin
      valid_362 <= _GEN_4496;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_363 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h16b == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_363 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_363 <= _GEN_4497;
      end
    end else begin
      valid_363 <= _GEN_4497;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_364 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h16c == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_364 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_364 <= _GEN_4498;
      end
    end else begin
      valid_364 <= _GEN_4498;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_365 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h16d == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_365 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_365 <= _GEN_4499;
      end
    end else begin
      valid_365 <= _GEN_4499;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_366 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h16e == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_366 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_366 <= _GEN_4500;
      end
    end else begin
      valid_366 <= _GEN_4500;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_367 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h16f == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_367 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_367 <= _GEN_4501;
      end
    end else begin
      valid_367 <= _GEN_4501;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_368 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h170 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_368 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_368 <= _GEN_4502;
      end
    end else begin
      valid_368 <= _GEN_4502;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_369 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h171 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_369 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_369 <= _GEN_4503;
      end
    end else begin
      valid_369 <= _GEN_4503;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_370 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h172 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_370 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_370 <= _GEN_4504;
      end
    end else begin
      valid_370 <= _GEN_4504;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_371 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h173 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_371 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_371 <= _GEN_4505;
      end
    end else begin
      valid_371 <= _GEN_4505;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_372 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h174 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_372 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_372 <= _GEN_4506;
      end
    end else begin
      valid_372 <= _GEN_4506;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_373 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h175 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_373 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_373 <= _GEN_4507;
      end
    end else begin
      valid_373 <= _GEN_4507;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_374 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h176 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_374 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_374 <= _GEN_4508;
      end
    end else begin
      valid_374 <= _GEN_4508;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_375 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h177 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_375 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_375 <= _GEN_4509;
      end
    end else begin
      valid_375 <= _GEN_4509;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_376 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h178 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_376 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_376 <= _GEN_4510;
      end
    end else begin
      valid_376 <= _GEN_4510;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_377 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h179 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_377 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_377 <= _GEN_4511;
      end
    end else begin
      valid_377 <= _GEN_4511;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_378 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h17a == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_378 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_378 <= _GEN_4512;
      end
    end else begin
      valid_378 <= _GEN_4512;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_379 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h17b == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_379 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_379 <= _GEN_4513;
      end
    end else begin
      valid_379 <= _GEN_4513;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_380 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h17c == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_380 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_380 <= _GEN_4514;
      end
    end else begin
      valid_380 <= _GEN_4514;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_381 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h17d == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_381 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_381 <= _GEN_4515;
      end
    end else begin
      valid_381 <= _GEN_4515;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_382 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h17e == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_382 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_382 <= _GEN_4516;
      end
    end else begin
      valid_382 <= _GEN_4516;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_383 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h17f == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_383 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_383 <= _GEN_4517;
      end
    end else begin
      valid_383 <= _GEN_4517;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_384 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h180 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_384 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_384 <= _GEN_4518;
      end
    end else begin
      valid_384 <= _GEN_4518;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_385 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h181 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_385 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_385 <= _GEN_4519;
      end
    end else begin
      valid_385 <= _GEN_4519;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_386 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h182 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_386 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_386 <= _GEN_4520;
      end
    end else begin
      valid_386 <= _GEN_4520;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_387 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h183 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_387 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_387 <= _GEN_4521;
      end
    end else begin
      valid_387 <= _GEN_4521;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_388 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h184 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_388 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_388 <= _GEN_4522;
      end
    end else begin
      valid_388 <= _GEN_4522;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_389 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h185 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_389 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_389 <= _GEN_4523;
      end
    end else begin
      valid_389 <= _GEN_4523;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_390 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h186 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_390 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_390 <= _GEN_4524;
      end
    end else begin
      valid_390 <= _GEN_4524;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_391 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h187 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_391 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_391 <= _GEN_4525;
      end
    end else begin
      valid_391 <= _GEN_4525;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_392 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h188 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_392 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_392 <= _GEN_4526;
      end
    end else begin
      valid_392 <= _GEN_4526;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_393 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h189 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_393 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_393 <= _GEN_4527;
      end
    end else begin
      valid_393 <= _GEN_4527;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_394 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h18a == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_394 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_394 <= _GEN_4528;
      end
    end else begin
      valid_394 <= _GEN_4528;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_395 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h18b == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_395 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_395 <= _GEN_4529;
      end
    end else begin
      valid_395 <= _GEN_4529;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_396 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h18c == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_396 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_396 <= _GEN_4530;
      end
    end else begin
      valid_396 <= _GEN_4530;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_397 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h18d == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_397 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_397 <= _GEN_4531;
      end
    end else begin
      valid_397 <= _GEN_4531;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_398 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h18e == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_398 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_398 <= _GEN_4532;
      end
    end else begin
      valid_398 <= _GEN_4532;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_399 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h18f == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_399 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_399 <= _GEN_4533;
      end
    end else begin
      valid_399 <= _GEN_4533;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_400 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h190 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_400 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_400 <= _GEN_4534;
      end
    end else begin
      valid_400 <= _GEN_4534;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_401 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h191 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_401 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_401 <= _GEN_4535;
      end
    end else begin
      valid_401 <= _GEN_4535;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_402 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h192 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_402 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_402 <= _GEN_4536;
      end
    end else begin
      valid_402 <= _GEN_4536;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_403 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h193 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_403 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_403 <= _GEN_4537;
      end
    end else begin
      valid_403 <= _GEN_4537;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_404 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h194 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_404 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_404 <= _GEN_4538;
      end
    end else begin
      valid_404 <= _GEN_4538;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_405 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h195 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_405 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_405 <= _GEN_4539;
      end
    end else begin
      valid_405 <= _GEN_4539;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_406 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h196 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_406 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_406 <= _GEN_4540;
      end
    end else begin
      valid_406 <= _GEN_4540;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_407 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h197 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_407 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_407 <= _GEN_4541;
      end
    end else begin
      valid_407 <= _GEN_4541;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_408 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h198 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_408 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_408 <= _GEN_4542;
      end
    end else begin
      valid_408 <= _GEN_4542;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_409 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h199 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_409 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_409 <= _GEN_4543;
      end
    end else begin
      valid_409 <= _GEN_4543;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_410 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h19a == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_410 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_410 <= _GEN_4544;
      end
    end else begin
      valid_410 <= _GEN_4544;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_411 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h19b == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_411 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_411 <= _GEN_4545;
      end
    end else begin
      valid_411 <= _GEN_4545;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_412 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h19c == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_412 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_412 <= _GEN_4546;
      end
    end else begin
      valid_412 <= _GEN_4546;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_413 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h19d == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_413 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_413 <= _GEN_4547;
      end
    end else begin
      valid_413 <= _GEN_4547;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_414 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h19e == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_414 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_414 <= _GEN_4548;
      end
    end else begin
      valid_414 <= _GEN_4548;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_415 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h19f == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_415 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_415 <= _GEN_4549;
      end
    end else begin
      valid_415 <= _GEN_4549;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_416 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1a0 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_416 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_416 <= _GEN_4550;
      end
    end else begin
      valid_416 <= _GEN_4550;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_417 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1a1 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_417 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_417 <= _GEN_4551;
      end
    end else begin
      valid_417 <= _GEN_4551;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_418 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1a2 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_418 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_418 <= _GEN_4552;
      end
    end else begin
      valid_418 <= _GEN_4552;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_419 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1a3 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_419 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_419 <= _GEN_4553;
      end
    end else begin
      valid_419 <= _GEN_4553;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_420 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1a4 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_420 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_420 <= _GEN_4554;
      end
    end else begin
      valid_420 <= _GEN_4554;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_421 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1a5 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_421 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_421 <= _GEN_4555;
      end
    end else begin
      valid_421 <= _GEN_4555;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_422 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1a6 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_422 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_422 <= _GEN_4556;
      end
    end else begin
      valid_422 <= _GEN_4556;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_423 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1a7 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_423 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_423 <= _GEN_4557;
      end
    end else begin
      valid_423 <= _GEN_4557;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_424 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1a8 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_424 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_424 <= _GEN_4558;
      end
    end else begin
      valid_424 <= _GEN_4558;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_425 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1a9 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_425 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_425 <= _GEN_4559;
      end
    end else begin
      valid_425 <= _GEN_4559;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_426 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1aa == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_426 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_426 <= _GEN_4560;
      end
    end else begin
      valid_426 <= _GEN_4560;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_427 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1ab == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_427 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_427 <= _GEN_4561;
      end
    end else begin
      valid_427 <= _GEN_4561;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_428 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1ac == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_428 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_428 <= _GEN_4562;
      end
    end else begin
      valid_428 <= _GEN_4562;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_429 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1ad == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_429 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_429 <= _GEN_4563;
      end
    end else begin
      valid_429 <= _GEN_4563;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_430 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1ae == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_430 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_430 <= _GEN_4564;
      end
    end else begin
      valid_430 <= _GEN_4564;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_431 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1af == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_431 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_431 <= _GEN_4565;
      end
    end else begin
      valid_431 <= _GEN_4565;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_432 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1b0 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_432 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_432 <= _GEN_4566;
      end
    end else begin
      valid_432 <= _GEN_4566;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_433 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1b1 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_433 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_433 <= _GEN_4567;
      end
    end else begin
      valid_433 <= _GEN_4567;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_434 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1b2 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_434 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_434 <= _GEN_4568;
      end
    end else begin
      valid_434 <= _GEN_4568;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_435 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1b3 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_435 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_435 <= _GEN_4569;
      end
    end else begin
      valid_435 <= _GEN_4569;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_436 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1b4 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_436 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_436 <= _GEN_4570;
      end
    end else begin
      valid_436 <= _GEN_4570;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_437 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1b5 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_437 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_437 <= _GEN_4571;
      end
    end else begin
      valid_437 <= _GEN_4571;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_438 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1b6 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_438 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_438 <= _GEN_4572;
      end
    end else begin
      valid_438 <= _GEN_4572;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_439 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1b7 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_439 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_439 <= _GEN_4573;
      end
    end else begin
      valid_439 <= _GEN_4573;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_440 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1b8 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_440 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_440 <= _GEN_4574;
      end
    end else begin
      valid_440 <= _GEN_4574;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_441 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1b9 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_441 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_441 <= _GEN_4575;
      end
    end else begin
      valid_441 <= _GEN_4575;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_442 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1ba == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_442 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_442 <= _GEN_4576;
      end
    end else begin
      valid_442 <= _GEN_4576;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_443 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1bb == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_443 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_443 <= _GEN_4577;
      end
    end else begin
      valid_443 <= _GEN_4577;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_444 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1bc == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_444 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_444 <= _GEN_4578;
      end
    end else begin
      valid_444 <= _GEN_4578;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_445 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1bd == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_445 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_445 <= _GEN_4579;
      end
    end else begin
      valid_445 <= _GEN_4579;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_446 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1be == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_446 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_446 <= _GEN_4580;
      end
    end else begin
      valid_446 <= _GEN_4580;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_447 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1bf == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_447 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_447 <= _GEN_4581;
      end
    end else begin
      valid_447 <= _GEN_4581;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_448 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1c0 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_448 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_448 <= _GEN_4582;
      end
    end else begin
      valid_448 <= _GEN_4582;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_449 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1c1 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_449 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_449 <= _GEN_4583;
      end
    end else begin
      valid_449 <= _GEN_4583;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_450 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1c2 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_450 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_450 <= _GEN_4584;
      end
    end else begin
      valid_450 <= _GEN_4584;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_451 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1c3 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_451 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_451 <= _GEN_4585;
      end
    end else begin
      valid_451 <= _GEN_4585;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_452 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1c4 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_452 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_452 <= _GEN_4586;
      end
    end else begin
      valid_452 <= _GEN_4586;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_453 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1c5 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_453 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_453 <= _GEN_4587;
      end
    end else begin
      valid_453 <= _GEN_4587;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_454 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1c6 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_454 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_454 <= _GEN_4588;
      end
    end else begin
      valid_454 <= _GEN_4588;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_455 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1c7 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_455 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_455 <= _GEN_4589;
      end
    end else begin
      valid_455 <= _GEN_4589;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_456 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1c8 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_456 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_456 <= _GEN_4590;
      end
    end else begin
      valid_456 <= _GEN_4590;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_457 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1c9 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_457 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_457 <= _GEN_4591;
      end
    end else begin
      valid_457 <= _GEN_4591;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_458 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1ca == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_458 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_458 <= _GEN_4592;
      end
    end else begin
      valid_458 <= _GEN_4592;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_459 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1cb == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_459 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_459 <= _GEN_4593;
      end
    end else begin
      valid_459 <= _GEN_4593;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_460 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1cc == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_460 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_460 <= _GEN_4594;
      end
    end else begin
      valid_460 <= _GEN_4594;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_461 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1cd == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_461 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_461 <= _GEN_4595;
      end
    end else begin
      valid_461 <= _GEN_4595;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_462 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1ce == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_462 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_462 <= _GEN_4596;
      end
    end else begin
      valid_462 <= _GEN_4596;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_463 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1cf == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_463 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_463 <= _GEN_4597;
      end
    end else begin
      valid_463 <= _GEN_4597;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_464 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1d0 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_464 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_464 <= _GEN_4598;
      end
    end else begin
      valid_464 <= _GEN_4598;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_465 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1d1 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_465 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_465 <= _GEN_4599;
      end
    end else begin
      valid_465 <= _GEN_4599;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_466 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1d2 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_466 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_466 <= _GEN_4600;
      end
    end else begin
      valid_466 <= _GEN_4600;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_467 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1d3 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_467 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_467 <= _GEN_4601;
      end
    end else begin
      valid_467 <= _GEN_4601;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_468 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1d4 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_468 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_468 <= _GEN_4602;
      end
    end else begin
      valid_468 <= _GEN_4602;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_469 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1d5 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_469 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_469 <= _GEN_4603;
      end
    end else begin
      valid_469 <= _GEN_4603;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_470 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1d6 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_470 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_470 <= _GEN_4604;
      end
    end else begin
      valid_470 <= _GEN_4604;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_471 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1d7 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_471 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_471 <= _GEN_4605;
      end
    end else begin
      valid_471 <= _GEN_4605;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_472 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1d8 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_472 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_472 <= _GEN_4606;
      end
    end else begin
      valid_472 <= _GEN_4606;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_473 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1d9 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_473 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_473 <= _GEN_4607;
      end
    end else begin
      valid_473 <= _GEN_4607;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_474 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1da == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_474 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_474 <= _GEN_4608;
      end
    end else begin
      valid_474 <= _GEN_4608;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_475 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1db == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_475 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_475 <= _GEN_4609;
      end
    end else begin
      valid_475 <= _GEN_4609;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_476 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1dc == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_476 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_476 <= _GEN_4610;
      end
    end else begin
      valid_476 <= _GEN_4610;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_477 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1dd == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_477 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_477 <= _GEN_4611;
      end
    end else begin
      valid_477 <= _GEN_4611;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_478 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1de == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_478 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_478 <= _GEN_4612;
      end
    end else begin
      valid_478 <= _GEN_4612;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_479 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1df == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_479 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_479 <= _GEN_4613;
      end
    end else begin
      valid_479 <= _GEN_4613;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_480 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1e0 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_480 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_480 <= _GEN_4614;
      end
    end else begin
      valid_480 <= _GEN_4614;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_481 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1e1 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_481 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_481 <= _GEN_4615;
      end
    end else begin
      valid_481 <= _GEN_4615;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_482 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1e2 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_482 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_482 <= _GEN_4616;
      end
    end else begin
      valid_482 <= _GEN_4616;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_483 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1e3 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_483 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_483 <= _GEN_4617;
      end
    end else begin
      valid_483 <= _GEN_4617;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_484 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1e4 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_484 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_484 <= _GEN_4618;
      end
    end else begin
      valid_484 <= _GEN_4618;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_485 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1e5 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_485 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_485 <= _GEN_4619;
      end
    end else begin
      valid_485 <= _GEN_4619;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_486 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1e6 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_486 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_486 <= _GEN_4620;
      end
    end else begin
      valid_486 <= _GEN_4620;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_487 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1e7 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_487 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_487 <= _GEN_4621;
      end
    end else begin
      valid_487 <= _GEN_4621;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_488 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1e8 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_488 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_488 <= _GEN_4622;
      end
    end else begin
      valid_488 <= _GEN_4622;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_489 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1e9 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_489 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_489 <= _GEN_4623;
      end
    end else begin
      valid_489 <= _GEN_4623;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_490 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1ea == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_490 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_490 <= _GEN_4624;
      end
    end else begin
      valid_490 <= _GEN_4624;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_491 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1eb == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_491 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_491 <= _GEN_4625;
      end
    end else begin
      valid_491 <= _GEN_4625;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_492 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1ec == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_492 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_492 <= _GEN_4626;
      end
    end else begin
      valid_492 <= _GEN_4626;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_493 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1ed == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_493 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_493 <= _GEN_4627;
      end
    end else begin
      valid_493 <= _GEN_4627;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_494 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1ee == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_494 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_494 <= _GEN_4628;
      end
    end else begin
      valid_494 <= _GEN_4628;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_495 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1ef == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_495 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_495 <= _GEN_4629;
      end
    end else begin
      valid_495 <= _GEN_4629;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_496 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1f0 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_496 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_496 <= _GEN_4630;
      end
    end else begin
      valid_496 <= _GEN_4630;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_497 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1f1 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_497 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_497 <= _GEN_4631;
      end
    end else begin
      valid_497 <= _GEN_4631;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_498 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1f2 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_498 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_498 <= _GEN_4632;
      end
    end else begin
      valid_498 <= _GEN_4632;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_499 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1f3 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_499 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_499 <= _GEN_4633;
      end
    end else begin
      valid_499 <= _GEN_4633;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_500 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1f4 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_500 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_500 <= _GEN_4634;
      end
    end else begin
      valid_500 <= _GEN_4634;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_501 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1f5 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_501 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_501 <= _GEN_4635;
      end
    end else begin
      valid_501 <= _GEN_4635;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_502 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1f6 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_502 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_502 <= _GEN_4636;
      end
    end else begin
      valid_502 <= _GEN_4636;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_503 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1f7 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_503 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_503 <= _GEN_4637;
      end
    end else begin
      valid_503 <= _GEN_4637;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_504 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1f8 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_504 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_504 <= _GEN_4638;
      end
    end else begin
      valid_504 <= _GEN_4638;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_505 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1f9 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_505 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_505 <= _GEN_4639;
      end
    end else begin
      valid_505 <= _GEN_4639;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_506 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1fa == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_506 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_506 <= _GEN_4640;
      end
    end else begin
      valid_506 <= _GEN_4640;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_507 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1fb == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_507 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_507 <= _GEN_4641;
      end
    end else begin
      valid_507 <= _GEN_4641;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_508 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1fc == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_508 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_508 <= _GEN_4642;
      end
    end else begin
      valid_508 <= _GEN_4642;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_509 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1fd == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_509 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_509 <= _GEN_4643;
      end
    end else begin
      valid_509 <= _GEN_4643;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_510 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1fe == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_510 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_510 <= _GEN_4644;
      end
    end else begin
      valid_510 <= _GEN_4644;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_511 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h1ff == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_511 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_511 <= _GEN_4645;
      end
    end else begin
      valid_511 <= _GEN_4645;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_512 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h200 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_512 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_512 <= _GEN_4646;
      end
    end else begin
      valid_512 <= _GEN_4646;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_513 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h201 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_513 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_513 <= _GEN_4647;
      end
    end else begin
      valid_513 <= _GEN_4647;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_514 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h202 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_514 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_514 <= _GEN_4648;
      end
    end else begin
      valid_514 <= _GEN_4648;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_515 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h203 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_515 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_515 <= _GEN_4649;
      end
    end else begin
      valid_515 <= _GEN_4649;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_516 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h204 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_516 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_516 <= _GEN_4650;
      end
    end else begin
      valid_516 <= _GEN_4650;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_517 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h205 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_517 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_517 <= _GEN_4651;
      end
    end else begin
      valid_517 <= _GEN_4651;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_518 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h206 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_518 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_518 <= _GEN_4652;
      end
    end else begin
      valid_518 <= _GEN_4652;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_519 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h207 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_519 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_519 <= _GEN_4653;
      end
    end else begin
      valid_519 <= _GEN_4653;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_520 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h208 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_520 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_520 <= _GEN_4654;
      end
    end else begin
      valid_520 <= _GEN_4654;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_521 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h209 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_521 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_521 <= _GEN_4655;
      end
    end else begin
      valid_521 <= _GEN_4655;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_522 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h20a == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_522 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_522 <= _GEN_4656;
      end
    end else begin
      valid_522 <= _GEN_4656;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_523 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h20b == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_523 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_523 <= _GEN_4657;
      end
    end else begin
      valid_523 <= _GEN_4657;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_524 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h20c == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_524 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_524 <= _GEN_4658;
      end
    end else begin
      valid_524 <= _GEN_4658;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_525 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h20d == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_525 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_525 <= _GEN_4659;
      end
    end else begin
      valid_525 <= _GEN_4659;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_526 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h20e == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_526 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_526 <= _GEN_4660;
      end
    end else begin
      valid_526 <= _GEN_4660;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_527 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h20f == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_527 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_527 <= _GEN_4661;
      end
    end else begin
      valid_527 <= _GEN_4661;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_528 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h210 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_528 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_528 <= _GEN_4662;
      end
    end else begin
      valid_528 <= _GEN_4662;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_529 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h211 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_529 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_529 <= _GEN_4663;
      end
    end else begin
      valid_529 <= _GEN_4663;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_530 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h212 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_530 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_530 <= _GEN_4664;
      end
    end else begin
      valid_530 <= _GEN_4664;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_531 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h213 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_531 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_531 <= _GEN_4665;
      end
    end else begin
      valid_531 <= _GEN_4665;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_532 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h214 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_532 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_532 <= _GEN_4666;
      end
    end else begin
      valid_532 <= _GEN_4666;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_533 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h215 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_533 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_533 <= _GEN_4667;
      end
    end else begin
      valid_533 <= _GEN_4667;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_534 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h216 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_534 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_534 <= _GEN_4668;
      end
    end else begin
      valid_534 <= _GEN_4668;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_535 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h217 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_535 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_535 <= _GEN_4669;
      end
    end else begin
      valid_535 <= _GEN_4669;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_536 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h218 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_536 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_536 <= _GEN_4670;
      end
    end else begin
      valid_536 <= _GEN_4670;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_537 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h219 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_537 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_537 <= _GEN_4671;
      end
    end else begin
      valid_537 <= _GEN_4671;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_538 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h21a == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_538 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_538 <= _GEN_4672;
      end
    end else begin
      valid_538 <= _GEN_4672;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_539 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h21b == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_539 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_539 <= _GEN_4673;
      end
    end else begin
      valid_539 <= _GEN_4673;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_540 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h21c == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_540 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_540 <= _GEN_4674;
      end
    end else begin
      valid_540 <= _GEN_4674;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_541 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h21d == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_541 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_541 <= _GEN_4675;
      end
    end else begin
      valid_541 <= _GEN_4675;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_542 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h21e == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_542 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_542 <= _GEN_4676;
      end
    end else begin
      valid_542 <= _GEN_4676;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_543 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h21f == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_543 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_543 <= _GEN_4677;
      end
    end else begin
      valid_543 <= _GEN_4677;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_544 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h220 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_544 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_544 <= _GEN_4678;
      end
    end else begin
      valid_544 <= _GEN_4678;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_545 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h221 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_545 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_545 <= _GEN_4679;
      end
    end else begin
      valid_545 <= _GEN_4679;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_546 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h222 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_546 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_546 <= _GEN_4680;
      end
    end else begin
      valid_546 <= _GEN_4680;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_547 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h223 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_547 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_547 <= _GEN_4681;
      end
    end else begin
      valid_547 <= _GEN_4681;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_548 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h224 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_548 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_548 <= _GEN_4682;
      end
    end else begin
      valid_548 <= _GEN_4682;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_549 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h225 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_549 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_549 <= _GEN_4683;
      end
    end else begin
      valid_549 <= _GEN_4683;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_550 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h226 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_550 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_550 <= _GEN_4684;
      end
    end else begin
      valid_550 <= _GEN_4684;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_551 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h227 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_551 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_551 <= _GEN_4685;
      end
    end else begin
      valid_551 <= _GEN_4685;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_552 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h228 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_552 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_552 <= _GEN_4686;
      end
    end else begin
      valid_552 <= _GEN_4686;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_553 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h229 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_553 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_553 <= _GEN_4687;
      end
    end else begin
      valid_553 <= _GEN_4687;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_554 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h22a == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_554 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_554 <= _GEN_4688;
      end
    end else begin
      valid_554 <= _GEN_4688;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_555 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h22b == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_555 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_555 <= _GEN_4689;
      end
    end else begin
      valid_555 <= _GEN_4689;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_556 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h22c == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_556 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_556 <= _GEN_4690;
      end
    end else begin
      valid_556 <= _GEN_4690;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_557 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h22d == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_557 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_557 <= _GEN_4691;
      end
    end else begin
      valid_557 <= _GEN_4691;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_558 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h22e == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_558 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_558 <= _GEN_4692;
      end
    end else begin
      valid_558 <= _GEN_4692;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_559 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h22f == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_559 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_559 <= _GEN_4693;
      end
    end else begin
      valid_559 <= _GEN_4693;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_560 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h230 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_560 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_560 <= _GEN_4694;
      end
    end else begin
      valid_560 <= _GEN_4694;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_561 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h231 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_561 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_561 <= _GEN_4695;
      end
    end else begin
      valid_561 <= _GEN_4695;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_562 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h232 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_562 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_562 <= _GEN_4696;
      end
    end else begin
      valid_562 <= _GEN_4696;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_563 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h233 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_563 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_563 <= _GEN_4697;
      end
    end else begin
      valid_563 <= _GEN_4697;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_564 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h234 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_564 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_564 <= _GEN_4698;
      end
    end else begin
      valid_564 <= _GEN_4698;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_565 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h235 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_565 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_565 <= _GEN_4699;
      end
    end else begin
      valid_565 <= _GEN_4699;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_566 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h236 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_566 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_566 <= _GEN_4700;
      end
    end else begin
      valid_566 <= _GEN_4700;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_567 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h237 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_567 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_567 <= _GEN_4701;
      end
    end else begin
      valid_567 <= _GEN_4701;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_568 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h238 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_568 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_568 <= _GEN_4702;
      end
    end else begin
      valid_568 <= _GEN_4702;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_569 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h239 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_569 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_569 <= _GEN_4703;
      end
    end else begin
      valid_569 <= _GEN_4703;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_570 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h23a == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_570 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_570 <= _GEN_4704;
      end
    end else begin
      valid_570 <= _GEN_4704;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_571 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h23b == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_571 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_571 <= _GEN_4705;
      end
    end else begin
      valid_571 <= _GEN_4705;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_572 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h23c == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_572 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_572 <= _GEN_4706;
      end
    end else begin
      valid_572 <= _GEN_4706;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_573 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h23d == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_573 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_573 <= _GEN_4707;
      end
    end else begin
      valid_573 <= _GEN_4707;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_574 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h23e == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_574 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_574 <= _GEN_4708;
      end
    end else begin
      valid_574 <= _GEN_4708;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_575 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h23f == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_575 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_575 <= _GEN_4709;
      end
    end else begin
      valid_575 <= _GEN_4709;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_576 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h240 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_576 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_576 <= _GEN_4710;
      end
    end else begin
      valid_576 <= _GEN_4710;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_577 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h241 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_577 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_577 <= _GEN_4711;
      end
    end else begin
      valid_577 <= _GEN_4711;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_578 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h242 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_578 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_578 <= _GEN_4712;
      end
    end else begin
      valid_578 <= _GEN_4712;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_579 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h243 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_579 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_579 <= _GEN_4713;
      end
    end else begin
      valid_579 <= _GEN_4713;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_580 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h244 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_580 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_580 <= _GEN_4714;
      end
    end else begin
      valid_580 <= _GEN_4714;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_581 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h245 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_581 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_581 <= _GEN_4715;
      end
    end else begin
      valid_581 <= _GEN_4715;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_582 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h246 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_582 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_582 <= _GEN_4716;
      end
    end else begin
      valid_582 <= _GEN_4716;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_583 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h247 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_583 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_583 <= _GEN_4717;
      end
    end else begin
      valid_583 <= _GEN_4717;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_584 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h248 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_584 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_584 <= _GEN_4718;
      end
    end else begin
      valid_584 <= _GEN_4718;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_585 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h249 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_585 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_585 <= _GEN_4719;
      end
    end else begin
      valid_585 <= _GEN_4719;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_586 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h24a == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_586 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_586 <= _GEN_4720;
      end
    end else begin
      valid_586 <= _GEN_4720;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_587 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h24b == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_587 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_587 <= _GEN_4721;
      end
    end else begin
      valid_587 <= _GEN_4721;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_588 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h24c == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_588 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_588 <= _GEN_4722;
      end
    end else begin
      valid_588 <= _GEN_4722;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_589 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h24d == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_589 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_589 <= _GEN_4723;
      end
    end else begin
      valid_589 <= _GEN_4723;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_590 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h24e == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_590 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_590 <= _GEN_4724;
      end
    end else begin
      valid_590 <= _GEN_4724;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_591 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h24f == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_591 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_591 <= _GEN_4725;
      end
    end else begin
      valid_591 <= _GEN_4725;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_592 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h250 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_592 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_592 <= _GEN_4726;
      end
    end else begin
      valid_592 <= _GEN_4726;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_593 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h251 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_593 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_593 <= _GEN_4727;
      end
    end else begin
      valid_593 <= _GEN_4727;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_594 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h252 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_594 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_594 <= _GEN_4728;
      end
    end else begin
      valid_594 <= _GEN_4728;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_595 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h253 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_595 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_595 <= _GEN_4729;
      end
    end else begin
      valid_595 <= _GEN_4729;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_596 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h254 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_596 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_596 <= _GEN_4730;
      end
    end else begin
      valid_596 <= _GEN_4730;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_597 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h255 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_597 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_597 <= _GEN_4731;
      end
    end else begin
      valid_597 <= _GEN_4731;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_598 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h256 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_598 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_598 <= _GEN_4732;
      end
    end else begin
      valid_598 <= _GEN_4732;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_599 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h257 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_599 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_599 <= _GEN_4733;
      end
    end else begin
      valid_599 <= _GEN_4733;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_600 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h258 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_600 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_600 <= _GEN_4734;
      end
    end else begin
      valid_600 <= _GEN_4734;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_601 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h259 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_601 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_601 <= _GEN_4735;
      end
    end else begin
      valid_601 <= _GEN_4735;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_602 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h25a == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_602 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_602 <= _GEN_4736;
      end
    end else begin
      valid_602 <= _GEN_4736;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_603 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h25b == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_603 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_603 <= _GEN_4737;
      end
    end else begin
      valid_603 <= _GEN_4737;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_604 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h25c == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_604 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_604 <= _GEN_4738;
      end
    end else begin
      valid_604 <= _GEN_4738;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_605 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h25d == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_605 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_605 <= _GEN_4739;
      end
    end else begin
      valid_605 <= _GEN_4739;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_606 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h25e == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_606 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_606 <= _GEN_4740;
      end
    end else begin
      valid_606 <= _GEN_4740;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_607 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h25f == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_607 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_607 <= _GEN_4741;
      end
    end else begin
      valid_607 <= _GEN_4741;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_608 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h260 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_608 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_608 <= _GEN_4742;
      end
    end else begin
      valid_608 <= _GEN_4742;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_609 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h261 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_609 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_609 <= _GEN_4743;
      end
    end else begin
      valid_609 <= _GEN_4743;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_610 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h262 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_610 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_610 <= _GEN_4744;
      end
    end else begin
      valid_610 <= _GEN_4744;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_611 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h263 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_611 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_611 <= _GEN_4745;
      end
    end else begin
      valid_611 <= _GEN_4745;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_612 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h264 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_612 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_612 <= _GEN_4746;
      end
    end else begin
      valid_612 <= _GEN_4746;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_613 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h265 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_613 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_613 <= _GEN_4747;
      end
    end else begin
      valid_613 <= _GEN_4747;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_614 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h266 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_614 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_614 <= _GEN_4748;
      end
    end else begin
      valid_614 <= _GEN_4748;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_615 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h267 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_615 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_615 <= _GEN_4749;
      end
    end else begin
      valid_615 <= _GEN_4749;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_616 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h268 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_616 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_616 <= _GEN_4750;
      end
    end else begin
      valid_616 <= _GEN_4750;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_617 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h269 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_617 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_617 <= _GEN_4751;
      end
    end else begin
      valid_617 <= _GEN_4751;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_618 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h26a == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_618 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_618 <= _GEN_4752;
      end
    end else begin
      valid_618 <= _GEN_4752;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_619 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h26b == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_619 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_619 <= _GEN_4753;
      end
    end else begin
      valid_619 <= _GEN_4753;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_620 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h26c == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_620 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_620 <= _GEN_4754;
      end
    end else begin
      valid_620 <= _GEN_4754;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_621 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h26d == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_621 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_621 <= _GEN_4755;
      end
    end else begin
      valid_621 <= _GEN_4755;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_622 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h26e == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_622 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_622 <= _GEN_4756;
      end
    end else begin
      valid_622 <= _GEN_4756;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_623 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h26f == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_623 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_623 <= _GEN_4757;
      end
    end else begin
      valid_623 <= _GEN_4757;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_624 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h270 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_624 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_624 <= _GEN_4758;
      end
    end else begin
      valid_624 <= _GEN_4758;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_625 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h271 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_625 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_625 <= _GEN_4759;
      end
    end else begin
      valid_625 <= _GEN_4759;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_626 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h272 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_626 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_626 <= _GEN_4760;
      end
    end else begin
      valid_626 <= _GEN_4760;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_627 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h273 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_627 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_627 <= _GEN_4761;
      end
    end else begin
      valid_627 <= _GEN_4761;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_628 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h274 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_628 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_628 <= _GEN_4762;
      end
    end else begin
      valid_628 <= _GEN_4762;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_629 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h275 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_629 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_629 <= _GEN_4763;
      end
    end else begin
      valid_629 <= _GEN_4763;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_630 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h276 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_630 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_630 <= _GEN_4764;
      end
    end else begin
      valid_630 <= _GEN_4764;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_631 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h277 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_631 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_631 <= _GEN_4765;
      end
    end else begin
      valid_631 <= _GEN_4765;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_632 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h278 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_632 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_632 <= _GEN_4766;
      end
    end else begin
      valid_632 <= _GEN_4766;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_633 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h279 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_633 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_633 <= _GEN_4767;
      end
    end else begin
      valid_633 <= _GEN_4767;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_634 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h27a == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_634 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_634 <= _GEN_4768;
      end
    end else begin
      valid_634 <= _GEN_4768;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_635 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h27b == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_635 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_635 <= _GEN_4769;
      end
    end else begin
      valid_635 <= _GEN_4769;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_636 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h27c == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_636 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_636 <= _GEN_4770;
      end
    end else begin
      valid_636 <= _GEN_4770;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_637 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h27d == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_637 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_637 <= _GEN_4771;
      end
    end else begin
      valid_637 <= _GEN_4771;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_638 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h27e == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_638 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_638 <= _GEN_4772;
      end
    end else begin
      valid_638 <= _GEN_4772;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_639 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h27f == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_639 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_639 <= _GEN_4773;
      end
    end else begin
      valid_639 <= _GEN_4773;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_640 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h280 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_640 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_640 <= _GEN_4774;
      end
    end else begin
      valid_640 <= _GEN_4774;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_641 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h281 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_641 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_641 <= _GEN_4775;
      end
    end else begin
      valid_641 <= _GEN_4775;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_642 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h282 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_642 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_642 <= _GEN_4776;
      end
    end else begin
      valid_642 <= _GEN_4776;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_643 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h283 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_643 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_643 <= _GEN_4777;
      end
    end else begin
      valid_643 <= _GEN_4777;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_644 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h284 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_644 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_644 <= _GEN_4778;
      end
    end else begin
      valid_644 <= _GEN_4778;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_645 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h285 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_645 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_645 <= _GEN_4779;
      end
    end else begin
      valid_645 <= _GEN_4779;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_646 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h286 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_646 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_646 <= _GEN_4780;
      end
    end else begin
      valid_646 <= _GEN_4780;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_647 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h287 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_647 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_647 <= _GEN_4781;
      end
    end else begin
      valid_647 <= _GEN_4781;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_648 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h288 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_648 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_648 <= _GEN_4782;
      end
    end else begin
      valid_648 <= _GEN_4782;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_649 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h289 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_649 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_649 <= _GEN_4783;
      end
    end else begin
      valid_649 <= _GEN_4783;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_650 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h28a == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_650 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_650 <= _GEN_4784;
      end
    end else begin
      valid_650 <= _GEN_4784;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_651 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h28b == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_651 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_651 <= _GEN_4785;
      end
    end else begin
      valid_651 <= _GEN_4785;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_652 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h28c == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_652 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_652 <= _GEN_4786;
      end
    end else begin
      valid_652 <= _GEN_4786;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_653 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h28d == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_653 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_653 <= _GEN_4787;
      end
    end else begin
      valid_653 <= _GEN_4787;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_654 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h28e == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_654 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_654 <= _GEN_4788;
      end
    end else begin
      valid_654 <= _GEN_4788;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_655 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h28f == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_655 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_655 <= _GEN_4789;
      end
    end else begin
      valid_655 <= _GEN_4789;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_656 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h290 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_656 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_656 <= _GEN_4790;
      end
    end else begin
      valid_656 <= _GEN_4790;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_657 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h291 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_657 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_657 <= _GEN_4791;
      end
    end else begin
      valid_657 <= _GEN_4791;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_658 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h292 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_658 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_658 <= _GEN_4792;
      end
    end else begin
      valid_658 <= _GEN_4792;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_659 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h293 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_659 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_659 <= _GEN_4793;
      end
    end else begin
      valid_659 <= _GEN_4793;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_660 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h294 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_660 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_660 <= _GEN_4794;
      end
    end else begin
      valid_660 <= _GEN_4794;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_661 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h295 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_661 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_661 <= _GEN_4795;
      end
    end else begin
      valid_661 <= _GEN_4795;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_662 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h296 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_662 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_662 <= _GEN_4796;
      end
    end else begin
      valid_662 <= _GEN_4796;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_663 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h297 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_663 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_663 <= _GEN_4797;
      end
    end else begin
      valid_663 <= _GEN_4797;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_664 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h298 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_664 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_664 <= _GEN_4798;
      end
    end else begin
      valid_664 <= _GEN_4798;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_665 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h299 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_665 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_665 <= _GEN_4799;
      end
    end else begin
      valid_665 <= _GEN_4799;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_666 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h29a == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_666 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_666 <= _GEN_4800;
      end
    end else begin
      valid_666 <= _GEN_4800;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_667 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h29b == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_667 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_667 <= _GEN_4801;
      end
    end else begin
      valid_667 <= _GEN_4801;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_668 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h29c == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_668 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_668 <= _GEN_4802;
      end
    end else begin
      valid_668 <= _GEN_4802;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_669 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h29d == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_669 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_669 <= _GEN_4803;
      end
    end else begin
      valid_669 <= _GEN_4803;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_670 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h29e == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_670 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_670 <= _GEN_4804;
      end
    end else begin
      valid_670 <= _GEN_4804;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_671 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h29f == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_671 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_671 <= _GEN_4805;
      end
    end else begin
      valid_671 <= _GEN_4805;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_672 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2a0 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_672 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_672 <= _GEN_4806;
      end
    end else begin
      valid_672 <= _GEN_4806;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_673 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2a1 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_673 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_673 <= _GEN_4807;
      end
    end else begin
      valid_673 <= _GEN_4807;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_674 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2a2 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_674 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_674 <= _GEN_4808;
      end
    end else begin
      valid_674 <= _GEN_4808;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_675 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2a3 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_675 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_675 <= _GEN_4809;
      end
    end else begin
      valid_675 <= _GEN_4809;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_676 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2a4 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_676 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_676 <= _GEN_4810;
      end
    end else begin
      valid_676 <= _GEN_4810;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_677 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2a5 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_677 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_677 <= _GEN_4811;
      end
    end else begin
      valid_677 <= _GEN_4811;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_678 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2a6 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_678 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_678 <= _GEN_4812;
      end
    end else begin
      valid_678 <= _GEN_4812;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_679 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2a7 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_679 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_679 <= _GEN_4813;
      end
    end else begin
      valid_679 <= _GEN_4813;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_680 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2a8 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_680 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_680 <= _GEN_4814;
      end
    end else begin
      valid_680 <= _GEN_4814;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_681 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2a9 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_681 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_681 <= _GEN_4815;
      end
    end else begin
      valid_681 <= _GEN_4815;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_682 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2aa == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_682 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_682 <= _GEN_4816;
      end
    end else begin
      valid_682 <= _GEN_4816;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_683 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2ab == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_683 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_683 <= _GEN_4817;
      end
    end else begin
      valid_683 <= _GEN_4817;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_684 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2ac == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_684 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_684 <= _GEN_4818;
      end
    end else begin
      valid_684 <= _GEN_4818;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_685 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2ad == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_685 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_685 <= _GEN_4819;
      end
    end else begin
      valid_685 <= _GEN_4819;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_686 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2ae == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_686 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_686 <= _GEN_4820;
      end
    end else begin
      valid_686 <= _GEN_4820;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_687 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2af == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_687 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_687 <= _GEN_4821;
      end
    end else begin
      valid_687 <= _GEN_4821;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_688 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2b0 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_688 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_688 <= _GEN_4822;
      end
    end else begin
      valid_688 <= _GEN_4822;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_689 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2b1 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_689 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_689 <= _GEN_4823;
      end
    end else begin
      valid_689 <= _GEN_4823;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_690 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2b2 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_690 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_690 <= _GEN_4824;
      end
    end else begin
      valid_690 <= _GEN_4824;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_691 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2b3 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_691 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_691 <= _GEN_4825;
      end
    end else begin
      valid_691 <= _GEN_4825;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_692 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2b4 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_692 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_692 <= _GEN_4826;
      end
    end else begin
      valid_692 <= _GEN_4826;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_693 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2b5 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_693 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_693 <= _GEN_4827;
      end
    end else begin
      valid_693 <= _GEN_4827;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_694 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2b6 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_694 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_694 <= _GEN_4828;
      end
    end else begin
      valid_694 <= _GEN_4828;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_695 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2b7 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_695 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_695 <= _GEN_4829;
      end
    end else begin
      valid_695 <= _GEN_4829;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_696 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2b8 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_696 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_696 <= _GEN_4830;
      end
    end else begin
      valid_696 <= _GEN_4830;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_697 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2b9 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_697 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_697 <= _GEN_4831;
      end
    end else begin
      valid_697 <= _GEN_4831;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_698 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2ba == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_698 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_698 <= _GEN_4832;
      end
    end else begin
      valid_698 <= _GEN_4832;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_699 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2bb == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_699 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_699 <= _GEN_4833;
      end
    end else begin
      valid_699 <= _GEN_4833;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_700 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2bc == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_700 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_700 <= _GEN_4834;
      end
    end else begin
      valid_700 <= _GEN_4834;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_701 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2bd == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_701 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_701 <= _GEN_4835;
      end
    end else begin
      valid_701 <= _GEN_4835;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_702 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2be == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_702 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_702 <= _GEN_4836;
      end
    end else begin
      valid_702 <= _GEN_4836;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_703 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2bf == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_703 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_703 <= _GEN_4837;
      end
    end else begin
      valid_703 <= _GEN_4837;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_704 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2c0 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_704 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_704 <= _GEN_4838;
      end
    end else begin
      valid_704 <= _GEN_4838;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_705 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2c1 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_705 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_705 <= _GEN_4839;
      end
    end else begin
      valid_705 <= _GEN_4839;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_706 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2c2 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_706 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_706 <= _GEN_4840;
      end
    end else begin
      valid_706 <= _GEN_4840;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_707 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2c3 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_707 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_707 <= _GEN_4841;
      end
    end else begin
      valid_707 <= _GEN_4841;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_708 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2c4 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_708 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_708 <= _GEN_4842;
      end
    end else begin
      valid_708 <= _GEN_4842;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_709 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2c5 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_709 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_709 <= _GEN_4843;
      end
    end else begin
      valid_709 <= _GEN_4843;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_710 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2c6 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_710 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_710 <= _GEN_4844;
      end
    end else begin
      valid_710 <= _GEN_4844;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_711 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2c7 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_711 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_711 <= _GEN_4845;
      end
    end else begin
      valid_711 <= _GEN_4845;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_712 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2c8 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_712 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_712 <= _GEN_4846;
      end
    end else begin
      valid_712 <= _GEN_4846;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_713 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2c9 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_713 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_713 <= _GEN_4847;
      end
    end else begin
      valid_713 <= _GEN_4847;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_714 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2ca == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_714 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_714 <= _GEN_4848;
      end
    end else begin
      valid_714 <= _GEN_4848;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_715 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2cb == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_715 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_715 <= _GEN_4849;
      end
    end else begin
      valid_715 <= _GEN_4849;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_716 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2cc == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_716 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_716 <= _GEN_4850;
      end
    end else begin
      valid_716 <= _GEN_4850;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_717 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2cd == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_717 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_717 <= _GEN_4851;
      end
    end else begin
      valid_717 <= _GEN_4851;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_718 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2ce == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_718 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_718 <= _GEN_4852;
      end
    end else begin
      valid_718 <= _GEN_4852;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_719 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2cf == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_719 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_719 <= _GEN_4853;
      end
    end else begin
      valid_719 <= _GEN_4853;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_720 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2d0 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_720 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_720 <= _GEN_4854;
      end
    end else begin
      valid_720 <= _GEN_4854;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_721 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2d1 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_721 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_721 <= _GEN_4855;
      end
    end else begin
      valid_721 <= _GEN_4855;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_722 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2d2 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_722 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_722 <= _GEN_4856;
      end
    end else begin
      valid_722 <= _GEN_4856;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_723 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2d3 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_723 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_723 <= _GEN_4857;
      end
    end else begin
      valid_723 <= _GEN_4857;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_724 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2d4 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_724 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_724 <= _GEN_4858;
      end
    end else begin
      valid_724 <= _GEN_4858;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_725 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2d5 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_725 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_725 <= _GEN_4859;
      end
    end else begin
      valid_725 <= _GEN_4859;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_726 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2d6 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_726 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_726 <= _GEN_4860;
      end
    end else begin
      valid_726 <= _GEN_4860;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_727 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2d7 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_727 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_727 <= _GEN_4861;
      end
    end else begin
      valid_727 <= _GEN_4861;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_728 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2d8 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_728 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_728 <= _GEN_4862;
      end
    end else begin
      valid_728 <= _GEN_4862;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_729 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2d9 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_729 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_729 <= _GEN_4863;
      end
    end else begin
      valid_729 <= _GEN_4863;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_730 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2da == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_730 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_730 <= _GEN_4864;
      end
    end else begin
      valid_730 <= _GEN_4864;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_731 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2db == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_731 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_731 <= _GEN_4865;
      end
    end else begin
      valid_731 <= _GEN_4865;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_732 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2dc == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_732 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_732 <= _GEN_4866;
      end
    end else begin
      valid_732 <= _GEN_4866;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_733 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2dd == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_733 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_733 <= _GEN_4867;
      end
    end else begin
      valid_733 <= _GEN_4867;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_734 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2de == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_734 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_734 <= _GEN_4868;
      end
    end else begin
      valid_734 <= _GEN_4868;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_735 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2df == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_735 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_735 <= _GEN_4869;
      end
    end else begin
      valid_735 <= _GEN_4869;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_736 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2e0 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_736 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_736 <= _GEN_4870;
      end
    end else begin
      valid_736 <= _GEN_4870;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_737 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2e1 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_737 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_737 <= _GEN_4871;
      end
    end else begin
      valid_737 <= _GEN_4871;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_738 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2e2 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_738 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_738 <= _GEN_4872;
      end
    end else begin
      valid_738 <= _GEN_4872;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_739 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2e3 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_739 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_739 <= _GEN_4873;
      end
    end else begin
      valid_739 <= _GEN_4873;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_740 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2e4 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_740 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_740 <= _GEN_4874;
      end
    end else begin
      valid_740 <= _GEN_4874;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_741 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2e5 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_741 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_741 <= _GEN_4875;
      end
    end else begin
      valid_741 <= _GEN_4875;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_742 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2e6 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_742 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_742 <= _GEN_4876;
      end
    end else begin
      valid_742 <= _GEN_4876;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_743 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2e7 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_743 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_743 <= _GEN_4877;
      end
    end else begin
      valid_743 <= _GEN_4877;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_744 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2e8 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_744 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_744 <= _GEN_4878;
      end
    end else begin
      valid_744 <= _GEN_4878;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_745 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2e9 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_745 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_745 <= _GEN_4879;
      end
    end else begin
      valid_745 <= _GEN_4879;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_746 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2ea == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_746 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_746 <= _GEN_4880;
      end
    end else begin
      valid_746 <= _GEN_4880;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_747 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2eb == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_747 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_747 <= _GEN_4881;
      end
    end else begin
      valid_747 <= _GEN_4881;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_748 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2ec == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_748 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_748 <= _GEN_4882;
      end
    end else begin
      valid_748 <= _GEN_4882;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_749 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2ed == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_749 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_749 <= _GEN_4883;
      end
    end else begin
      valid_749 <= _GEN_4883;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_750 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2ee == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_750 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_750 <= _GEN_4884;
      end
    end else begin
      valid_750 <= _GEN_4884;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_751 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2ef == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_751 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_751 <= _GEN_4885;
      end
    end else begin
      valid_751 <= _GEN_4885;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_752 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2f0 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_752 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_752 <= _GEN_4886;
      end
    end else begin
      valid_752 <= _GEN_4886;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_753 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2f1 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_753 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_753 <= _GEN_4887;
      end
    end else begin
      valid_753 <= _GEN_4887;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_754 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2f2 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_754 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_754 <= _GEN_4888;
      end
    end else begin
      valid_754 <= _GEN_4888;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_755 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2f3 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_755 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_755 <= _GEN_4889;
      end
    end else begin
      valid_755 <= _GEN_4889;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_756 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2f4 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_756 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_756 <= _GEN_4890;
      end
    end else begin
      valid_756 <= _GEN_4890;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_757 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2f5 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_757 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_757 <= _GEN_4891;
      end
    end else begin
      valid_757 <= _GEN_4891;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_758 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2f6 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_758 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_758 <= _GEN_4892;
      end
    end else begin
      valid_758 <= _GEN_4892;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_759 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2f7 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_759 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_759 <= _GEN_4893;
      end
    end else begin
      valid_759 <= _GEN_4893;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_760 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2f8 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_760 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_760 <= _GEN_4894;
      end
    end else begin
      valid_760 <= _GEN_4894;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_761 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2f9 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_761 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_761 <= _GEN_4895;
      end
    end else begin
      valid_761 <= _GEN_4895;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_762 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2fa == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_762 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_762 <= _GEN_4896;
      end
    end else begin
      valid_762 <= _GEN_4896;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_763 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2fb == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_763 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_763 <= _GEN_4897;
      end
    end else begin
      valid_763 <= _GEN_4897;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_764 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2fc == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_764 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_764 <= _GEN_4898;
      end
    end else begin
      valid_764 <= _GEN_4898;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_765 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2fd == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_765 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_765 <= _GEN_4899;
      end
    end else begin
      valid_765 <= _GEN_4899;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_766 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2fe == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_766 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_766 <= _GEN_4900;
      end
    end else begin
      valid_766 <= _GEN_4900;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_767 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h2ff == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_767 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_767 <= _GEN_4901;
      end
    end else begin
      valid_767 <= _GEN_4901;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_768 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h300 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_768 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_768 <= _GEN_4902;
      end
    end else begin
      valid_768 <= _GEN_4902;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_769 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h301 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_769 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_769 <= _GEN_4903;
      end
    end else begin
      valid_769 <= _GEN_4903;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_770 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h302 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_770 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_770 <= _GEN_4904;
      end
    end else begin
      valid_770 <= _GEN_4904;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_771 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h303 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_771 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_771 <= _GEN_4905;
      end
    end else begin
      valid_771 <= _GEN_4905;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_772 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h304 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_772 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_772 <= _GEN_4906;
      end
    end else begin
      valid_772 <= _GEN_4906;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_773 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h305 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_773 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_773 <= _GEN_4907;
      end
    end else begin
      valid_773 <= _GEN_4907;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_774 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h306 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_774 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_774 <= _GEN_4908;
      end
    end else begin
      valid_774 <= _GEN_4908;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_775 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h307 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_775 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_775 <= _GEN_4909;
      end
    end else begin
      valid_775 <= _GEN_4909;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_776 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h308 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_776 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_776 <= _GEN_4910;
      end
    end else begin
      valid_776 <= _GEN_4910;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_777 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h309 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_777 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_777 <= _GEN_4911;
      end
    end else begin
      valid_777 <= _GEN_4911;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_778 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h30a == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_778 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_778 <= _GEN_4912;
      end
    end else begin
      valid_778 <= _GEN_4912;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_779 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h30b == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_779 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_779 <= _GEN_4913;
      end
    end else begin
      valid_779 <= _GEN_4913;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_780 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h30c == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_780 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_780 <= _GEN_4914;
      end
    end else begin
      valid_780 <= _GEN_4914;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_781 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h30d == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_781 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_781 <= _GEN_4915;
      end
    end else begin
      valid_781 <= _GEN_4915;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_782 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h30e == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_782 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_782 <= _GEN_4916;
      end
    end else begin
      valid_782 <= _GEN_4916;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_783 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h30f == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_783 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_783 <= _GEN_4917;
      end
    end else begin
      valid_783 <= _GEN_4917;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_784 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h310 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_784 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_784 <= _GEN_4918;
      end
    end else begin
      valid_784 <= _GEN_4918;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_785 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h311 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_785 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_785 <= _GEN_4919;
      end
    end else begin
      valid_785 <= _GEN_4919;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_786 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h312 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_786 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_786 <= _GEN_4920;
      end
    end else begin
      valid_786 <= _GEN_4920;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_787 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h313 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_787 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_787 <= _GEN_4921;
      end
    end else begin
      valid_787 <= _GEN_4921;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_788 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h314 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_788 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_788 <= _GEN_4922;
      end
    end else begin
      valid_788 <= _GEN_4922;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_789 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h315 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_789 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_789 <= _GEN_4923;
      end
    end else begin
      valid_789 <= _GEN_4923;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_790 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h316 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_790 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_790 <= _GEN_4924;
      end
    end else begin
      valid_790 <= _GEN_4924;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_791 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h317 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_791 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_791 <= _GEN_4925;
      end
    end else begin
      valid_791 <= _GEN_4925;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_792 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h318 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_792 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_792 <= _GEN_4926;
      end
    end else begin
      valid_792 <= _GEN_4926;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_793 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h319 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_793 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_793 <= _GEN_4927;
      end
    end else begin
      valid_793 <= _GEN_4927;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_794 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h31a == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_794 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_794 <= _GEN_4928;
      end
    end else begin
      valid_794 <= _GEN_4928;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_795 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h31b == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_795 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_795 <= _GEN_4929;
      end
    end else begin
      valid_795 <= _GEN_4929;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_796 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h31c == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_796 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_796 <= _GEN_4930;
      end
    end else begin
      valid_796 <= _GEN_4930;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_797 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h31d == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_797 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_797 <= _GEN_4931;
      end
    end else begin
      valid_797 <= _GEN_4931;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_798 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h31e == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_798 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_798 <= _GEN_4932;
      end
    end else begin
      valid_798 <= _GEN_4932;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_799 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h31f == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_799 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_799 <= _GEN_4933;
      end
    end else begin
      valid_799 <= _GEN_4933;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_800 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h320 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_800 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_800 <= _GEN_4934;
      end
    end else begin
      valid_800 <= _GEN_4934;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_801 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h321 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_801 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_801 <= _GEN_4935;
      end
    end else begin
      valid_801 <= _GEN_4935;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_802 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h322 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_802 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_802 <= _GEN_4936;
      end
    end else begin
      valid_802 <= _GEN_4936;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_803 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h323 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_803 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_803 <= _GEN_4937;
      end
    end else begin
      valid_803 <= _GEN_4937;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_804 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h324 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_804 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_804 <= _GEN_4938;
      end
    end else begin
      valid_804 <= _GEN_4938;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_805 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h325 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_805 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_805 <= _GEN_4939;
      end
    end else begin
      valid_805 <= _GEN_4939;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_806 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h326 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_806 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_806 <= _GEN_4940;
      end
    end else begin
      valid_806 <= _GEN_4940;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_807 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h327 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_807 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_807 <= _GEN_4941;
      end
    end else begin
      valid_807 <= _GEN_4941;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_808 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h328 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_808 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_808 <= _GEN_4942;
      end
    end else begin
      valid_808 <= _GEN_4942;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_809 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h329 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_809 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_809 <= _GEN_4943;
      end
    end else begin
      valid_809 <= _GEN_4943;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_810 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h32a == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_810 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_810 <= _GEN_4944;
      end
    end else begin
      valid_810 <= _GEN_4944;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_811 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h32b == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_811 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_811 <= _GEN_4945;
      end
    end else begin
      valid_811 <= _GEN_4945;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_812 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h32c == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_812 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_812 <= _GEN_4946;
      end
    end else begin
      valid_812 <= _GEN_4946;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_813 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h32d == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_813 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_813 <= _GEN_4947;
      end
    end else begin
      valid_813 <= _GEN_4947;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_814 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h32e == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_814 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_814 <= _GEN_4948;
      end
    end else begin
      valid_814 <= _GEN_4948;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_815 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h32f == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_815 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_815 <= _GEN_4949;
      end
    end else begin
      valid_815 <= _GEN_4949;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_816 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h330 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_816 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_816 <= _GEN_4950;
      end
    end else begin
      valid_816 <= _GEN_4950;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_817 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h331 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_817 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_817 <= _GEN_4951;
      end
    end else begin
      valid_817 <= _GEN_4951;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_818 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h332 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_818 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_818 <= _GEN_4952;
      end
    end else begin
      valid_818 <= _GEN_4952;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_819 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h333 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_819 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_819 <= _GEN_4953;
      end
    end else begin
      valid_819 <= _GEN_4953;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_820 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h334 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_820 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_820 <= _GEN_4954;
      end
    end else begin
      valid_820 <= _GEN_4954;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_821 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h335 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_821 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_821 <= _GEN_4955;
      end
    end else begin
      valid_821 <= _GEN_4955;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_822 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h336 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_822 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_822 <= _GEN_4956;
      end
    end else begin
      valid_822 <= _GEN_4956;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_823 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h337 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_823 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_823 <= _GEN_4957;
      end
    end else begin
      valid_823 <= _GEN_4957;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_824 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h338 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_824 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_824 <= _GEN_4958;
      end
    end else begin
      valid_824 <= _GEN_4958;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_825 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h339 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_825 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_825 <= _GEN_4959;
      end
    end else begin
      valid_825 <= _GEN_4959;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_826 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h33a == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_826 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_826 <= _GEN_4960;
      end
    end else begin
      valid_826 <= _GEN_4960;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_827 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h33b == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_827 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_827 <= _GEN_4961;
      end
    end else begin
      valid_827 <= _GEN_4961;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_828 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h33c == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_828 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_828 <= _GEN_4962;
      end
    end else begin
      valid_828 <= _GEN_4962;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_829 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h33d == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_829 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_829 <= _GEN_4963;
      end
    end else begin
      valid_829 <= _GEN_4963;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_830 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h33e == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_830 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_830 <= _GEN_4964;
      end
    end else begin
      valid_830 <= _GEN_4964;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_831 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h33f == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_831 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_831 <= _GEN_4965;
      end
    end else begin
      valid_831 <= _GEN_4965;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_832 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h340 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_832 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_832 <= _GEN_4966;
      end
    end else begin
      valid_832 <= _GEN_4966;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_833 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h341 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_833 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_833 <= _GEN_4967;
      end
    end else begin
      valid_833 <= _GEN_4967;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_834 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h342 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_834 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_834 <= _GEN_4968;
      end
    end else begin
      valid_834 <= _GEN_4968;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_835 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h343 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_835 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_835 <= _GEN_4969;
      end
    end else begin
      valid_835 <= _GEN_4969;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_836 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h344 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_836 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_836 <= _GEN_4970;
      end
    end else begin
      valid_836 <= _GEN_4970;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_837 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h345 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_837 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_837 <= _GEN_4971;
      end
    end else begin
      valid_837 <= _GEN_4971;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_838 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h346 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_838 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_838 <= _GEN_4972;
      end
    end else begin
      valid_838 <= _GEN_4972;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_839 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h347 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_839 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_839 <= _GEN_4973;
      end
    end else begin
      valid_839 <= _GEN_4973;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_840 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h348 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_840 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_840 <= _GEN_4974;
      end
    end else begin
      valid_840 <= _GEN_4974;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_841 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h349 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_841 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_841 <= _GEN_4975;
      end
    end else begin
      valid_841 <= _GEN_4975;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_842 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h34a == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_842 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_842 <= _GEN_4976;
      end
    end else begin
      valid_842 <= _GEN_4976;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_843 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h34b == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_843 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_843 <= _GEN_4977;
      end
    end else begin
      valid_843 <= _GEN_4977;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_844 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h34c == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_844 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_844 <= _GEN_4978;
      end
    end else begin
      valid_844 <= _GEN_4978;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_845 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h34d == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_845 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_845 <= _GEN_4979;
      end
    end else begin
      valid_845 <= _GEN_4979;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_846 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h34e == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_846 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_846 <= _GEN_4980;
      end
    end else begin
      valid_846 <= _GEN_4980;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_847 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h34f == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_847 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_847 <= _GEN_4981;
      end
    end else begin
      valid_847 <= _GEN_4981;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_848 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h350 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_848 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_848 <= _GEN_4982;
      end
    end else begin
      valid_848 <= _GEN_4982;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_849 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h351 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_849 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_849 <= _GEN_4983;
      end
    end else begin
      valid_849 <= _GEN_4983;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_850 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h352 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_850 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_850 <= _GEN_4984;
      end
    end else begin
      valid_850 <= _GEN_4984;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_851 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h353 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_851 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_851 <= _GEN_4985;
      end
    end else begin
      valid_851 <= _GEN_4985;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_852 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h354 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_852 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_852 <= _GEN_4986;
      end
    end else begin
      valid_852 <= _GEN_4986;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_853 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h355 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_853 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_853 <= _GEN_4987;
      end
    end else begin
      valid_853 <= _GEN_4987;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_854 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h356 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_854 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_854 <= _GEN_4988;
      end
    end else begin
      valid_854 <= _GEN_4988;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_855 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h357 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_855 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_855 <= _GEN_4989;
      end
    end else begin
      valid_855 <= _GEN_4989;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_856 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h358 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_856 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_856 <= _GEN_4990;
      end
    end else begin
      valid_856 <= _GEN_4990;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_857 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h359 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_857 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_857 <= _GEN_4991;
      end
    end else begin
      valid_857 <= _GEN_4991;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_858 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h35a == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_858 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_858 <= _GEN_4992;
      end
    end else begin
      valid_858 <= _GEN_4992;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_859 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h35b == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_859 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_859 <= _GEN_4993;
      end
    end else begin
      valid_859 <= _GEN_4993;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_860 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h35c == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_860 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_860 <= _GEN_4994;
      end
    end else begin
      valid_860 <= _GEN_4994;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_861 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h35d == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_861 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_861 <= _GEN_4995;
      end
    end else begin
      valid_861 <= _GEN_4995;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_862 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h35e == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_862 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_862 <= _GEN_4996;
      end
    end else begin
      valid_862 <= _GEN_4996;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_863 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h35f == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_863 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_863 <= _GEN_4997;
      end
    end else begin
      valid_863 <= _GEN_4997;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_864 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h360 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_864 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_864 <= _GEN_4998;
      end
    end else begin
      valid_864 <= _GEN_4998;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_865 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h361 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_865 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_865 <= _GEN_4999;
      end
    end else begin
      valid_865 <= _GEN_4999;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_866 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h362 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_866 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_866 <= _GEN_5000;
      end
    end else begin
      valid_866 <= _GEN_5000;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_867 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h363 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_867 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_867 <= _GEN_5001;
      end
    end else begin
      valid_867 <= _GEN_5001;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_868 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h364 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_868 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_868 <= _GEN_5002;
      end
    end else begin
      valid_868 <= _GEN_5002;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_869 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h365 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_869 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_869 <= _GEN_5003;
      end
    end else begin
      valid_869 <= _GEN_5003;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_870 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h366 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_870 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_870 <= _GEN_5004;
      end
    end else begin
      valid_870 <= _GEN_5004;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_871 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h367 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_871 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_871 <= _GEN_5005;
      end
    end else begin
      valid_871 <= _GEN_5005;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_872 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h368 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_872 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_872 <= _GEN_5006;
      end
    end else begin
      valid_872 <= _GEN_5006;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_873 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h369 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_873 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_873 <= _GEN_5007;
      end
    end else begin
      valid_873 <= _GEN_5007;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_874 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h36a == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_874 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_874 <= _GEN_5008;
      end
    end else begin
      valid_874 <= _GEN_5008;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_875 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h36b == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_875 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_875 <= _GEN_5009;
      end
    end else begin
      valid_875 <= _GEN_5009;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_876 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h36c == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_876 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_876 <= _GEN_5010;
      end
    end else begin
      valid_876 <= _GEN_5010;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_877 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h36d == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_877 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_877 <= _GEN_5011;
      end
    end else begin
      valid_877 <= _GEN_5011;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_878 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h36e == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_878 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_878 <= _GEN_5012;
      end
    end else begin
      valid_878 <= _GEN_5012;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_879 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h36f == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_879 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_879 <= _GEN_5013;
      end
    end else begin
      valid_879 <= _GEN_5013;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_880 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h370 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_880 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_880 <= _GEN_5014;
      end
    end else begin
      valid_880 <= _GEN_5014;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_881 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h371 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_881 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_881 <= _GEN_5015;
      end
    end else begin
      valid_881 <= _GEN_5015;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_882 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h372 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_882 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_882 <= _GEN_5016;
      end
    end else begin
      valid_882 <= _GEN_5016;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_883 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h373 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_883 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_883 <= _GEN_5017;
      end
    end else begin
      valid_883 <= _GEN_5017;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_884 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h374 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_884 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_884 <= _GEN_5018;
      end
    end else begin
      valid_884 <= _GEN_5018;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_885 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h375 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_885 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_885 <= _GEN_5019;
      end
    end else begin
      valid_885 <= _GEN_5019;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_886 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h376 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_886 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_886 <= _GEN_5020;
      end
    end else begin
      valid_886 <= _GEN_5020;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_887 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h377 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_887 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_887 <= _GEN_5021;
      end
    end else begin
      valid_887 <= _GEN_5021;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_888 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h378 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_888 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_888 <= _GEN_5022;
      end
    end else begin
      valid_888 <= _GEN_5022;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_889 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h379 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_889 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_889 <= _GEN_5023;
      end
    end else begin
      valid_889 <= _GEN_5023;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_890 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h37a == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_890 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_890 <= _GEN_5024;
      end
    end else begin
      valid_890 <= _GEN_5024;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_891 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h37b == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_891 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_891 <= _GEN_5025;
      end
    end else begin
      valid_891 <= _GEN_5025;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_892 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h37c == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_892 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_892 <= _GEN_5026;
      end
    end else begin
      valid_892 <= _GEN_5026;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_893 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h37d == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_893 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_893 <= _GEN_5027;
      end
    end else begin
      valid_893 <= _GEN_5027;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_894 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h37e == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_894 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_894 <= _GEN_5028;
      end
    end else begin
      valid_894 <= _GEN_5028;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_895 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h37f == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_895 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_895 <= _GEN_5029;
      end
    end else begin
      valid_895 <= _GEN_5029;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_896 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h380 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_896 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_896 <= _GEN_5030;
      end
    end else begin
      valid_896 <= _GEN_5030;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_897 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h381 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_897 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_897 <= _GEN_5031;
      end
    end else begin
      valid_897 <= _GEN_5031;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_898 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h382 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_898 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_898 <= _GEN_5032;
      end
    end else begin
      valid_898 <= _GEN_5032;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_899 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h383 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_899 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_899 <= _GEN_5033;
      end
    end else begin
      valid_899 <= _GEN_5033;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_900 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h384 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_900 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_900 <= _GEN_5034;
      end
    end else begin
      valid_900 <= _GEN_5034;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_901 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h385 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_901 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_901 <= _GEN_5035;
      end
    end else begin
      valid_901 <= _GEN_5035;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_902 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h386 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_902 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_902 <= _GEN_5036;
      end
    end else begin
      valid_902 <= _GEN_5036;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_903 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h387 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_903 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_903 <= _GEN_5037;
      end
    end else begin
      valid_903 <= _GEN_5037;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_904 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h388 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_904 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_904 <= _GEN_5038;
      end
    end else begin
      valid_904 <= _GEN_5038;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_905 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h389 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_905 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_905 <= _GEN_5039;
      end
    end else begin
      valid_905 <= _GEN_5039;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_906 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h38a == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_906 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_906 <= _GEN_5040;
      end
    end else begin
      valid_906 <= _GEN_5040;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_907 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h38b == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_907 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_907 <= _GEN_5041;
      end
    end else begin
      valid_907 <= _GEN_5041;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_908 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h38c == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_908 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_908 <= _GEN_5042;
      end
    end else begin
      valid_908 <= _GEN_5042;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_909 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h38d == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_909 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_909 <= _GEN_5043;
      end
    end else begin
      valid_909 <= _GEN_5043;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_910 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h38e == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_910 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_910 <= _GEN_5044;
      end
    end else begin
      valid_910 <= _GEN_5044;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_911 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h38f == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_911 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_911 <= _GEN_5045;
      end
    end else begin
      valid_911 <= _GEN_5045;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_912 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h390 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_912 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_912 <= _GEN_5046;
      end
    end else begin
      valid_912 <= _GEN_5046;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_913 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h391 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_913 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_913 <= _GEN_5047;
      end
    end else begin
      valid_913 <= _GEN_5047;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_914 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h392 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_914 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_914 <= _GEN_5048;
      end
    end else begin
      valid_914 <= _GEN_5048;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_915 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h393 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_915 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_915 <= _GEN_5049;
      end
    end else begin
      valid_915 <= _GEN_5049;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_916 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h394 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_916 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_916 <= _GEN_5050;
      end
    end else begin
      valid_916 <= _GEN_5050;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_917 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h395 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_917 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_917 <= _GEN_5051;
      end
    end else begin
      valid_917 <= _GEN_5051;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_918 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h396 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_918 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_918 <= _GEN_5052;
      end
    end else begin
      valid_918 <= _GEN_5052;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_919 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h397 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_919 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_919 <= _GEN_5053;
      end
    end else begin
      valid_919 <= _GEN_5053;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_920 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h398 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_920 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_920 <= _GEN_5054;
      end
    end else begin
      valid_920 <= _GEN_5054;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_921 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h399 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_921 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_921 <= _GEN_5055;
      end
    end else begin
      valid_921 <= _GEN_5055;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_922 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h39a == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_922 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_922 <= _GEN_5056;
      end
    end else begin
      valid_922 <= _GEN_5056;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_923 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h39b == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_923 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_923 <= _GEN_5057;
      end
    end else begin
      valid_923 <= _GEN_5057;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_924 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h39c == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_924 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_924 <= _GEN_5058;
      end
    end else begin
      valid_924 <= _GEN_5058;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_925 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h39d == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_925 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_925 <= _GEN_5059;
      end
    end else begin
      valid_925 <= _GEN_5059;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_926 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h39e == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_926 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_926 <= _GEN_5060;
      end
    end else begin
      valid_926 <= _GEN_5060;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_927 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h39f == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_927 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_927 <= _GEN_5061;
      end
    end else begin
      valid_927 <= _GEN_5061;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_928 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3a0 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_928 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_928 <= _GEN_5062;
      end
    end else begin
      valid_928 <= _GEN_5062;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_929 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3a1 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_929 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_929 <= _GEN_5063;
      end
    end else begin
      valid_929 <= _GEN_5063;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_930 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3a2 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_930 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_930 <= _GEN_5064;
      end
    end else begin
      valid_930 <= _GEN_5064;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_931 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3a3 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_931 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_931 <= _GEN_5065;
      end
    end else begin
      valid_931 <= _GEN_5065;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_932 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3a4 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_932 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_932 <= _GEN_5066;
      end
    end else begin
      valid_932 <= _GEN_5066;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_933 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3a5 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_933 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_933 <= _GEN_5067;
      end
    end else begin
      valid_933 <= _GEN_5067;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_934 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3a6 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_934 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_934 <= _GEN_5068;
      end
    end else begin
      valid_934 <= _GEN_5068;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_935 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3a7 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_935 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_935 <= _GEN_5069;
      end
    end else begin
      valid_935 <= _GEN_5069;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_936 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3a8 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_936 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_936 <= _GEN_5070;
      end
    end else begin
      valid_936 <= _GEN_5070;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_937 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3a9 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_937 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_937 <= _GEN_5071;
      end
    end else begin
      valid_937 <= _GEN_5071;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_938 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3aa == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_938 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_938 <= _GEN_5072;
      end
    end else begin
      valid_938 <= _GEN_5072;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_939 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3ab == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_939 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_939 <= _GEN_5073;
      end
    end else begin
      valid_939 <= _GEN_5073;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_940 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3ac == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_940 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_940 <= _GEN_5074;
      end
    end else begin
      valid_940 <= _GEN_5074;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_941 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3ad == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_941 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_941 <= _GEN_5075;
      end
    end else begin
      valid_941 <= _GEN_5075;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_942 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3ae == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_942 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_942 <= _GEN_5076;
      end
    end else begin
      valid_942 <= _GEN_5076;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_943 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3af == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_943 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_943 <= _GEN_5077;
      end
    end else begin
      valid_943 <= _GEN_5077;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_944 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3b0 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_944 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_944 <= _GEN_5078;
      end
    end else begin
      valid_944 <= _GEN_5078;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_945 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3b1 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_945 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_945 <= _GEN_5079;
      end
    end else begin
      valid_945 <= _GEN_5079;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_946 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3b2 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_946 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_946 <= _GEN_5080;
      end
    end else begin
      valid_946 <= _GEN_5080;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_947 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3b3 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_947 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_947 <= _GEN_5081;
      end
    end else begin
      valid_947 <= _GEN_5081;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_948 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3b4 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_948 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_948 <= _GEN_5082;
      end
    end else begin
      valid_948 <= _GEN_5082;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_949 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3b5 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_949 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_949 <= _GEN_5083;
      end
    end else begin
      valid_949 <= _GEN_5083;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_950 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3b6 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_950 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_950 <= _GEN_5084;
      end
    end else begin
      valid_950 <= _GEN_5084;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_951 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3b7 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_951 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_951 <= _GEN_5085;
      end
    end else begin
      valid_951 <= _GEN_5085;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_952 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3b8 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_952 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_952 <= _GEN_5086;
      end
    end else begin
      valid_952 <= _GEN_5086;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_953 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3b9 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_953 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_953 <= _GEN_5087;
      end
    end else begin
      valid_953 <= _GEN_5087;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_954 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3ba == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_954 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_954 <= _GEN_5088;
      end
    end else begin
      valid_954 <= _GEN_5088;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_955 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3bb == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_955 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_955 <= _GEN_5089;
      end
    end else begin
      valid_955 <= _GEN_5089;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_956 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3bc == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_956 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_956 <= _GEN_5090;
      end
    end else begin
      valid_956 <= _GEN_5090;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_957 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3bd == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_957 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_957 <= _GEN_5091;
      end
    end else begin
      valid_957 <= _GEN_5091;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_958 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3be == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_958 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_958 <= _GEN_5092;
      end
    end else begin
      valid_958 <= _GEN_5092;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_959 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3bf == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_959 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_959 <= _GEN_5093;
      end
    end else begin
      valid_959 <= _GEN_5093;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_960 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3c0 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_960 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_960 <= _GEN_5094;
      end
    end else begin
      valid_960 <= _GEN_5094;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_961 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3c1 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_961 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_961 <= _GEN_5095;
      end
    end else begin
      valid_961 <= _GEN_5095;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_962 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3c2 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_962 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_962 <= _GEN_5096;
      end
    end else begin
      valid_962 <= _GEN_5096;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_963 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3c3 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_963 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_963 <= _GEN_5097;
      end
    end else begin
      valid_963 <= _GEN_5097;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_964 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3c4 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_964 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_964 <= _GEN_5098;
      end
    end else begin
      valid_964 <= _GEN_5098;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_965 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3c5 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_965 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_965 <= _GEN_5099;
      end
    end else begin
      valid_965 <= _GEN_5099;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_966 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3c6 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_966 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_966 <= _GEN_5100;
      end
    end else begin
      valid_966 <= _GEN_5100;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_967 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3c7 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_967 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_967 <= _GEN_5101;
      end
    end else begin
      valid_967 <= _GEN_5101;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_968 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3c8 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_968 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_968 <= _GEN_5102;
      end
    end else begin
      valid_968 <= _GEN_5102;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_969 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3c9 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_969 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_969 <= _GEN_5103;
      end
    end else begin
      valid_969 <= _GEN_5103;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_970 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3ca == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_970 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_970 <= _GEN_5104;
      end
    end else begin
      valid_970 <= _GEN_5104;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_971 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3cb == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_971 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_971 <= _GEN_5105;
      end
    end else begin
      valid_971 <= _GEN_5105;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_972 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3cc == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_972 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_972 <= _GEN_5106;
      end
    end else begin
      valid_972 <= _GEN_5106;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_973 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3cd == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_973 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_973 <= _GEN_5107;
      end
    end else begin
      valid_973 <= _GEN_5107;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_974 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3ce == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_974 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_974 <= _GEN_5108;
      end
    end else begin
      valid_974 <= _GEN_5108;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_975 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3cf == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_975 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_975 <= _GEN_5109;
      end
    end else begin
      valid_975 <= _GEN_5109;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_976 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3d0 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_976 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_976 <= _GEN_5110;
      end
    end else begin
      valid_976 <= _GEN_5110;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_977 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3d1 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_977 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_977 <= _GEN_5111;
      end
    end else begin
      valid_977 <= _GEN_5111;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_978 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3d2 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_978 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_978 <= _GEN_5112;
      end
    end else begin
      valid_978 <= _GEN_5112;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_979 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3d3 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_979 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_979 <= _GEN_5113;
      end
    end else begin
      valid_979 <= _GEN_5113;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_980 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3d4 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_980 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_980 <= _GEN_5114;
      end
    end else begin
      valid_980 <= _GEN_5114;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_981 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3d5 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_981 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_981 <= _GEN_5115;
      end
    end else begin
      valid_981 <= _GEN_5115;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_982 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3d6 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_982 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_982 <= _GEN_5116;
      end
    end else begin
      valid_982 <= _GEN_5116;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_983 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3d7 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_983 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_983 <= _GEN_5117;
      end
    end else begin
      valid_983 <= _GEN_5117;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_984 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3d8 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_984 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_984 <= _GEN_5118;
      end
    end else begin
      valid_984 <= _GEN_5118;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_985 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3d9 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_985 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_985 <= _GEN_5119;
      end
    end else begin
      valid_985 <= _GEN_5119;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_986 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3da == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_986 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_986 <= _GEN_5120;
      end
    end else begin
      valid_986 <= _GEN_5120;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_987 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3db == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_987 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_987 <= _GEN_5121;
      end
    end else begin
      valid_987 <= _GEN_5121;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_988 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3dc == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_988 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_988 <= _GEN_5122;
      end
    end else begin
      valid_988 <= _GEN_5122;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_989 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3dd == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_989 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_989 <= _GEN_5123;
      end
    end else begin
      valid_989 <= _GEN_5123;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_990 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3de == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_990 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_990 <= _GEN_5124;
      end
    end else begin
      valid_990 <= _GEN_5124;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_991 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3df == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_991 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_991 <= _GEN_5125;
      end
    end else begin
      valid_991 <= _GEN_5125;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_992 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3e0 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_992 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_992 <= _GEN_5126;
      end
    end else begin
      valid_992 <= _GEN_5126;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_993 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3e1 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_993 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_993 <= _GEN_5127;
      end
    end else begin
      valid_993 <= _GEN_5127;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_994 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3e2 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_994 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_994 <= _GEN_5128;
      end
    end else begin
      valid_994 <= _GEN_5128;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_995 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3e3 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_995 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_995 <= _GEN_5129;
      end
    end else begin
      valid_995 <= _GEN_5129;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_996 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3e4 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_996 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_996 <= _GEN_5130;
      end
    end else begin
      valid_996 <= _GEN_5130;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_997 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3e5 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_997 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_997 <= _GEN_5131;
      end
    end else begin
      valid_997 <= _GEN_5131;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_998 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3e6 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_998 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_998 <= _GEN_5132;
      end
    end else begin
      valid_998 <= _GEN_5132;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_999 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3e7 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_999 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_999 <= _GEN_5133;
      end
    end else begin
      valid_999 <= _GEN_5133;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_1000 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3e8 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_1000 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_1000 <= _GEN_5134;
      end
    end else begin
      valid_1000 <= _GEN_5134;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_1001 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3e9 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_1001 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_1001 <= _GEN_5135;
      end
    end else begin
      valid_1001 <= _GEN_5135;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_1002 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3ea == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_1002 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_1002 <= _GEN_5136;
      end
    end else begin
      valid_1002 <= _GEN_5136;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_1003 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3eb == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_1003 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_1003 <= _GEN_5137;
      end
    end else begin
      valid_1003 <= _GEN_5137;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_1004 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3ec == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_1004 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_1004 <= _GEN_5138;
      end
    end else begin
      valid_1004 <= _GEN_5138;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_1005 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3ed == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_1005 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_1005 <= _GEN_5139;
      end
    end else begin
      valid_1005 <= _GEN_5139;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_1006 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3ee == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_1006 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_1006 <= _GEN_5140;
      end
    end else begin
      valid_1006 <= _GEN_5140;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_1007 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3ef == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_1007 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_1007 <= _GEN_5141;
      end
    end else begin
      valid_1007 <= _GEN_5141;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_1008 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3f0 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_1008 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_1008 <= _GEN_5142;
      end
    end else begin
      valid_1008 <= _GEN_5142;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_1009 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3f1 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_1009 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_1009 <= _GEN_5143;
      end
    end else begin
      valid_1009 <= _GEN_5143;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_1010 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3f2 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_1010 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_1010 <= _GEN_5144;
      end
    end else begin
      valid_1010 <= _GEN_5144;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_1011 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3f3 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_1011 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_1011 <= _GEN_5145;
      end
    end else begin
      valid_1011 <= _GEN_5145;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_1012 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3f4 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_1012 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_1012 <= _GEN_5146;
      end
    end else begin
      valid_1012 <= _GEN_5146;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_1013 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3f5 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_1013 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_1013 <= _GEN_5147;
      end
    end else begin
      valid_1013 <= _GEN_5147;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_1014 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3f6 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_1014 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_1014 <= _GEN_5148;
      end
    end else begin
      valid_1014 <= _GEN_5148;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_1015 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3f7 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_1015 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_1015 <= _GEN_5149;
      end
    end else begin
      valid_1015 <= _GEN_5149;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_1016 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3f8 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_1016 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_1016 <= _GEN_5150;
      end
    end else begin
      valid_1016 <= _GEN_5150;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_1017 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3f9 == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_1017 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_1017 <= _GEN_5151;
      end
    end else begin
      valid_1017 <= _GEN_5151;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_1018 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3fa == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_1018 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_1018 <= _GEN_5152;
      end
    end else begin
      valid_1018 <= _GEN_5152;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_1019 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3fb == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_1019 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_1019 <= _GEN_5153;
      end
    end else begin
      valid_1019 <= _GEN_5153;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_1020 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3fc == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_1020 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_1020 <= _GEN_5154;
      end
    end else begin
      valid_1020 <= _GEN_5154;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_1021 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3fd == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_1021 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_1021 <= _GEN_5155;
      end
    end else begin
      valid_1021 <= _GEN_5155;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_1022 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3fe == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_1022 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_1022 <= _GEN_5156;
      end
    end else begin
      valid_1022 <= _GEN_5156;
    end
    if (reset) begin // @[DCache.scala 56:22]
      valid_1023 <= 1'h0; // @[DCache.scala 56:22]
    end else if (probing & _probing_T_1 & probe_hit) begin // @[DCache.scala 240:43]
      if (10'h3ff == _GEN_4[14:5]) begin // @[DCache.scala 241:33]
        valid_1023 <= 1'h0; // @[DCache.scala 241:33]
      end else begin
        valid_1023 <= _GEN_5157;
      end
    end else begin
      valid_1023 <= _GEN_5157;
    end
    array_out_REG <= io_cache_req_ready & io_cache_req_valid; // @[Decoupled.scala 51:35]
    if (reset) begin // @[Reg.scala 35:20]
      array_out_r <= 273'h0; // @[Reg.scala 35:20]
    end else if (array_out_REG) begin // @[Utils.scala 50:8]
      array_out_r <= array_io_rdata;
    end
    if (reset) begin // @[DCache.scala 128:30]
      lrsc_addr <= 27'h0; // @[DCache.scala 128:30]
    end else if (_array_io_en_T_1 & is_lr_r) begin // @[DCache.scala 132:30]
      lrsc_addr <= req_r_addr[31:5]; // @[DCache.scala 134:19]
    end
    if (reset) begin // @[Reg.scala 35:20]
      sc_fail_r <= 1'h0; // @[Reg.scala 35:20]
    end else if (_req_r_T) begin // @[Reg.scala 36:18]
      sc_fail_r <= sc_fail; // @[Reg.scala 36:22]
    end
    probe_out_REG <= tl_b_ready & auto_out_b_valid; // @[Decoupled.scala 51:35]
    if (reset) begin // @[Reg.scala 35:20]
      probe_out_r <= 273'h0; // @[Reg.scala 35:20]
    end else if (probe_out_REG) begin // @[Reg.scala 36:18]
      probe_out_r <= array_io_rdata; // @[Reg.scala 36:22]
    end
    release_addr_aligned_REG <= array_io_addr; // @[DCache.scala 245:56]
    if (reset) begin // @[Counter.scala 61:40]
      source <= 2'h0; // @[Counter.scala 61:40]
    end else if (_source_T_2) begin // @[Counter.scala 118:16]
      source <= _source_wrap_value_T_1; // @[Counter.scala 77:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  probing = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  lrsc_reserved = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  lrsc_counter = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  tl_b_bits_r_size = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  tl_b_bits_r_source = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  tl_b_bits_r_address = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  state = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  tl_d_bits_r_sink = _RAND_7[5:0];
  _RAND_8 = {8{`RANDOM}};
  tl_d_bits_r_data = _RAND_8[255:0];
  _RAND_9 = {2{`RANDOM}};
  req_r_addr = _RAND_9[38:0];
  _RAND_10 = {2{`RANDOM}};
  req_r_wdata = _RAND_10[63:0];
  _RAND_11 = {1{`RANDOM}};
  req_r_wmask = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  req_r_wen = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  req_r_len = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  req_r_lrsc = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  req_r_amo = _RAND_15[4:0];
  _RAND_16 = {1{`RANDOM}};
  valid_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  valid_1 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  valid_2 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  valid_3 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  valid_4 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  valid_5 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  valid_6 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  valid_7 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  valid_8 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  valid_9 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  valid_10 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  valid_11 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  valid_12 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  valid_13 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  valid_14 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  valid_15 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  valid_16 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  valid_17 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  valid_18 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  valid_19 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  valid_20 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  valid_21 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  valid_22 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  valid_23 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  valid_24 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  valid_25 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  valid_26 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  valid_27 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  valid_28 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  valid_29 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  valid_30 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  valid_31 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  valid_32 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  valid_33 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  valid_34 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  valid_35 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  valid_36 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  valid_37 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  valid_38 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  valid_39 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  valid_40 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  valid_41 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  valid_42 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  valid_43 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  valid_44 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  valid_45 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  valid_46 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  valid_47 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  valid_48 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  valid_49 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  valid_50 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  valid_51 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  valid_52 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  valid_53 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  valid_54 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  valid_55 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  valid_56 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  valid_57 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  valid_58 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  valid_59 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  valid_60 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  valid_61 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  valid_62 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  valid_63 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  valid_64 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  valid_65 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  valid_66 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  valid_67 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  valid_68 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  valid_69 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  valid_70 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  valid_71 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  valid_72 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  valid_73 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  valid_74 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  valid_75 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  valid_76 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  valid_77 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  valid_78 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  valid_79 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  valid_80 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  valid_81 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  valid_82 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  valid_83 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  valid_84 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  valid_85 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  valid_86 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  valid_87 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  valid_88 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  valid_89 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  valid_90 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  valid_91 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  valid_92 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  valid_93 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  valid_94 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  valid_95 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  valid_96 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  valid_97 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  valid_98 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  valid_99 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  valid_100 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  valid_101 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  valid_102 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  valid_103 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  valid_104 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  valid_105 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  valid_106 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  valid_107 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  valid_108 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  valid_109 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  valid_110 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  valid_111 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  valid_112 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  valid_113 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  valid_114 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  valid_115 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  valid_116 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  valid_117 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  valid_118 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  valid_119 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  valid_120 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  valid_121 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  valid_122 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  valid_123 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  valid_124 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  valid_125 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  valid_126 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  valid_127 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  valid_128 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  valid_129 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  valid_130 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  valid_131 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  valid_132 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  valid_133 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  valid_134 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  valid_135 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  valid_136 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  valid_137 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  valid_138 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  valid_139 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  valid_140 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  valid_141 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  valid_142 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  valid_143 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  valid_144 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  valid_145 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  valid_146 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  valid_147 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  valid_148 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  valid_149 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  valid_150 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  valid_151 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  valid_152 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  valid_153 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  valid_154 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  valid_155 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  valid_156 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  valid_157 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  valid_158 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  valid_159 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  valid_160 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  valid_161 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  valid_162 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  valid_163 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  valid_164 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  valid_165 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  valid_166 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  valid_167 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  valid_168 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  valid_169 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  valid_170 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  valid_171 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  valid_172 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  valid_173 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  valid_174 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  valid_175 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  valid_176 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  valid_177 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  valid_178 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  valid_179 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  valid_180 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  valid_181 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  valid_182 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  valid_183 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  valid_184 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  valid_185 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  valid_186 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  valid_187 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  valid_188 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  valid_189 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  valid_190 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  valid_191 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  valid_192 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  valid_193 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  valid_194 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  valid_195 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  valid_196 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  valid_197 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  valid_198 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  valid_199 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  valid_200 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  valid_201 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  valid_202 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  valid_203 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  valid_204 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  valid_205 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  valid_206 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  valid_207 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  valid_208 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  valid_209 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  valid_210 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  valid_211 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  valid_212 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  valid_213 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  valid_214 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  valid_215 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  valid_216 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  valid_217 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  valid_218 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  valid_219 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  valid_220 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  valid_221 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  valid_222 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  valid_223 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  valid_224 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  valid_225 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  valid_226 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  valid_227 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  valid_228 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  valid_229 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  valid_230 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  valid_231 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  valid_232 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  valid_233 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  valid_234 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  valid_235 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  valid_236 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  valid_237 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  valid_238 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  valid_239 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  valid_240 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  valid_241 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  valid_242 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  valid_243 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  valid_244 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  valid_245 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  valid_246 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  valid_247 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  valid_248 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  valid_249 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  valid_250 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  valid_251 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  valid_252 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  valid_253 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  valid_254 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  valid_255 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  valid_256 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  valid_257 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  valid_258 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  valid_259 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  valid_260 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  valid_261 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  valid_262 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  valid_263 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  valid_264 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  valid_265 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  valid_266 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  valid_267 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  valid_268 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  valid_269 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  valid_270 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  valid_271 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  valid_272 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  valid_273 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  valid_274 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  valid_275 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  valid_276 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  valid_277 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  valid_278 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  valid_279 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  valid_280 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  valid_281 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  valid_282 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  valid_283 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  valid_284 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  valid_285 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  valid_286 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  valid_287 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  valid_288 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  valid_289 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  valid_290 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  valid_291 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  valid_292 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  valid_293 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  valid_294 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  valid_295 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  valid_296 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  valid_297 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  valid_298 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  valid_299 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  valid_300 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  valid_301 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  valid_302 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  valid_303 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  valid_304 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  valid_305 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  valid_306 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  valid_307 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  valid_308 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  valid_309 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  valid_310 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  valid_311 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  valid_312 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  valid_313 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  valid_314 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  valid_315 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  valid_316 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  valid_317 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  valid_318 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  valid_319 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  valid_320 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  valid_321 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  valid_322 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  valid_323 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  valid_324 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  valid_325 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  valid_326 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  valid_327 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  valid_328 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  valid_329 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  valid_330 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  valid_331 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  valid_332 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  valid_333 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  valid_334 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  valid_335 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  valid_336 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  valid_337 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  valid_338 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  valid_339 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  valid_340 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  valid_341 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  valid_342 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  valid_343 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  valid_344 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  valid_345 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  valid_346 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  valid_347 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  valid_348 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  valid_349 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  valid_350 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  valid_351 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  valid_352 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  valid_353 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  valid_354 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  valid_355 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  valid_356 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  valid_357 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  valid_358 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  valid_359 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  valid_360 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  valid_361 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  valid_362 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  valid_363 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  valid_364 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  valid_365 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  valid_366 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  valid_367 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  valid_368 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  valid_369 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  valid_370 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  valid_371 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  valid_372 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  valid_373 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  valid_374 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  valid_375 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  valid_376 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  valid_377 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  valid_378 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  valid_379 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  valid_380 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  valid_381 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  valid_382 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  valid_383 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  valid_384 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  valid_385 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  valid_386 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  valid_387 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  valid_388 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  valid_389 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  valid_390 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  valid_391 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  valid_392 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  valid_393 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  valid_394 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  valid_395 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  valid_396 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  valid_397 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  valid_398 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  valid_399 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  valid_400 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  valid_401 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  valid_402 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  valid_403 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  valid_404 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  valid_405 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  valid_406 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  valid_407 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  valid_408 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  valid_409 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  valid_410 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  valid_411 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  valid_412 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  valid_413 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  valid_414 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  valid_415 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  valid_416 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  valid_417 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  valid_418 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  valid_419 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  valid_420 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  valid_421 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  valid_422 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  valid_423 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  valid_424 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  valid_425 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  valid_426 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  valid_427 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  valid_428 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  valid_429 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  valid_430 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  valid_431 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  valid_432 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  valid_433 = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  valid_434 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  valid_435 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  valid_436 = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  valid_437 = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  valid_438 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  valid_439 = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  valid_440 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  valid_441 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  valid_442 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  valid_443 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  valid_444 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  valid_445 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  valid_446 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  valid_447 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  valid_448 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  valid_449 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  valid_450 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  valid_451 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  valid_452 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  valid_453 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  valid_454 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  valid_455 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  valid_456 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  valid_457 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  valid_458 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  valid_459 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  valid_460 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  valid_461 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  valid_462 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  valid_463 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  valid_464 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  valid_465 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  valid_466 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  valid_467 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  valid_468 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  valid_469 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  valid_470 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  valid_471 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  valid_472 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  valid_473 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  valid_474 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  valid_475 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  valid_476 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  valid_477 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  valid_478 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  valid_479 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  valid_480 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  valid_481 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  valid_482 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  valid_483 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  valid_484 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  valid_485 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  valid_486 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  valid_487 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  valid_488 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  valid_489 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  valid_490 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  valid_491 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  valid_492 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  valid_493 = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  valid_494 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  valid_495 = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  valid_496 = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  valid_497 = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  valid_498 = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  valid_499 = _RAND_515[0:0];
  _RAND_516 = {1{`RANDOM}};
  valid_500 = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  valid_501 = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  valid_502 = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  valid_503 = _RAND_519[0:0];
  _RAND_520 = {1{`RANDOM}};
  valid_504 = _RAND_520[0:0];
  _RAND_521 = {1{`RANDOM}};
  valid_505 = _RAND_521[0:0];
  _RAND_522 = {1{`RANDOM}};
  valid_506 = _RAND_522[0:0];
  _RAND_523 = {1{`RANDOM}};
  valid_507 = _RAND_523[0:0];
  _RAND_524 = {1{`RANDOM}};
  valid_508 = _RAND_524[0:0];
  _RAND_525 = {1{`RANDOM}};
  valid_509 = _RAND_525[0:0];
  _RAND_526 = {1{`RANDOM}};
  valid_510 = _RAND_526[0:0];
  _RAND_527 = {1{`RANDOM}};
  valid_511 = _RAND_527[0:0];
  _RAND_528 = {1{`RANDOM}};
  valid_512 = _RAND_528[0:0];
  _RAND_529 = {1{`RANDOM}};
  valid_513 = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  valid_514 = _RAND_530[0:0];
  _RAND_531 = {1{`RANDOM}};
  valid_515 = _RAND_531[0:0];
  _RAND_532 = {1{`RANDOM}};
  valid_516 = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  valid_517 = _RAND_533[0:0];
  _RAND_534 = {1{`RANDOM}};
  valid_518 = _RAND_534[0:0];
  _RAND_535 = {1{`RANDOM}};
  valid_519 = _RAND_535[0:0];
  _RAND_536 = {1{`RANDOM}};
  valid_520 = _RAND_536[0:0];
  _RAND_537 = {1{`RANDOM}};
  valid_521 = _RAND_537[0:0];
  _RAND_538 = {1{`RANDOM}};
  valid_522 = _RAND_538[0:0];
  _RAND_539 = {1{`RANDOM}};
  valid_523 = _RAND_539[0:0];
  _RAND_540 = {1{`RANDOM}};
  valid_524 = _RAND_540[0:0];
  _RAND_541 = {1{`RANDOM}};
  valid_525 = _RAND_541[0:0];
  _RAND_542 = {1{`RANDOM}};
  valid_526 = _RAND_542[0:0];
  _RAND_543 = {1{`RANDOM}};
  valid_527 = _RAND_543[0:0];
  _RAND_544 = {1{`RANDOM}};
  valid_528 = _RAND_544[0:0];
  _RAND_545 = {1{`RANDOM}};
  valid_529 = _RAND_545[0:0];
  _RAND_546 = {1{`RANDOM}};
  valid_530 = _RAND_546[0:0];
  _RAND_547 = {1{`RANDOM}};
  valid_531 = _RAND_547[0:0];
  _RAND_548 = {1{`RANDOM}};
  valid_532 = _RAND_548[0:0];
  _RAND_549 = {1{`RANDOM}};
  valid_533 = _RAND_549[0:0];
  _RAND_550 = {1{`RANDOM}};
  valid_534 = _RAND_550[0:0];
  _RAND_551 = {1{`RANDOM}};
  valid_535 = _RAND_551[0:0];
  _RAND_552 = {1{`RANDOM}};
  valid_536 = _RAND_552[0:0];
  _RAND_553 = {1{`RANDOM}};
  valid_537 = _RAND_553[0:0];
  _RAND_554 = {1{`RANDOM}};
  valid_538 = _RAND_554[0:0];
  _RAND_555 = {1{`RANDOM}};
  valid_539 = _RAND_555[0:0];
  _RAND_556 = {1{`RANDOM}};
  valid_540 = _RAND_556[0:0];
  _RAND_557 = {1{`RANDOM}};
  valid_541 = _RAND_557[0:0];
  _RAND_558 = {1{`RANDOM}};
  valid_542 = _RAND_558[0:0];
  _RAND_559 = {1{`RANDOM}};
  valid_543 = _RAND_559[0:0];
  _RAND_560 = {1{`RANDOM}};
  valid_544 = _RAND_560[0:0];
  _RAND_561 = {1{`RANDOM}};
  valid_545 = _RAND_561[0:0];
  _RAND_562 = {1{`RANDOM}};
  valid_546 = _RAND_562[0:0];
  _RAND_563 = {1{`RANDOM}};
  valid_547 = _RAND_563[0:0];
  _RAND_564 = {1{`RANDOM}};
  valid_548 = _RAND_564[0:0];
  _RAND_565 = {1{`RANDOM}};
  valid_549 = _RAND_565[0:0];
  _RAND_566 = {1{`RANDOM}};
  valid_550 = _RAND_566[0:0];
  _RAND_567 = {1{`RANDOM}};
  valid_551 = _RAND_567[0:0];
  _RAND_568 = {1{`RANDOM}};
  valid_552 = _RAND_568[0:0];
  _RAND_569 = {1{`RANDOM}};
  valid_553 = _RAND_569[0:0];
  _RAND_570 = {1{`RANDOM}};
  valid_554 = _RAND_570[0:0];
  _RAND_571 = {1{`RANDOM}};
  valid_555 = _RAND_571[0:0];
  _RAND_572 = {1{`RANDOM}};
  valid_556 = _RAND_572[0:0];
  _RAND_573 = {1{`RANDOM}};
  valid_557 = _RAND_573[0:0];
  _RAND_574 = {1{`RANDOM}};
  valid_558 = _RAND_574[0:0];
  _RAND_575 = {1{`RANDOM}};
  valid_559 = _RAND_575[0:0];
  _RAND_576 = {1{`RANDOM}};
  valid_560 = _RAND_576[0:0];
  _RAND_577 = {1{`RANDOM}};
  valid_561 = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  valid_562 = _RAND_578[0:0];
  _RAND_579 = {1{`RANDOM}};
  valid_563 = _RAND_579[0:0];
  _RAND_580 = {1{`RANDOM}};
  valid_564 = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  valid_565 = _RAND_581[0:0];
  _RAND_582 = {1{`RANDOM}};
  valid_566 = _RAND_582[0:0];
  _RAND_583 = {1{`RANDOM}};
  valid_567 = _RAND_583[0:0];
  _RAND_584 = {1{`RANDOM}};
  valid_568 = _RAND_584[0:0];
  _RAND_585 = {1{`RANDOM}};
  valid_569 = _RAND_585[0:0];
  _RAND_586 = {1{`RANDOM}};
  valid_570 = _RAND_586[0:0];
  _RAND_587 = {1{`RANDOM}};
  valid_571 = _RAND_587[0:0];
  _RAND_588 = {1{`RANDOM}};
  valid_572 = _RAND_588[0:0];
  _RAND_589 = {1{`RANDOM}};
  valid_573 = _RAND_589[0:0];
  _RAND_590 = {1{`RANDOM}};
  valid_574 = _RAND_590[0:0];
  _RAND_591 = {1{`RANDOM}};
  valid_575 = _RAND_591[0:0];
  _RAND_592 = {1{`RANDOM}};
  valid_576 = _RAND_592[0:0];
  _RAND_593 = {1{`RANDOM}};
  valid_577 = _RAND_593[0:0];
  _RAND_594 = {1{`RANDOM}};
  valid_578 = _RAND_594[0:0];
  _RAND_595 = {1{`RANDOM}};
  valid_579 = _RAND_595[0:0];
  _RAND_596 = {1{`RANDOM}};
  valid_580 = _RAND_596[0:0];
  _RAND_597 = {1{`RANDOM}};
  valid_581 = _RAND_597[0:0];
  _RAND_598 = {1{`RANDOM}};
  valid_582 = _RAND_598[0:0];
  _RAND_599 = {1{`RANDOM}};
  valid_583 = _RAND_599[0:0];
  _RAND_600 = {1{`RANDOM}};
  valid_584 = _RAND_600[0:0];
  _RAND_601 = {1{`RANDOM}};
  valid_585 = _RAND_601[0:0];
  _RAND_602 = {1{`RANDOM}};
  valid_586 = _RAND_602[0:0];
  _RAND_603 = {1{`RANDOM}};
  valid_587 = _RAND_603[0:0];
  _RAND_604 = {1{`RANDOM}};
  valid_588 = _RAND_604[0:0];
  _RAND_605 = {1{`RANDOM}};
  valid_589 = _RAND_605[0:0];
  _RAND_606 = {1{`RANDOM}};
  valid_590 = _RAND_606[0:0];
  _RAND_607 = {1{`RANDOM}};
  valid_591 = _RAND_607[0:0];
  _RAND_608 = {1{`RANDOM}};
  valid_592 = _RAND_608[0:0];
  _RAND_609 = {1{`RANDOM}};
  valid_593 = _RAND_609[0:0];
  _RAND_610 = {1{`RANDOM}};
  valid_594 = _RAND_610[0:0];
  _RAND_611 = {1{`RANDOM}};
  valid_595 = _RAND_611[0:0];
  _RAND_612 = {1{`RANDOM}};
  valid_596 = _RAND_612[0:0];
  _RAND_613 = {1{`RANDOM}};
  valid_597 = _RAND_613[0:0];
  _RAND_614 = {1{`RANDOM}};
  valid_598 = _RAND_614[0:0];
  _RAND_615 = {1{`RANDOM}};
  valid_599 = _RAND_615[0:0];
  _RAND_616 = {1{`RANDOM}};
  valid_600 = _RAND_616[0:0];
  _RAND_617 = {1{`RANDOM}};
  valid_601 = _RAND_617[0:0];
  _RAND_618 = {1{`RANDOM}};
  valid_602 = _RAND_618[0:0];
  _RAND_619 = {1{`RANDOM}};
  valid_603 = _RAND_619[0:0];
  _RAND_620 = {1{`RANDOM}};
  valid_604 = _RAND_620[0:0];
  _RAND_621 = {1{`RANDOM}};
  valid_605 = _RAND_621[0:0];
  _RAND_622 = {1{`RANDOM}};
  valid_606 = _RAND_622[0:0];
  _RAND_623 = {1{`RANDOM}};
  valid_607 = _RAND_623[0:0];
  _RAND_624 = {1{`RANDOM}};
  valid_608 = _RAND_624[0:0];
  _RAND_625 = {1{`RANDOM}};
  valid_609 = _RAND_625[0:0];
  _RAND_626 = {1{`RANDOM}};
  valid_610 = _RAND_626[0:0];
  _RAND_627 = {1{`RANDOM}};
  valid_611 = _RAND_627[0:0];
  _RAND_628 = {1{`RANDOM}};
  valid_612 = _RAND_628[0:0];
  _RAND_629 = {1{`RANDOM}};
  valid_613 = _RAND_629[0:0];
  _RAND_630 = {1{`RANDOM}};
  valid_614 = _RAND_630[0:0];
  _RAND_631 = {1{`RANDOM}};
  valid_615 = _RAND_631[0:0];
  _RAND_632 = {1{`RANDOM}};
  valid_616 = _RAND_632[0:0];
  _RAND_633 = {1{`RANDOM}};
  valid_617 = _RAND_633[0:0];
  _RAND_634 = {1{`RANDOM}};
  valid_618 = _RAND_634[0:0];
  _RAND_635 = {1{`RANDOM}};
  valid_619 = _RAND_635[0:0];
  _RAND_636 = {1{`RANDOM}};
  valid_620 = _RAND_636[0:0];
  _RAND_637 = {1{`RANDOM}};
  valid_621 = _RAND_637[0:0];
  _RAND_638 = {1{`RANDOM}};
  valid_622 = _RAND_638[0:0];
  _RAND_639 = {1{`RANDOM}};
  valid_623 = _RAND_639[0:0];
  _RAND_640 = {1{`RANDOM}};
  valid_624 = _RAND_640[0:0];
  _RAND_641 = {1{`RANDOM}};
  valid_625 = _RAND_641[0:0];
  _RAND_642 = {1{`RANDOM}};
  valid_626 = _RAND_642[0:0];
  _RAND_643 = {1{`RANDOM}};
  valid_627 = _RAND_643[0:0];
  _RAND_644 = {1{`RANDOM}};
  valid_628 = _RAND_644[0:0];
  _RAND_645 = {1{`RANDOM}};
  valid_629 = _RAND_645[0:0];
  _RAND_646 = {1{`RANDOM}};
  valid_630 = _RAND_646[0:0];
  _RAND_647 = {1{`RANDOM}};
  valid_631 = _RAND_647[0:0];
  _RAND_648 = {1{`RANDOM}};
  valid_632 = _RAND_648[0:0];
  _RAND_649 = {1{`RANDOM}};
  valid_633 = _RAND_649[0:0];
  _RAND_650 = {1{`RANDOM}};
  valid_634 = _RAND_650[0:0];
  _RAND_651 = {1{`RANDOM}};
  valid_635 = _RAND_651[0:0];
  _RAND_652 = {1{`RANDOM}};
  valid_636 = _RAND_652[0:0];
  _RAND_653 = {1{`RANDOM}};
  valid_637 = _RAND_653[0:0];
  _RAND_654 = {1{`RANDOM}};
  valid_638 = _RAND_654[0:0];
  _RAND_655 = {1{`RANDOM}};
  valid_639 = _RAND_655[0:0];
  _RAND_656 = {1{`RANDOM}};
  valid_640 = _RAND_656[0:0];
  _RAND_657 = {1{`RANDOM}};
  valid_641 = _RAND_657[0:0];
  _RAND_658 = {1{`RANDOM}};
  valid_642 = _RAND_658[0:0];
  _RAND_659 = {1{`RANDOM}};
  valid_643 = _RAND_659[0:0];
  _RAND_660 = {1{`RANDOM}};
  valid_644 = _RAND_660[0:0];
  _RAND_661 = {1{`RANDOM}};
  valid_645 = _RAND_661[0:0];
  _RAND_662 = {1{`RANDOM}};
  valid_646 = _RAND_662[0:0];
  _RAND_663 = {1{`RANDOM}};
  valid_647 = _RAND_663[0:0];
  _RAND_664 = {1{`RANDOM}};
  valid_648 = _RAND_664[0:0];
  _RAND_665 = {1{`RANDOM}};
  valid_649 = _RAND_665[0:0];
  _RAND_666 = {1{`RANDOM}};
  valid_650 = _RAND_666[0:0];
  _RAND_667 = {1{`RANDOM}};
  valid_651 = _RAND_667[0:0];
  _RAND_668 = {1{`RANDOM}};
  valid_652 = _RAND_668[0:0];
  _RAND_669 = {1{`RANDOM}};
  valid_653 = _RAND_669[0:0];
  _RAND_670 = {1{`RANDOM}};
  valid_654 = _RAND_670[0:0];
  _RAND_671 = {1{`RANDOM}};
  valid_655 = _RAND_671[0:0];
  _RAND_672 = {1{`RANDOM}};
  valid_656 = _RAND_672[0:0];
  _RAND_673 = {1{`RANDOM}};
  valid_657 = _RAND_673[0:0];
  _RAND_674 = {1{`RANDOM}};
  valid_658 = _RAND_674[0:0];
  _RAND_675 = {1{`RANDOM}};
  valid_659 = _RAND_675[0:0];
  _RAND_676 = {1{`RANDOM}};
  valid_660 = _RAND_676[0:0];
  _RAND_677 = {1{`RANDOM}};
  valid_661 = _RAND_677[0:0];
  _RAND_678 = {1{`RANDOM}};
  valid_662 = _RAND_678[0:0];
  _RAND_679 = {1{`RANDOM}};
  valid_663 = _RAND_679[0:0];
  _RAND_680 = {1{`RANDOM}};
  valid_664 = _RAND_680[0:0];
  _RAND_681 = {1{`RANDOM}};
  valid_665 = _RAND_681[0:0];
  _RAND_682 = {1{`RANDOM}};
  valid_666 = _RAND_682[0:0];
  _RAND_683 = {1{`RANDOM}};
  valid_667 = _RAND_683[0:0];
  _RAND_684 = {1{`RANDOM}};
  valid_668 = _RAND_684[0:0];
  _RAND_685 = {1{`RANDOM}};
  valid_669 = _RAND_685[0:0];
  _RAND_686 = {1{`RANDOM}};
  valid_670 = _RAND_686[0:0];
  _RAND_687 = {1{`RANDOM}};
  valid_671 = _RAND_687[0:0];
  _RAND_688 = {1{`RANDOM}};
  valid_672 = _RAND_688[0:0];
  _RAND_689 = {1{`RANDOM}};
  valid_673 = _RAND_689[0:0];
  _RAND_690 = {1{`RANDOM}};
  valid_674 = _RAND_690[0:0];
  _RAND_691 = {1{`RANDOM}};
  valid_675 = _RAND_691[0:0];
  _RAND_692 = {1{`RANDOM}};
  valid_676 = _RAND_692[0:0];
  _RAND_693 = {1{`RANDOM}};
  valid_677 = _RAND_693[0:0];
  _RAND_694 = {1{`RANDOM}};
  valid_678 = _RAND_694[0:0];
  _RAND_695 = {1{`RANDOM}};
  valid_679 = _RAND_695[0:0];
  _RAND_696 = {1{`RANDOM}};
  valid_680 = _RAND_696[0:0];
  _RAND_697 = {1{`RANDOM}};
  valid_681 = _RAND_697[0:0];
  _RAND_698 = {1{`RANDOM}};
  valid_682 = _RAND_698[0:0];
  _RAND_699 = {1{`RANDOM}};
  valid_683 = _RAND_699[0:0];
  _RAND_700 = {1{`RANDOM}};
  valid_684 = _RAND_700[0:0];
  _RAND_701 = {1{`RANDOM}};
  valid_685 = _RAND_701[0:0];
  _RAND_702 = {1{`RANDOM}};
  valid_686 = _RAND_702[0:0];
  _RAND_703 = {1{`RANDOM}};
  valid_687 = _RAND_703[0:0];
  _RAND_704 = {1{`RANDOM}};
  valid_688 = _RAND_704[0:0];
  _RAND_705 = {1{`RANDOM}};
  valid_689 = _RAND_705[0:0];
  _RAND_706 = {1{`RANDOM}};
  valid_690 = _RAND_706[0:0];
  _RAND_707 = {1{`RANDOM}};
  valid_691 = _RAND_707[0:0];
  _RAND_708 = {1{`RANDOM}};
  valid_692 = _RAND_708[0:0];
  _RAND_709 = {1{`RANDOM}};
  valid_693 = _RAND_709[0:0];
  _RAND_710 = {1{`RANDOM}};
  valid_694 = _RAND_710[0:0];
  _RAND_711 = {1{`RANDOM}};
  valid_695 = _RAND_711[0:0];
  _RAND_712 = {1{`RANDOM}};
  valid_696 = _RAND_712[0:0];
  _RAND_713 = {1{`RANDOM}};
  valid_697 = _RAND_713[0:0];
  _RAND_714 = {1{`RANDOM}};
  valid_698 = _RAND_714[0:0];
  _RAND_715 = {1{`RANDOM}};
  valid_699 = _RAND_715[0:0];
  _RAND_716 = {1{`RANDOM}};
  valid_700 = _RAND_716[0:0];
  _RAND_717 = {1{`RANDOM}};
  valid_701 = _RAND_717[0:0];
  _RAND_718 = {1{`RANDOM}};
  valid_702 = _RAND_718[0:0];
  _RAND_719 = {1{`RANDOM}};
  valid_703 = _RAND_719[0:0];
  _RAND_720 = {1{`RANDOM}};
  valid_704 = _RAND_720[0:0];
  _RAND_721 = {1{`RANDOM}};
  valid_705 = _RAND_721[0:0];
  _RAND_722 = {1{`RANDOM}};
  valid_706 = _RAND_722[0:0];
  _RAND_723 = {1{`RANDOM}};
  valid_707 = _RAND_723[0:0];
  _RAND_724 = {1{`RANDOM}};
  valid_708 = _RAND_724[0:0];
  _RAND_725 = {1{`RANDOM}};
  valid_709 = _RAND_725[0:0];
  _RAND_726 = {1{`RANDOM}};
  valid_710 = _RAND_726[0:0];
  _RAND_727 = {1{`RANDOM}};
  valid_711 = _RAND_727[0:0];
  _RAND_728 = {1{`RANDOM}};
  valid_712 = _RAND_728[0:0];
  _RAND_729 = {1{`RANDOM}};
  valid_713 = _RAND_729[0:0];
  _RAND_730 = {1{`RANDOM}};
  valid_714 = _RAND_730[0:0];
  _RAND_731 = {1{`RANDOM}};
  valid_715 = _RAND_731[0:0];
  _RAND_732 = {1{`RANDOM}};
  valid_716 = _RAND_732[0:0];
  _RAND_733 = {1{`RANDOM}};
  valid_717 = _RAND_733[0:0];
  _RAND_734 = {1{`RANDOM}};
  valid_718 = _RAND_734[0:0];
  _RAND_735 = {1{`RANDOM}};
  valid_719 = _RAND_735[0:0];
  _RAND_736 = {1{`RANDOM}};
  valid_720 = _RAND_736[0:0];
  _RAND_737 = {1{`RANDOM}};
  valid_721 = _RAND_737[0:0];
  _RAND_738 = {1{`RANDOM}};
  valid_722 = _RAND_738[0:0];
  _RAND_739 = {1{`RANDOM}};
  valid_723 = _RAND_739[0:0];
  _RAND_740 = {1{`RANDOM}};
  valid_724 = _RAND_740[0:0];
  _RAND_741 = {1{`RANDOM}};
  valid_725 = _RAND_741[0:0];
  _RAND_742 = {1{`RANDOM}};
  valid_726 = _RAND_742[0:0];
  _RAND_743 = {1{`RANDOM}};
  valid_727 = _RAND_743[0:0];
  _RAND_744 = {1{`RANDOM}};
  valid_728 = _RAND_744[0:0];
  _RAND_745 = {1{`RANDOM}};
  valid_729 = _RAND_745[0:0];
  _RAND_746 = {1{`RANDOM}};
  valid_730 = _RAND_746[0:0];
  _RAND_747 = {1{`RANDOM}};
  valid_731 = _RAND_747[0:0];
  _RAND_748 = {1{`RANDOM}};
  valid_732 = _RAND_748[0:0];
  _RAND_749 = {1{`RANDOM}};
  valid_733 = _RAND_749[0:0];
  _RAND_750 = {1{`RANDOM}};
  valid_734 = _RAND_750[0:0];
  _RAND_751 = {1{`RANDOM}};
  valid_735 = _RAND_751[0:0];
  _RAND_752 = {1{`RANDOM}};
  valid_736 = _RAND_752[0:0];
  _RAND_753 = {1{`RANDOM}};
  valid_737 = _RAND_753[0:0];
  _RAND_754 = {1{`RANDOM}};
  valid_738 = _RAND_754[0:0];
  _RAND_755 = {1{`RANDOM}};
  valid_739 = _RAND_755[0:0];
  _RAND_756 = {1{`RANDOM}};
  valid_740 = _RAND_756[0:0];
  _RAND_757 = {1{`RANDOM}};
  valid_741 = _RAND_757[0:0];
  _RAND_758 = {1{`RANDOM}};
  valid_742 = _RAND_758[0:0];
  _RAND_759 = {1{`RANDOM}};
  valid_743 = _RAND_759[0:0];
  _RAND_760 = {1{`RANDOM}};
  valid_744 = _RAND_760[0:0];
  _RAND_761 = {1{`RANDOM}};
  valid_745 = _RAND_761[0:0];
  _RAND_762 = {1{`RANDOM}};
  valid_746 = _RAND_762[0:0];
  _RAND_763 = {1{`RANDOM}};
  valid_747 = _RAND_763[0:0];
  _RAND_764 = {1{`RANDOM}};
  valid_748 = _RAND_764[0:0];
  _RAND_765 = {1{`RANDOM}};
  valid_749 = _RAND_765[0:0];
  _RAND_766 = {1{`RANDOM}};
  valid_750 = _RAND_766[0:0];
  _RAND_767 = {1{`RANDOM}};
  valid_751 = _RAND_767[0:0];
  _RAND_768 = {1{`RANDOM}};
  valid_752 = _RAND_768[0:0];
  _RAND_769 = {1{`RANDOM}};
  valid_753 = _RAND_769[0:0];
  _RAND_770 = {1{`RANDOM}};
  valid_754 = _RAND_770[0:0];
  _RAND_771 = {1{`RANDOM}};
  valid_755 = _RAND_771[0:0];
  _RAND_772 = {1{`RANDOM}};
  valid_756 = _RAND_772[0:0];
  _RAND_773 = {1{`RANDOM}};
  valid_757 = _RAND_773[0:0];
  _RAND_774 = {1{`RANDOM}};
  valid_758 = _RAND_774[0:0];
  _RAND_775 = {1{`RANDOM}};
  valid_759 = _RAND_775[0:0];
  _RAND_776 = {1{`RANDOM}};
  valid_760 = _RAND_776[0:0];
  _RAND_777 = {1{`RANDOM}};
  valid_761 = _RAND_777[0:0];
  _RAND_778 = {1{`RANDOM}};
  valid_762 = _RAND_778[0:0];
  _RAND_779 = {1{`RANDOM}};
  valid_763 = _RAND_779[0:0];
  _RAND_780 = {1{`RANDOM}};
  valid_764 = _RAND_780[0:0];
  _RAND_781 = {1{`RANDOM}};
  valid_765 = _RAND_781[0:0];
  _RAND_782 = {1{`RANDOM}};
  valid_766 = _RAND_782[0:0];
  _RAND_783 = {1{`RANDOM}};
  valid_767 = _RAND_783[0:0];
  _RAND_784 = {1{`RANDOM}};
  valid_768 = _RAND_784[0:0];
  _RAND_785 = {1{`RANDOM}};
  valid_769 = _RAND_785[0:0];
  _RAND_786 = {1{`RANDOM}};
  valid_770 = _RAND_786[0:0];
  _RAND_787 = {1{`RANDOM}};
  valid_771 = _RAND_787[0:0];
  _RAND_788 = {1{`RANDOM}};
  valid_772 = _RAND_788[0:0];
  _RAND_789 = {1{`RANDOM}};
  valid_773 = _RAND_789[0:0];
  _RAND_790 = {1{`RANDOM}};
  valid_774 = _RAND_790[0:0];
  _RAND_791 = {1{`RANDOM}};
  valid_775 = _RAND_791[0:0];
  _RAND_792 = {1{`RANDOM}};
  valid_776 = _RAND_792[0:0];
  _RAND_793 = {1{`RANDOM}};
  valid_777 = _RAND_793[0:0];
  _RAND_794 = {1{`RANDOM}};
  valid_778 = _RAND_794[0:0];
  _RAND_795 = {1{`RANDOM}};
  valid_779 = _RAND_795[0:0];
  _RAND_796 = {1{`RANDOM}};
  valid_780 = _RAND_796[0:0];
  _RAND_797 = {1{`RANDOM}};
  valid_781 = _RAND_797[0:0];
  _RAND_798 = {1{`RANDOM}};
  valid_782 = _RAND_798[0:0];
  _RAND_799 = {1{`RANDOM}};
  valid_783 = _RAND_799[0:0];
  _RAND_800 = {1{`RANDOM}};
  valid_784 = _RAND_800[0:0];
  _RAND_801 = {1{`RANDOM}};
  valid_785 = _RAND_801[0:0];
  _RAND_802 = {1{`RANDOM}};
  valid_786 = _RAND_802[0:0];
  _RAND_803 = {1{`RANDOM}};
  valid_787 = _RAND_803[0:0];
  _RAND_804 = {1{`RANDOM}};
  valid_788 = _RAND_804[0:0];
  _RAND_805 = {1{`RANDOM}};
  valid_789 = _RAND_805[0:0];
  _RAND_806 = {1{`RANDOM}};
  valid_790 = _RAND_806[0:0];
  _RAND_807 = {1{`RANDOM}};
  valid_791 = _RAND_807[0:0];
  _RAND_808 = {1{`RANDOM}};
  valid_792 = _RAND_808[0:0];
  _RAND_809 = {1{`RANDOM}};
  valid_793 = _RAND_809[0:0];
  _RAND_810 = {1{`RANDOM}};
  valid_794 = _RAND_810[0:0];
  _RAND_811 = {1{`RANDOM}};
  valid_795 = _RAND_811[0:0];
  _RAND_812 = {1{`RANDOM}};
  valid_796 = _RAND_812[0:0];
  _RAND_813 = {1{`RANDOM}};
  valid_797 = _RAND_813[0:0];
  _RAND_814 = {1{`RANDOM}};
  valid_798 = _RAND_814[0:0];
  _RAND_815 = {1{`RANDOM}};
  valid_799 = _RAND_815[0:0];
  _RAND_816 = {1{`RANDOM}};
  valid_800 = _RAND_816[0:0];
  _RAND_817 = {1{`RANDOM}};
  valid_801 = _RAND_817[0:0];
  _RAND_818 = {1{`RANDOM}};
  valid_802 = _RAND_818[0:0];
  _RAND_819 = {1{`RANDOM}};
  valid_803 = _RAND_819[0:0];
  _RAND_820 = {1{`RANDOM}};
  valid_804 = _RAND_820[0:0];
  _RAND_821 = {1{`RANDOM}};
  valid_805 = _RAND_821[0:0];
  _RAND_822 = {1{`RANDOM}};
  valid_806 = _RAND_822[0:0];
  _RAND_823 = {1{`RANDOM}};
  valid_807 = _RAND_823[0:0];
  _RAND_824 = {1{`RANDOM}};
  valid_808 = _RAND_824[0:0];
  _RAND_825 = {1{`RANDOM}};
  valid_809 = _RAND_825[0:0];
  _RAND_826 = {1{`RANDOM}};
  valid_810 = _RAND_826[0:0];
  _RAND_827 = {1{`RANDOM}};
  valid_811 = _RAND_827[0:0];
  _RAND_828 = {1{`RANDOM}};
  valid_812 = _RAND_828[0:0];
  _RAND_829 = {1{`RANDOM}};
  valid_813 = _RAND_829[0:0];
  _RAND_830 = {1{`RANDOM}};
  valid_814 = _RAND_830[0:0];
  _RAND_831 = {1{`RANDOM}};
  valid_815 = _RAND_831[0:0];
  _RAND_832 = {1{`RANDOM}};
  valid_816 = _RAND_832[0:0];
  _RAND_833 = {1{`RANDOM}};
  valid_817 = _RAND_833[0:0];
  _RAND_834 = {1{`RANDOM}};
  valid_818 = _RAND_834[0:0];
  _RAND_835 = {1{`RANDOM}};
  valid_819 = _RAND_835[0:0];
  _RAND_836 = {1{`RANDOM}};
  valid_820 = _RAND_836[0:0];
  _RAND_837 = {1{`RANDOM}};
  valid_821 = _RAND_837[0:0];
  _RAND_838 = {1{`RANDOM}};
  valid_822 = _RAND_838[0:0];
  _RAND_839 = {1{`RANDOM}};
  valid_823 = _RAND_839[0:0];
  _RAND_840 = {1{`RANDOM}};
  valid_824 = _RAND_840[0:0];
  _RAND_841 = {1{`RANDOM}};
  valid_825 = _RAND_841[0:0];
  _RAND_842 = {1{`RANDOM}};
  valid_826 = _RAND_842[0:0];
  _RAND_843 = {1{`RANDOM}};
  valid_827 = _RAND_843[0:0];
  _RAND_844 = {1{`RANDOM}};
  valid_828 = _RAND_844[0:0];
  _RAND_845 = {1{`RANDOM}};
  valid_829 = _RAND_845[0:0];
  _RAND_846 = {1{`RANDOM}};
  valid_830 = _RAND_846[0:0];
  _RAND_847 = {1{`RANDOM}};
  valid_831 = _RAND_847[0:0];
  _RAND_848 = {1{`RANDOM}};
  valid_832 = _RAND_848[0:0];
  _RAND_849 = {1{`RANDOM}};
  valid_833 = _RAND_849[0:0];
  _RAND_850 = {1{`RANDOM}};
  valid_834 = _RAND_850[0:0];
  _RAND_851 = {1{`RANDOM}};
  valid_835 = _RAND_851[0:0];
  _RAND_852 = {1{`RANDOM}};
  valid_836 = _RAND_852[0:0];
  _RAND_853 = {1{`RANDOM}};
  valid_837 = _RAND_853[0:0];
  _RAND_854 = {1{`RANDOM}};
  valid_838 = _RAND_854[0:0];
  _RAND_855 = {1{`RANDOM}};
  valid_839 = _RAND_855[0:0];
  _RAND_856 = {1{`RANDOM}};
  valid_840 = _RAND_856[0:0];
  _RAND_857 = {1{`RANDOM}};
  valid_841 = _RAND_857[0:0];
  _RAND_858 = {1{`RANDOM}};
  valid_842 = _RAND_858[0:0];
  _RAND_859 = {1{`RANDOM}};
  valid_843 = _RAND_859[0:0];
  _RAND_860 = {1{`RANDOM}};
  valid_844 = _RAND_860[0:0];
  _RAND_861 = {1{`RANDOM}};
  valid_845 = _RAND_861[0:0];
  _RAND_862 = {1{`RANDOM}};
  valid_846 = _RAND_862[0:0];
  _RAND_863 = {1{`RANDOM}};
  valid_847 = _RAND_863[0:0];
  _RAND_864 = {1{`RANDOM}};
  valid_848 = _RAND_864[0:0];
  _RAND_865 = {1{`RANDOM}};
  valid_849 = _RAND_865[0:0];
  _RAND_866 = {1{`RANDOM}};
  valid_850 = _RAND_866[0:0];
  _RAND_867 = {1{`RANDOM}};
  valid_851 = _RAND_867[0:0];
  _RAND_868 = {1{`RANDOM}};
  valid_852 = _RAND_868[0:0];
  _RAND_869 = {1{`RANDOM}};
  valid_853 = _RAND_869[0:0];
  _RAND_870 = {1{`RANDOM}};
  valid_854 = _RAND_870[0:0];
  _RAND_871 = {1{`RANDOM}};
  valid_855 = _RAND_871[0:0];
  _RAND_872 = {1{`RANDOM}};
  valid_856 = _RAND_872[0:0];
  _RAND_873 = {1{`RANDOM}};
  valid_857 = _RAND_873[0:0];
  _RAND_874 = {1{`RANDOM}};
  valid_858 = _RAND_874[0:0];
  _RAND_875 = {1{`RANDOM}};
  valid_859 = _RAND_875[0:0];
  _RAND_876 = {1{`RANDOM}};
  valid_860 = _RAND_876[0:0];
  _RAND_877 = {1{`RANDOM}};
  valid_861 = _RAND_877[0:0];
  _RAND_878 = {1{`RANDOM}};
  valid_862 = _RAND_878[0:0];
  _RAND_879 = {1{`RANDOM}};
  valid_863 = _RAND_879[0:0];
  _RAND_880 = {1{`RANDOM}};
  valid_864 = _RAND_880[0:0];
  _RAND_881 = {1{`RANDOM}};
  valid_865 = _RAND_881[0:0];
  _RAND_882 = {1{`RANDOM}};
  valid_866 = _RAND_882[0:0];
  _RAND_883 = {1{`RANDOM}};
  valid_867 = _RAND_883[0:0];
  _RAND_884 = {1{`RANDOM}};
  valid_868 = _RAND_884[0:0];
  _RAND_885 = {1{`RANDOM}};
  valid_869 = _RAND_885[0:0];
  _RAND_886 = {1{`RANDOM}};
  valid_870 = _RAND_886[0:0];
  _RAND_887 = {1{`RANDOM}};
  valid_871 = _RAND_887[0:0];
  _RAND_888 = {1{`RANDOM}};
  valid_872 = _RAND_888[0:0];
  _RAND_889 = {1{`RANDOM}};
  valid_873 = _RAND_889[0:0];
  _RAND_890 = {1{`RANDOM}};
  valid_874 = _RAND_890[0:0];
  _RAND_891 = {1{`RANDOM}};
  valid_875 = _RAND_891[0:0];
  _RAND_892 = {1{`RANDOM}};
  valid_876 = _RAND_892[0:0];
  _RAND_893 = {1{`RANDOM}};
  valid_877 = _RAND_893[0:0];
  _RAND_894 = {1{`RANDOM}};
  valid_878 = _RAND_894[0:0];
  _RAND_895 = {1{`RANDOM}};
  valid_879 = _RAND_895[0:0];
  _RAND_896 = {1{`RANDOM}};
  valid_880 = _RAND_896[0:0];
  _RAND_897 = {1{`RANDOM}};
  valid_881 = _RAND_897[0:0];
  _RAND_898 = {1{`RANDOM}};
  valid_882 = _RAND_898[0:0];
  _RAND_899 = {1{`RANDOM}};
  valid_883 = _RAND_899[0:0];
  _RAND_900 = {1{`RANDOM}};
  valid_884 = _RAND_900[0:0];
  _RAND_901 = {1{`RANDOM}};
  valid_885 = _RAND_901[0:0];
  _RAND_902 = {1{`RANDOM}};
  valid_886 = _RAND_902[0:0];
  _RAND_903 = {1{`RANDOM}};
  valid_887 = _RAND_903[0:0];
  _RAND_904 = {1{`RANDOM}};
  valid_888 = _RAND_904[0:0];
  _RAND_905 = {1{`RANDOM}};
  valid_889 = _RAND_905[0:0];
  _RAND_906 = {1{`RANDOM}};
  valid_890 = _RAND_906[0:0];
  _RAND_907 = {1{`RANDOM}};
  valid_891 = _RAND_907[0:0];
  _RAND_908 = {1{`RANDOM}};
  valid_892 = _RAND_908[0:0];
  _RAND_909 = {1{`RANDOM}};
  valid_893 = _RAND_909[0:0];
  _RAND_910 = {1{`RANDOM}};
  valid_894 = _RAND_910[0:0];
  _RAND_911 = {1{`RANDOM}};
  valid_895 = _RAND_911[0:0];
  _RAND_912 = {1{`RANDOM}};
  valid_896 = _RAND_912[0:0];
  _RAND_913 = {1{`RANDOM}};
  valid_897 = _RAND_913[0:0];
  _RAND_914 = {1{`RANDOM}};
  valid_898 = _RAND_914[0:0];
  _RAND_915 = {1{`RANDOM}};
  valid_899 = _RAND_915[0:0];
  _RAND_916 = {1{`RANDOM}};
  valid_900 = _RAND_916[0:0];
  _RAND_917 = {1{`RANDOM}};
  valid_901 = _RAND_917[0:0];
  _RAND_918 = {1{`RANDOM}};
  valid_902 = _RAND_918[0:0];
  _RAND_919 = {1{`RANDOM}};
  valid_903 = _RAND_919[0:0];
  _RAND_920 = {1{`RANDOM}};
  valid_904 = _RAND_920[0:0];
  _RAND_921 = {1{`RANDOM}};
  valid_905 = _RAND_921[0:0];
  _RAND_922 = {1{`RANDOM}};
  valid_906 = _RAND_922[0:0];
  _RAND_923 = {1{`RANDOM}};
  valid_907 = _RAND_923[0:0];
  _RAND_924 = {1{`RANDOM}};
  valid_908 = _RAND_924[0:0];
  _RAND_925 = {1{`RANDOM}};
  valid_909 = _RAND_925[0:0];
  _RAND_926 = {1{`RANDOM}};
  valid_910 = _RAND_926[0:0];
  _RAND_927 = {1{`RANDOM}};
  valid_911 = _RAND_927[0:0];
  _RAND_928 = {1{`RANDOM}};
  valid_912 = _RAND_928[0:0];
  _RAND_929 = {1{`RANDOM}};
  valid_913 = _RAND_929[0:0];
  _RAND_930 = {1{`RANDOM}};
  valid_914 = _RAND_930[0:0];
  _RAND_931 = {1{`RANDOM}};
  valid_915 = _RAND_931[0:0];
  _RAND_932 = {1{`RANDOM}};
  valid_916 = _RAND_932[0:0];
  _RAND_933 = {1{`RANDOM}};
  valid_917 = _RAND_933[0:0];
  _RAND_934 = {1{`RANDOM}};
  valid_918 = _RAND_934[0:0];
  _RAND_935 = {1{`RANDOM}};
  valid_919 = _RAND_935[0:0];
  _RAND_936 = {1{`RANDOM}};
  valid_920 = _RAND_936[0:0];
  _RAND_937 = {1{`RANDOM}};
  valid_921 = _RAND_937[0:0];
  _RAND_938 = {1{`RANDOM}};
  valid_922 = _RAND_938[0:0];
  _RAND_939 = {1{`RANDOM}};
  valid_923 = _RAND_939[0:0];
  _RAND_940 = {1{`RANDOM}};
  valid_924 = _RAND_940[0:0];
  _RAND_941 = {1{`RANDOM}};
  valid_925 = _RAND_941[0:0];
  _RAND_942 = {1{`RANDOM}};
  valid_926 = _RAND_942[0:0];
  _RAND_943 = {1{`RANDOM}};
  valid_927 = _RAND_943[0:0];
  _RAND_944 = {1{`RANDOM}};
  valid_928 = _RAND_944[0:0];
  _RAND_945 = {1{`RANDOM}};
  valid_929 = _RAND_945[0:0];
  _RAND_946 = {1{`RANDOM}};
  valid_930 = _RAND_946[0:0];
  _RAND_947 = {1{`RANDOM}};
  valid_931 = _RAND_947[0:0];
  _RAND_948 = {1{`RANDOM}};
  valid_932 = _RAND_948[0:0];
  _RAND_949 = {1{`RANDOM}};
  valid_933 = _RAND_949[0:0];
  _RAND_950 = {1{`RANDOM}};
  valid_934 = _RAND_950[0:0];
  _RAND_951 = {1{`RANDOM}};
  valid_935 = _RAND_951[0:0];
  _RAND_952 = {1{`RANDOM}};
  valid_936 = _RAND_952[0:0];
  _RAND_953 = {1{`RANDOM}};
  valid_937 = _RAND_953[0:0];
  _RAND_954 = {1{`RANDOM}};
  valid_938 = _RAND_954[0:0];
  _RAND_955 = {1{`RANDOM}};
  valid_939 = _RAND_955[0:0];
  _RAND_956 = {1{`RANDOM}};
  valid_940 = _RAND_956[0:0];
  _RAND_957 = {1{`RANDOM}};
  valid_941 = _RAND_957[0:0];
  _RAND_958 = {1{`RANDOM}};
  valid_942 = _RAND_958[0:0];
  _RAND_959 = {1{`RANDOM}};
  valid_943 = _RAND_959[0:0];
  _RAND_960 = {1{`RANDOM}};
  valid_944 = _RAND_960[0:0];
  _RAND_961 = {1{`RANDOM}};
  valid_945 = _RAND_961[0:0];
  _RAND_962 = {1{`RANDOM}};
  valid_946 = _RAND_962[0:0];
  _RAND_963 = {1{`RANDOM}};
  valid_947 = _RAND_963[0:0];
  _RAND_964 = {1{`RANDOM}};
  valid_948 = _RAND_964[0:0];
  _RAND_965 = {1{`RANDOM}};
  valid_949 = _RAND_965[0:0];
  _RAND_966 = {1{`RANDOM}};
  valid_950 = _RAND_966[0:0];
  _RAND_967 = {1{`RANDOM}};
  valid_951 = _RAND_967[0:0];
  _RAND_968 = {1{`RANDOM}};
  valid_952 = _RAND_968[0:0];
  _RAND_969 = {1{`RANDOM}};
  valid_953 = _RAND_969[0:0];
  _RAND_970 = {1{`RANDOM}};
  valid_954 = _RAND_970[0:0];
  _RAND_971 = {1{`RANDOM}};
  valid_955 = _RAND_971[0:0];
  _RAND_972 = {1{`RANDOM}};
  valid_956 = _RAND_972[0:0];
  _RAND_973 = {1{`RANDOM}};
  valid_957 = _RAND_973[0:0];
  _RAND_974 = {1{`RANDOM}};
  valid_958 = _RAND_974[0:0];
  _RAND_975 = {1{`RANDOM}};
  valid_959 = _RAND_975[0:0];
  _RAND_976 = {1{`RANDOM}};
  valid_960 = _RAND_976[0:0];
  _RAND_977 = {1{`RANDOM}};
  valid_961 = _RAND_977[0:0];
  _RAND_978 = {1{`RANDOM}};
  valid_962 = _RAND_978[0:0];
  _RAND_979 = {1{`RANDOM}};
  valid_963 = _RAND_979[0:0];
  _RAND_980 = {1{`RANDOM}};
  valid_964 = _RAND_980[0:0];
  _RAND_981 = {1{`RANDOM}};
  valid_965 = _RAND_981[0:0];
  _RAND_982 = {1{`RANDOM}};
  valid_966 = _RAND_982[0:0];
  _RAND_983 = {1{`RANDOM}};
  valid_967 = _RAND_983[0:0];
  _RAND_984 = {1{`RANDOM}};
  valid_968 = _RAND_984[0:0];
  _RAND_985 = {1{`RANDOM}};
  valid_969 = _RAND_985[0:0];
  _RAND_986 = {1{`RANDOM}};
  valid_970 = _RAND_986[0:0];
  _RAND_987 = {1{`RANDOM}};
  valid_971 = _RAND_987[0:0];
  _RAND_988 = {1{`RANDOM}};
  valid_972 = _RAND_988[0:0];
  _RAND_989 = {1{`RANDOM}};
  valid_973 = _RAND_989[0:0];
  _RAND_990 = {1{`RANDOM}};
  valid_974 = _RAND_990[0:0];
  _RAND_991 = {1{`RANDOM}};
  valid_975 = _RAND_991[0:0];
  _RAND_992 = {1{`RANDOM}};
  valid_976 = _RAND_992[0:0];
  _RAND_993 = {1{`RANDOM}};
  valid_977 = _RAND_993[0:0];
  _RAND_994 = {1{`RANDOM}};
  valid_978 = _RAND_994[0:0];
  _RAND_995 = {1{`RANDOM}};
  valid_979 = _RAND_995[0:0];
  _RAND_996 = {1{`RANDOM}};
  valid_980 = _RAND_996[0:0];
  _RAND_997 = {1{`RANDOM}};
  valid_981 = _RAND_997[0:0];
  _RAND_998 = {1{`RANDOM}};
  valid_982 = _RAND_998[0:0];
  _RAND_999 = {1{`RANDOM}};
  valid_983 = _RAND_999[0:0];
  _RAND_1000 = {1{`RANDOM}};
  valid_984 = _RAND_1000[0:0];
  _RAND_1001 = {1{`RANDOM}};
  valid_985 = _RAND_1001[0:0];
  _RAND_1002 = {1{`RANDOM}};
  valid_986 = _RAND_1002[0:0];
  _RAND_1003 = {1{`RANDOM}};
  valid_987 = _RAND_1003[0:0];
  _RAND_1004 = {1{`RANDOM}};
  valid_988 = _RAND_1004[0:0];
  _RAND_1005 = {1{`RANDOM}};
  valid_989 = _RAND_1005[0:0];
  _RAND_1006 = {1{`RANDOM}};
  valid_990 = _RAND_1006[0:0];
  _RAND_1007 = {1{`RANDOM}};
  valid_991 = _RAND_1007[0:0];
  _RAND_1008 = {1{`RANDOM}};
  valid_992 = _RAND_1008[0:0];
  _RAND_1009 = {1{`RANDOM}};
  valid_993 = _RAND_1009[0:0];
  _RAND_1010 = {1{`RANDOM}};
  valid_994 = _RAND_1010[0:0];
  _RAND_1011 = {1{`RANDOM}};
  valid_995 = _RAND_1011[0:0];
  _RAND_1012 = {1{`RANDOM}};
  valid_996 = _RAND_1012[0:0];
  _RAND_1013 = {1{`RANDOM}};
  valid_997 = _RAND_1013[0:0];
  _RAND_1014 = {1{`RANDOM}};
  valid_998 = _RAND_1014[0:0];
  _RAND_1015 = {1{`RANDOM}};
  valid_999 = _RAND_1015[0:0];
  _RAND_1016 = {1{`RANDOM}};
  valid_1000 = _RAND_1016[0:0];
  _RAND_1017 = {1{`RANDOM}};
  valid_1001 = _RAND_1017[0:0];
  _RAND_1018 = {1{`RANDOM}};
  valid_1002 = _RAND_1018[0:0];
  _RAND_1019 = {1{`RANDOM}};
  valid_1003 = _RAND_1019[0:0];
  _RAND_1020 = {1{`RANDOM}};
  valid_1004 = _RAND_1020[0:0];
  _RAND_1021 = {1{`RANDOM}};
  valid_1005 = _RAND_1021[0:0];
  _RAND_1022 = {1{`RANDOM}};
  valid_1006 = _RAND_1022[0:0];
  _RAND_1023 = {1{`RANDOM}};
  valid_1007 = _RAND_1023[0:0];
  _RAND_1024 = {1{`RANDOM}};
  valid_1008 = _RAND_1024[0:0];
  _RAND_1025 = {1{`RANDOM}};
  valid_1009 = _RAND_1025[0:0];
  _RAND_1026 = {1{`RANDOM}};
  valid_1010 = _RAND_1026[0:0];
  _RAND_1027 = {1{`RANDOM}};
  valid_1011 = _RAND_1027[0:0];
  _RAND_1028 = {1{`RANDOM}};
  valid_1012 = _RAND_1028[0:0];
  _RAND_1029 = {1{`RANDOM}};
  valid_1013 = _RAND_1029[0:0];
  _RAND_1030 = {1{`RANDOM}};
  valid_1014 = _RAND_1030[0:0];
  _RAND_1031 = {1{`RANDOM}};
  valid_1015 = _RAND_1031[0:0];
  _RAND_1032 = {1{`RANDOM}};
  valid_1016 = _RAND_1032[0:0];
  _RAND_1033 = {1{`RANDOM}};
  valid_1017 = _RAND_1033[0:0];
  _RAND_1034 = {1{`RANDOM}};
  valid_1018 = _RAND_1034[0:0];
  _RAND_1035 = {1{`RANDOM}};
  valid_1019 = _RAND_1035[0:0];
  _RAND_1036 = {1{`RANDOM}};
  valid_1020 = _RAND_1036[0:0];
  _RAND_1037 = {1{`RANDOM}};
  valid_1021 = _RAND_1037[0:0];
  _RAND_1038 = {1{`RANDOM}};
  valid_1022 = _RAND_1038[0:0];
  _RAND_1039 = {1{`RANDOM}};
  valid_1023 = _RAND_1039[0:0];
  _RAND_1040 = {1{`RANDOM}};
  array_out_REG = _RAND_1040[0:0];
  _RAND_1041 = {9{`RANDOM}};
  array_out_r = _RAND_1041[272:0];
  _RAND_1042 = {1{`RANDOM}};
  lrsc_addr = _RAND_1042[26:0];
  _RAND_1043 = {1{`RANDOM}};
  sc_fail_r = _RAND_1043[0:0];
  _RAND_1044 = {1{`RANDOM}};
  probe_out_REG = _RAND_1044[0:0];
  _RAND_1045 = {9{`RANDOM}};
  probe_out_r = _RAND_1045[272:0];
  _RAND_1046 = {1{`RANDOM}};
  release_addr_aligned_REG = _RAND_1046[9:0];
  _RAND_1047 = {1{`RANDOM}};
  source = _RAND_1047[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Uncache(
  input         clock,
  input         reset,
  input         auto_out_a_ready,
  output        auto_out_a_valid,
  output [2:0]  auto_out_a_bits_opcode,
  output [2:0]  auto_out_a_bits_size,
  output [1:0]  auto_out_a_bits_source,
  output [31:0] auto_out_a_bits_address,
  output [7:0]  auto_out_a_bits_mask,
  output [63:0] auto_out_a_bits_data,
  output        auto_out_d_ready,
  input         auto_out_d_valid,
  input  [63:0] auto_out_d_bits_data,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [38:0] io_in_req_bits_addr,
  input  [63:0] io_in_req_bits_wdata,
  input  [7:0]  io_in_req_bits_wmask,
  input         io_in_req_bits_wen,
  input  [1:0]  io_in_req_bits_len,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [63:0] io_in_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  _source_T = auto_out_a_ready & io_in_req_valid; // @[Decoupled.scala 51:35]
  reg [1:0] source; // @[Counter.scala 61:40]
  wire [1:0] _source_wrap_value_T_1 = source + 2'h1; // @[Counter.scala 77:24]
  wire [2:0] _get_bits_a_mask_sizeOH_T = {{1'd0}, io_in_req_bits_len}; // @[Misc.scala 201:34]
  wire [1:0] get_bits_a_mask_sizeOH_shiftAmount = _get_bits_a_mask_sizeOH_T[1:0]; // @[OneHot.scala 63:49]
  wire [3:0] _get_bits_a_mask_sizeOH_T_1 = 4'h1 << get_bits_a_mask_sizeOH_shiftAmount; // @[OneHot.scala 64:12]
  wire [2:0] get_bits_a_mask_sizeOH = _get_bits_a_mask_sizeOH_T_1[2:0] | 3'h1; // @[Misc.scala 201:81]
  wire  _get_bits_a_mask_T = io_in_req_bits_len >= 2'h3; // @[Misc.scala 205:21]
  wire  get_bits_a_mask_size = get_bits_a_mask_sizeOH[2]; // @[Misc.scala 208:26]
  wire  get_bits_a_mask_bit = io_in_req_bits_addr[2]; // @[Misc.scala 209:26]
  wire  get_bits_a_mask_nbit = ~get_bits_a_mask_bit; // @[Misc.scala 210:20]
  wire  get_bits_a_mask_acc = _get_bits_a_mask_T | get_bits_a_mask_size & get_bits_a_mask_nbit; // @[Misc.scala 214:29]
  wire  get_bits_a_mask_acc_1 = _get_bits_a_mask_T | get_bits_a_mask_size & get_bits_a_mask_bit; // @[Misc.scala 214:29]
  wire  get_bits_a_mask_size_1 = get_bits_a_mask_sizeOH[1]; // @[Misc.scala 208:26]
  wire  get_bits_a_mask_bit_1 = io_in_req_bits_addr[1]; // @[Misc.scala 209:26]
  wire  get_bits_a_mask_nbit_1 = ~get_bits_a_mask_bit_1; // @[Misc.scala 210:20]
  wire  get_bits_a_mask_eq_2 = get_bits_a_mask_nbit & get_bits_a_mask_nbit_1; // @[Misc.scala 213:27]
  wire  get_bits_a_mask_acc_2 = get_bits_a_mask_acc | get_bits_a_mask_size_1 & get_bits_a_mask_eq_2; // @[Misc.scala 214:29]
  wire  get_bits_a_mask_eq_3 = get_bits_a_mask_nbit & get_bits_a_mask_bit_1; // @[Misc.scala 213:27]
  wire  get_bits_a_mask_acc_3 = get_bits_a_mask_acc | get_bits_a_mask_size_1 & get_bits_a_mask_eq_3; // @[Misc.scala 214:29]
  wire  get_bits_a_mask_eq_4 = get_bits_a_mask_bit & get_bits_a_mask_nbit_1; // @[Misc.scala 213:27]
  wire  get_bits_a_mask_acc_4 = get_bits_a_mask_acc_1 | get_bits_a_mask_size_1 & get_bits_a_mask_eq_4; // @[Misc.scala 214:29]
  wire  get_bits_a_mask_eq_5 = get_bits_a_mask_bit & get_bits_a_mask_bit_1; // @[Misc.scala 213:27]
  wire  get_bits_a_mask_acc_5 = get_bits_a_mask_acc_1 | get_bits_a_mask_size_1 & get_bits_a_mask_eq_5; // @[Misc.scala 214:29]
  wire  get_bits_a_mask_size_2 = get_bits_a_mask_sizeOH[0]; // @[Misc.scala 208:26]
  wire  get_bits_a_mask_bit_2 = io_in_req_bits_addr[0]; // @[Misc.scala 209:26]
  wire  get_bits_a_mask_nbit_2 = ~get_bits_a_mask_bit_2; // @[Misc.scala 210:20]
  wire  get_bits_a_mask_eq_6 = get_bits_a_mask_eq_2 & get_bits_a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  get_bits_a_mask_acc_6 = get_bits_a_mask_acc_2 | get_bits_a_mask_size_2 & get_bits_a_mask_eq_6; // @[Misc.scala 214:29]
  wire  get_bits_a_mask_eq_7 = get_bits_a_mask_eq_2 & get_bits_a_mask_bit_2; // @[Misc.scala 213:27]
  wire  get_bits_a_mask_acc_7 = get_bits_a_mask_acc_2 | get_bits_a_mask_size_2 & get_bits_a_mask_eq_7; // @[Misc.scala 214:29]
  wire  get_bits_a_mask_eq_8 = get_bits_a_mask_eq_3 & get_bits_a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  get_bits_a_mask_acc_8 = get_bits_a_mask_acc_3 | get_bits_a_mask_size_2 & get_bits_a_mask_eq_8; // @[Misc.scala 214:29]
  wire  get_bits_a_mask_eq_9 = get_bits_a_mask_eq_3 & get_bits_a_mask_bit_2; // @[Misc.scala 213:27]
  wire  get_bits_a_mask_acc_9 = get_bits_a_mask_acc_3 | get_bits_a_mask_size_2 & get_bits_a_mask_eq_9; // @[Misc.scala 214:29]
  wire  get_bits_a_mask_eq_10 = get_bits_a_mask_eq_4 & get_bits_a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  get_bits_a_mask_acc_10 = get_bits_a_mask_acc_4 | get_bits_a_mask_size_2 & get_bits_a_mask_eq_10; // @[Misc.scala 214:29]
  wire  get_bits_a_mask_eq_11 = get_bits_a_mask_eq_4 & get_bits_a_mask_bit_2; // @[Misc.scala 213:27]
  wire  get_bits_a_mask_acc_11 = get_bits_a_mask_acc_4 | get_bits_a_mask_size_2 & get_bits_a_mask_eq_11; // @[Misc.scala 214:29]
  wire  get_bits_a_mask_eq_12 = get_bits_a_mask_eq_5 & get_bits_a_mask_nbit_2; // @[Misc.scala 213:27]
  wire  get_bits_a_mask_acc_12 = get_bits_a_mask_acc_5 | get_bits_a_mask_size_2 & get_bits_a_mask_eq_12; // @[Misc.scala 214:29]
  wire  get_bits_a_mask_eq_13 = get_bits_a_mask_eq_5 & get_bits_a_mask_bit_2; // @[Misc.scala 213:27]
  wire  get_bits_a_mask_acc_13 = get_bits_a_mask_acc_5 | get_bits_a_mask_size_2 & get_bits_a_mask_eq_13; // @[Misc.scala 214:29]
  wire [7:0] get_bits_mask = {get_bits_a_mask_acc_13,get_bits_a_mask_acc_12,get_bits_a_mask_acc_11,
    get_bits_a_mask_acc_10,get_bits_a_mask_acc_9,get_bits_a_mask_acc_8,get_bits_a_mask_acc_7,get_bits_a_mask_acc_6}; // @[Cat.scala 33:92]
  wire [31:0] put_bits_address = io_in_req_bits_addr[31:0]; // @[Edges.scala 483:17 488:15]
  assign auto_out_a_valid = io_in_req_valid; // @[Nodes.scala 1212:84 Bus.scala 140:14]
  assign auto_out_a_bits_opcode = io_in_req_bits_wen ? 3'h1 : 3'h4; // @[Bus.scala 150:25]
  assign auto_out_a_bits_size = io_in_req_bits_wen ? _get_bits_a_mask_sizeOH_T : _get_bits_a_mask_sizeOH_T; // @[Bus.scala 150:25]
  assign auto_out_a_bits_source = source; // @[Bus.scala 150:25]
  assign auto_out_a_bits_address = io_in_req_bits_wen ? put_bits_address : put_bits_address; // @[Bus.scala 150:25]
  assign auto_out_a_bits_mask = io_in_req_bits_wen ? io_in_req_bits_wmask : get_bits_mask; // @[Bus.scala 150:25]
  assign auto_out_a_bits_data = io_in_req_bits_wen ? io_in_req_bits_wdata : 64'h0; // @[Bus.scala 150:25]
  assign auto_out_d_ready = io_in_resp_ready; // @[Nodes.scala 1212:84 Bus.scala 143:14]
  assign io_in_req_ready = auto_out_a_ready; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign io_in_resp_valid = auto_out_d_valid; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign io_in_resp_bits_rdata = auto_out_d_bits_data; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  always @(posedge clock) begin
    if (reset) begin // @[Counter.scala 61:40]
      source <= 2'h0; // @[Counter.scala 61:40]
    end else if (_source_T) begin // @[Counter.scala 118:16]
      source <= _source_wrap_value_T_1; // @[Counter.scala 77:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  source = _RAND_0[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLXbar(
  input          clock,
  input          reset,
  output         auto_in_2_a_ready,
  input          auto_in_2_a_valid,
  input  [1:0]   auto_in_2_a_bits_source,
  input  [31:0]  auto_in_2_a_bits_address,
  input          auto_in_2_b_ready,
  output         auto_in_2_b_valid,
  output [2:0]   auto_in_2_b_bits_size,
  output [1:0]   auto_in_2_b_bits_source,
  output [31:0]  auto_in_2_b_bits_address,
  output         auto_in_2_c_ready,
  input          auto_in_2_c_valid,
  input  [2:0]   auto_in_2_c_bits_opcode,
  input  [2:0]   auto_in_2_c_bits_param,
  input  [2:0]   auto_in_2_c_bits_size,
  input  [1:0]   auto_in_2_c_bits_source,
  input  [31:0]  auto_in_2_c_bits_address,
  input  [255:0] auto_in_2_c_bits_data,
  input          auto_in_2_d_ready,
  output         auto_in_2_d_valid,
  output [5:0]   auto_in_2_d_bits_sink,
  output [255:0] auto_in_2_d_bits_data,
  output         auto_in_2_e_ready,
  input          auto_in_2_e_valid,
  input  [5:0]   auto_in_2_e_bits_sink,
  output         auto_in_1_a_ready,
  input          auto_in_1_a_valid,
  input  [2:0]   auto_in_1_a_bits_opcode,
  input  [2:0]   auto_in_1_a_bits_size,
  input  [1:0]   auto_in_1_a_bits_source,
  input  [31:0]  auto_in_1_a_bits_address,
  input  [31:0]  auto_in_1_a_bits_mask,
  input  [255:0] auto_in_1_a_bits_data,
  input          auto_in_1_d_ready,
  output         auto_in_1_d_valid,
  output [2:0]   auto_in_1_d_bits_opcode,
  output [2:0]   auto_in_1_d_bits_size,
  output [1:0]   auto_in_1_d_bits_source,
  output [255:0] auto_in_1_d_bits_data,
  output         auto_in_0_a_ready,
  input          auto_in_0_a_valid,
  input  [1:0]   auto_in_0_a_bits_source,
  input  [31:0]  auto_in_0_a_bits_address,
  input          auto_in_0_d_ready,
  output         auto_in_0_d_valid,
  output [255:0] auto_in_0_d_bits_data,
  input          auto_out_a_ready,
  output         auto_out_a_valid,
  output [2:0]   auto_out_a_bits_opcode,
  output [2:0]   auto_out_a_bits_param,
  output [2:0]   auto_out_a_bits_size,
  output [3:0]   auto_out_a_bits_source,
  output [31:0]  auto_out_a_bits_address,
  output [31:0]  auto_out_a_bits_mask,
  output [255:0] auto_out_a_bits_data,
  output         auto_out_b_ready,
  input          auto_out_b_valid,
  input  [2:0]   auto_out_b_bits_size,
  input  [3:0]   auto_out_b_bits_source,
  input  [31:0]  auto_out_b_bits_address,
  input          auto_out_c_ready,
  output         auto_out_c_valid,
  output [2:0]   auto_out_c_bits_opcode,
  output [2:0]   auto_out_c_bits_param,
  output [2:0]   auto_out_c_bits_size,
  output [3:0]   auto_out_c_bits_source,
  output [31:0]  auto_out_c_bits_address,
  output [255:0] auto_out_c_bits_data,
  output         auto_out_d_ready,
  input          auto_out_d_valid,
  input  [2:0]   auto_out_d_bits_opcode,
  input  [2:0]   auto_out_d_bits_size,
  input  [3:0]   auto_out_d_bits_source,
  input  [5:0]   auto_out_d_bits_sink,
  input  [255:0] auto_out_d_bits_data,
  input          auto_out_e_ready,
  output         auto_out_e_valid,
  output [5:0]   auto_out_e_bits_sink
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire [3:0] _GEN_0 = {{2'd0}, auto_in_0_a_bits_source}; // @[Xbar.scala 240:55]
  wire [3:0] in_0_a_bits_source = _GEN_0 | 4'h8; // @[Xbar.scala 240:55]
  wire [2:0] _GEN_1 = {{1'd0}, auto_in_1_a_bits_source}; // @[Xbar.scala 240:55]
  wire [2:0] _in_1_a_bits_source_T = _GEN_1 | 3'h4; // @[Xbar.scala 240:55]
  wire  requestBOI_0_2 = auto_out_b_bits_source[3:2] == 2'h0; // @[Parameters.scala 54:32]
  wire  requestDOI_0_0 = auto_out_d_bits_source[3:2] == 2'h2; // @[Parameters.scala 54:32]
  wire  requestDOI_0_1 = auto_out_d_bits_source[3:2] == 2'h1; // @[Parameters.scala 54:32]
  wire  requestDOI_0_2 = auto_out_d_bits_source[3:2] == 2'h0; // @[Parameters.scala 54:32]
  reg  beatsLeft; // @[Arbiter.scala 88:30]
  wire  idle = ~beatsLeft; // @[Arbiter.scala 89:28]
  wire  latch = idle & auto_out_a_ready; // @[Arbiter.scala 90:24]
  wire [2:0] _readys_T = {auto_in_2_a_valid,auto_in_1_a_valid,auto_in_0_a_valid}; // @[Cat.scala 33:92]
  wire [2:0] _GEN_2 = {{1'd0}, _readys_T[2:1]}; // @[package.scala 254:43]
  wire [2:0] _readys_T_2 = _readys_T | _GEN_2; // @[package.scala 254:43]
  wire [2:0] _GEN_3 = {{2'd0}, _readys_T_2[2]}; // @[package.scala 254:43]
  wire [2:0] _readys_T_4 = _readys_T_2 | _GEN_3; // @[package.scala 254:43]
  wire [2:0] _readys_T_7 = {{1'd0}, _readys_T_4[2:1]}; // @[Arbiter.scala 19:90]
  wire [2:0] _readys_T_8 = ~_readys_T_7; // @[Arbiter.scala 19:62]
  wire  readys_0 = _readys_T_8[0]; // @[Arbiter.scala 96:86]
  wire  readys_1 = _readys_T_8[1]; // @[Arbiter.scala 96:86]
  wire  readys_2 = _readys_T_8[2]; // @[Arbiter.scala 96:86]
  wire  earlyWinner_0 = readys_0 & auto_in_0_a_valid; // @[Arbiter.scala 98:79]
  wire  earlyWinner_1 = readys_1 & auto_in_1_a_valid; // @[Arbiter.scala 98:79]
  wire  earlyWinner_2 = readys_2 & auto_in_2_a_valid; // @[Arbiter.scala 98:79]
  wire  prefixOR_2 = earlyWinner_0 | earlyWinner_1; // @[Arbiter.scala 105:53]
  wire  _prefixOR_T = prefixOR_2 | earlyWinner_2; // @[Arbiter.scala 105:53]
  wire  _T_13 = ~reset; // @[Arbiter.scala 106:13]
  wire  _T_16 = auto_in_0_a_valid | auto_in_1_a_valid | auto_in_2_a_valid; // @[Arbiter.scala 108:36]
  wire  _T_17 = ~(auto_in_0_a_valid | auto_in_1_a_valid | auto_in_2_a_valid); // @[Arbiter.scala 108:15]
  reg  state_0; // @[Arbiter.scala 117:26]
  wire  muxStateEarly_0 = idle ? earlyWinner_0 : state_0; // @[Arbiter.scala 118:30]
  reg  state_1; // @[Arbiter.scala 117:26]
  wire  muxStateEarly_1 = idle ? earlyWinner_1 : state_1; // @[Arbiter.scala 118:30]
  reg  state_2; // @[Arbiter.scala 117:26]
  wire  muxStateEarly_2 = idle ? earlyWinner_2 : state_2; // @[Arbiter.scala 118:30]
  wire  _out_0_a_earlyValid_T_6 = state_0 & auto_in_0_a_valid | state_1 & auto_in_1_a_valid | state_2 &
    auto_in_2_a_valid; // @[Mux.scala 27:73]
  wire  out_3_0_a_earlyValid = idle ? _T_16 : _out_0_a_earlyValid_T_6; // @[Arbiter.scala 126:29]
  wire  _beatsLeft_T_2 = auto_out_a_ready & out_3_0_a_earlyValid; // @[ReadyValidCancel.scala 49:33]
  wire  allowed_0 = idle ? readys_0 : state_0; // @[Arbiter.scala 122:24]
  wire  allowed_1 = idle ? readys_1 : state_1; // @[Arbiter.scala 122:24]
  wire  allowed_2 = idle ? readys_2 : state_2; // @[Arbiter.scala 122:24]
  wire [31:0] _T_43 = muxStateEarly_0 ? 32'hffffffff : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _T_44 = muxStateEarly_1 ? auto_in_1_a_bits_mask : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _T_45 = muxStateEarly_2 ? 32'hffffffff : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _T_46 = _T_43 | _T_44; // @[Mux.scala 27:73]
  wire [31:0] _T_48 = muxStateEarly_0 ? auto_in_0_a_bits_address : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _T_49 = muxStateEarly_1 ? auto_in_1_a_bits_address : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _T_50 = muxStateEarly_2 ? auto_in_2_a_bits_address : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _T_51 = _T_48 | _T_49; // @[Mux.scala 27:73]
  wire [3:0] _T_53 = muxStateEarly_0 ? in_0_a_bits_source : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] in_1_a_bits_source = {{1'd0}, _in_1_a_bits_source_T}; // @[Xbar.scala 234:18 240:29]
  wire [3:0] _T_54 = muxStateEarly_1 ? in_1_a_bits_source : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] in_2_a_bits_source = {{2'd0}, auto_in_2_a_bits_source}; // @[Xbar.scala 234:18 240:29]
  wire [3:0] _T_55 = muxStateEarly_2 ? in_2_a_bits_source : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _T_56 = _T_53 | _T_54; // @[Mux.scala 27:73]
  wire [2:0] _T_58 = muxStateEarly_0 ? 3'h5 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_59 = muxStateEarly_1 ? auto_in_1_a_bits_size : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_60 = muxStateEarly_2 ? 3'h5 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_61 = _T_58 | _T_59; // @[Mux.scala 27:73]
  wire [2:0] _T_68 = muxStateEarly_0 ? 3'h4 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_69 = muxStateEarly_1 ? auto_in_1_a_bits_opcode : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_70 = muxStateEarly_2 ? 3'h6 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_71 = _T_68 | _T_69; // @[Mux.scala 27:73]
  assign auto_in_2_a_ready = auto_out_a_ready & allowed_2; // @[Arbiter.scala 124:31]
  assign auto_in_2_b_valid = auto_out_b_valid & requestBOI_0_2; // @[Xbar.scala 182:40]
  assign auto_in_2_b_bits_size = auto_out_b_bits_size; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_2_b_bits_source = auto_out_b_bits_source[1:0]; // @[Xbar.scala 231:69]
  assign auto_in_2_b_bits_address = auto_out_b_bits_address; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_2_c_ready = auto_out_c_ready; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_2_d_valid = auto_out_d_valid & requestDOI_0_2; // @[Xbar.scala 182:40]
  assign auto_in_2_d_bits_sink = auto_out_d_bits_sink; // @[Xbar.scala 326:53]
  assign auto_in_2_d_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_2_e_ready = auto_out_e_ready; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_1_a_ready = auto_out_a_ready & allowed_1; // @[Arbiter.scala 124:31]
  assign auto_in_1_d_valid = auto_out_d_valid & requestDOI_0_1; // @[Xbar.scala 182:40]
  assign auto_in_1_d_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_1_d_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_1_d_bits_source = auto_out_d_bits_source[1:0]; // @[Xbar.scala 231:69]
  assign auto_in_1_d_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_in_0_a_ready = auto_out_a_ready & allowed_0; // @[Arbiter.scala 124:31]
  assign auto_in_0_d_valid = auto_out_d_valid & requestDOI_0_0; // @[Xbar.scala 182:40]
  assign auto_in_0_d_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign auto_out_a_valid = idle ? _T_16 : _out_0_a_earlyValid_T_6; // @[Arbiter.scala 126:29]
  assign auto_out_a_bits_opcode = _T_71 | _T_70; // @[Mux.scala 27:73]
  assign auto_out_a_bits_param = muxStateEarly_2 ? 3'h1 : 3'h0; // @[Mux.scala 27:73]
  assign auto_out_a_bits_size = _T_61 | _T_60; // @[Mux.scala 27:73]
  assign auto_out_a_bits_source = _T_56 | _T_55; // @[Mux.scala 27:73]
  assign auto_out_a_bits_address = _T_51 | _T_50; // @[Mux.scala 27:73]
  assign auto_out_a_bits_mask = _T_46 | _T_45; // @[Mux.scala 27:73]
  assign auto_out_a_bits_data = muxStateEarly_1 ? auto_in_1_a_bits_data : 256'h0; // @[Mux.scala 27:73]
  assign auto_out_b_ready = requestBOI_0_2 & auto_in_2_b_ready; // @[Mux.scala 27:73]
  assign auto_out_c_valid = auto_in_2_c_valid; // @[ReadyValidCancel.scala 21:38]
  assign auto_out_c_bits_opcode = auto_in_2_c_bits_opcode; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_c_bits_param = auto_in_2_c_bits_param; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_c_bits_size = auto_in_2_c_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_c_bits_source = {{2'd0}, auto_in_2_c_bits_source}; // @[Xbar.scala 234:18 262:29]
  assign auto_out_c_bits_address = auto_in_2_c_bits_address; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_c_bits_data = auto_in_2_c_bits_data; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_d_ready = requestDOI_0_0 & auto_in_0_d_ready | requestDOI_0_1 & auto_in_1_d_ready | requestDOI_0_2 &
    auto_in_2_d_ready; // @[Mux.scala 27:73]
  assign auto_out_e_valid = auto_in_2_e_valid; // @[ReadyValidCancel.scala 21:38]
  assign auto_out_e_bits_sink = auto_in_2_e_bits_sink; // @[Xbar.scala 231:69]
  always @(posedge clock) begin
    if (reset) begin // @[Arbiter.scala 88:30]
      beatsLeft <= 1'h0; // @[Arbiter.scala 88:30]
    end else if (latch) begin // @[Arbiter.scala 114:23]
      beatsLeft <= 1'h0;
    end else begin
      beatsLeft <= beatsLeft - _beatsLeft_T_2;
    end
    if (reset) begin // @[Arbiter.scala 117:26]
      state_0 <= 1'h0; // @[Arbiter.scala 117:26]
    end else if (idle) begin // @[Arbiter.scala 118:30]
      state_0 <= earlyWinner_0;
    end
    if (reset) begin // @[Arbiter.scala 117:26]
      state_1 <= 1'h0; // @[Arbiter.scala 117:26]
    end else if (idle) begin // @[Arbiter.scala 118:30]
      state_1 <= earlyWinner_1;
    end
    if (reset) begin // @[Arbiter.scala 117:26]
      state_2 <= 1'h0; // @[Arbiter.scala 117:26]
    end else if (idle) begin // @[Arbiter.scala 118:30]
      state_2 <= earlyWinner_2;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~((~earlyWinner_0 | ~earlyWinner_1) & (~prefixOR_2 | ~earlyWinner_2))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:106 assert((prefixOR zip earlyWinner) map { case (p,w) => !p || !w } reduce {_ && _})\n"
            ); // @[Arbiter.scala 106:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~((~earlyWinner_0 | ~earlyWinner_1) & (~prefixOR_2 | ~earlyWinner_2))) begin
          $fatal; // @[Arbiter.scala 106:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & ~(~(auto_in_0_a_valid | auto_in_1_a_valid | auto_in_2_a_valid) | _prefixOR_T)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:108 assert (!earlyValids.reduce(_||_) || earlyWinner.reduce(_||_))\n"
            ); // @[Arbiter.scala 108:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_13 & ~(~(auto_in_0_a_valid | auto_in_1_a_valid | auto_in_2_a_valid) | _prefixOR_T)) begin
          $fatal; // @[Arbiter.scala 108:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & ~(_T_17 | _T_16)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Arbiter.scala:109 assert (!validQuals .reduce(_||_) || validQuals .reduce(_||_))\n"
            ); // @[Arbiter.scala 109:14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_13 & ~(_T_17 | _T_16)) begin
          $fatal; // @[Arbiter.scala 109:14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  beatsLeft = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  state_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  state_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  state_2 = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Repeater(
  input          clock,
  input          reset,
  input          io_repeat,
  output         io_enq_ready,
  input          io_enq_valid,
  input  [2:0]   io_enq_bits_opcode,
  input  [2:0]   io_enq_bits_size,
  input  [1:0]   io_enq_bits_source,
  input  [255:0] io_enq_bits_data,
  input          io_deq_ready,
  output         io_deq_valid,
  output [2:0]   io_deq_bits_opcode,
  output [2:0]   io_deq_bits_size,
  output [1:0]   io_deq_bits_source,
  output [255:0] io_deq_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [255:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg  full; // @[Repeater.scala 19:21]
  reg [2:0] saved_opcode; // @[Repeater.scala 20:18]
  reg [2:0] saved_size; // @[Repeater.scala 20:18]
  reg [1:0] saved_source; // @[Repeater.scala 20:18]
  reg [255:0] saved_data; // @[Repeater.scala 20:18]
  wire  _T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  _GEN_0 = _T & io_repeat | full; // @[Repeater.scala 19:21 28:{38,45}]
  wire  _T_2 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  assign io_enq_ready = io_deq_ready & ~full; // @[Repeater.scala 24:32]
  assign io_deq_valid = io_enq_valid | full; // @[Repeater.scala 23:32]
  assign io_deq_bits_opcode = full ? saved_opcode : io_enq_bits_opcode; // @[Repeater.scala 25:21]
  assign io_deq_bits_size = full ? saved_size : io_enq_bits_size; // @[Repeater.scala 25:21]
  assign io_deq_bits_source = full ? saved_source : io_enq_bits_source; // @[Repeater.scala 25:21]
  assign io_deq_bits_data = full ? saved_data : io_enq_bits_data; // @[Repeater.scala 25:21]
  always @(posedge clock) begin
    if (reset) begin // @[Repeater.scala 19:21]
      full <= 1'h0; // @[Repeater.scala 19:21]
    end else if (_T_2 & ~io_repeat) begin // @[Repeater.scala 29:38]
      full <= 1'h0; // @[Repeater.scala 29:45]
    end else begin
      full <= _GEN_0;
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_opcode <= io_enq_bits_opcode; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_size <= io_enq_bits_size; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_source <= io_enq_bits_source; // @[Repeater.scala 28:62]
    end
    if (_T & io_repeat) begin // @[Repeater.scala 28:38]
      saved_data <= io_enq_bits_data; // @[Repeater.scala 28:62]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  full = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  saved_opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  saved_size = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  saved_source = _RAND_3[1:0];
  _RAND_4 = {8{`RANDOM}};
  saved_data = _RAND_4[255:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLWidthWidget(
  input          clock,
  input          reset,
  output         auto_in_a_ready,
  input          auto_in_a_valid,
  input  [2:0]   auto_in_a_bits_opcode,
  input  [2:0]   auto_in_a_bits_size,
  input  [1:0]   auto_in_a_bits_source,
  input  [31:0]  auto_in_a_bits_address,
  input  [7:0]   auto_in_a_bits_mask,
  input  [63:0]  auto_in_a_bits_data,
  input          auto_in_d_ready,
  output         auto_in_d_valid,
  output [63:0]  auto_in_d_bits_data,
  input          auto_out_a_ready,
  output         auto_out_a_valid,
  output [2:0]   auto_out_a_bits_opcode,
  output [2:0]   auto_out_a_bits_size,
  output [1:0]   auto_out_a_bits_source,
  output [31:0]  auto_out_a_bits_address,
  output [31:0]  auto_out_a_bits_mask,
  output [255:0] auto_out_a_bits_data,
  output         auto_out_d_ready,
  input          auto_out_d_valid,
  input  [2:0]   auto_out_d_bits_opcode,
  input  [2:0]   auto_out_d_bits_size,
  input  [1:0]   auto_out_d_bits_source,
  input  [255:0] auto_out_d_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
`endif // RANDOMIZE_REG_INIT
  wire  repeated_repeater_clock; // @[Repeater.scala 35:26]
  wire  repeated_repeater_reset; // @[Repeater.scala 35:26]
  wire  repeated_repeater_io_repeat; // @[Repeater.scala 35:26]
  wire  repeated_repeater_io_enq_ready; // @[Repeater.scala 35:26]
  wire  repeated_repeater_io_enq_valid; // @[Repeater.scala 35:26]
  wire [2:0] repeated_repeater_io_enq_bits_opcode; // @[Repeater.scala 35:26]
  wire [2:0] repeated_repeater_io_enq_bits_size; // @[Repeater.scala 35:26]
  wire [1:0] repeated_repeater_io_enq_bits_source; // @[Repeater.scala 35:26]
  wire [255:0] repeated_repeater_io_enq_bits_data; // @[Repeater.scala 35:26]
  wire  repeated_repeater_io_deq_ready; // @[Repeater.scala 35:26]
  wire  repeated_repeater_io_deq_valid; // @[Repeater.scala 35:26]
  wire [2:0] repeated_repeater_io_deq_bits_opcode; // @[Repeater.scala 35:26]
  wire [2:0] repeated_repeater_io_deq_bits_size; // @[Repeater.scala 35:26]
  wire [1:0] repeated_repeater_io_deq_bits_source; // @[Repeater.scala 35:26]
  wire [255:0] repeated_repeater_io_deq_bits_data; // @[Repeater.scala 35:26]
  wire  hasData = ~auto_in_a_bits_opcode[2]; // @[Edges.scala 91:28]
  wire [11:0] _limit_T_1 = 12'h1f << auto_in_a_bits_size; // @[package.scala 235:71]
  wire [4:0] _limit_T_3 = ~_limit_T_1[4:0]; // @[package.scala 235:46]
  wire [1:0] limit = _limit_T_3[4:3]; // @[WidthWidget.scala 33:47]
  reg [1:0] count; // @[WidthWidget.scala 35:27]
  wire  last = count == limit | ~hasData; // @[WidthWidget.scala 37:36]
  wire [1:0] _enable_T_1 = count & limit; // @[WidthWidget.scala 38:63]
  wire  enable_0 = ~(|_enable_T_1); // @[WidthWidget.scala 38:47]
  wire [1:0] _enable_T_3 = count ^ 2'h1; // @[WidthWidget.scala 38:56]
  wire [1:0] _enable_T_4 = _enable_T_3 & limit; // @[WidthWidget.scala 38:63]
  wire  enable_1 = ~(|_enable_T_4); // @[WidthWidget.scala 38:47]
  wire [1:0] _enable_T_6 = count ^ 2'h2; // @[WidthWidget.scala 38:56]
  wire [1:0] _enable_T_7 = _enable_T_6 & limit; // @[WidthWidget.scala 38:63]
  wire  enable_2 = ~(|_enable_T_7); // @[WidthWidget.scala 38:47]
  wire  _bundleIn_0_a_ready_T = ~last; // @[WidthWidget.scala 71:32]
  wire  bundleIn_0_a_ready = auto_out_a_ready | ~last; // @[WidthWidget.scala 71:29]
  wire  _T = bundleIn_0_a_ready & auto_in_a_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _count_T_1 = count + 2'h1; // @[WidthWidget.scala 45:24]
  reg  x1_a_bits_data_rdata_written_once; // @[WidthWidget.scala 57:41]
  wire  x1_a_bits_data_masked_enable_0 = enable_0 | ~x1_a_bits_data_rdata_written_once; // @[WidthWidget.scala 58:42]
  wire  x1_a_bits_data_masked_enable_1 = enable_1 | ~x1_a_bits_data_rdata_written_once; // @[WidthWidget.scala 58:42]
  wire  x1_a_bits_data_masked_enable_2 = enable_2 | ~x1_a_bits_data_rdata_written_once; // @[WidthWidget.scala 58:42]
  reg [63:0] x1_a_bits_data_rdata_0; // @[WidthWidget.scala 61:24]
  reg [63:0] x1_a_bits_data_rdata_1; // @[WidthWidget.scala 61:24]
  reg [63:0] x1_a_bits_data_rdata_2; // @[WidthWidget.scala 61:24]
  wire [63:0] x1_a_bits_data_mdata_0 = x1_a_bits_data_masked_enable_0 ? auto_in_a_bits_data : x1_a_bits_data_rdata_0; // @[WidthWidget.scala 63:88]
  wire [63:0] x1_a_bits_data_mdata_1 = x1_a_bits_data_masked_enable_1 ? auto_in_a_bits_data : x1_a_bits_data_rdata_1; // @[WidthWidget.scala 63:88]
  wire [63:0] x1_a_bits_data_mdata_2 = x1_a_bits_data_masked_enable_2 ? auto_in_a_bits_data : x1_a_bits_data_rdata_2; // @[WidthWidget.scala 63:88]
  wire  _GEN_4 = _T & _bundleIn_0_a_ready_T | x1_a_bits_data_rdata_written_once; // @[WidthWidget.scala 64:35 65:30 57:41]
  wire [127:0] x1_a_bits_data_lo = {x1_a_bits_data_mdata_1,x1_a_bits_data_mdata_0}; // @[Cat.scala 33:92]
  wire [127:0] x1_a_bits_data_hi = {auto_in_a_bits_data,x1_a_bits_data_mdata_2}; // @[Cat.scala 33:92]
  wire [4:0] _x1_a_bits_mask_sizeOH_T = {{2'd0}, auto_in_a_bits_size}; // @[Misc.scala 201:34]
  wire [2:0] x1_a_bits_mask_sizeOH_shiftAmount = _x1_a_bits_mask_sizeOH_T[2:0]; // @[OneHot.scala 63:49]
  wire [7:0] _x1_a_bits_mask_sizeOH_T_1 = 8'h1 << x1_a_bits_mask_sizeOH_shiftAmount; // @[OneHot.scala 64:12]
  wire [4:0] x1_a_bits_mask_sizeOH = _x1_a_bits_mask_sizeOH_T_1[4:0] | 5'h1; // @[Misc.scala 201:81]
  wire  _x1_a_bits_mask_T = auto_in_a_bits_size >= 3'h5; // @[Misc.scala 205:21]
  wire  x1_a_bits_mask_size = x1_a_bits_mask_sizeOH[4]; // @[Misc.scala 208:26]
  wire  x1_a_bits_mask_bit = auto_in_a_bits_address[4]; // @[Misc.scala 209:26]
  wire  x1_a_bits_mask_nbit = ~x1_a_bits_mask_bit; // @[Misc.scala 210:20]
  wire  x1_a_bits_mask_acc = _x1_a_bits_mask_T | x1_a_bits_mask_size & x1_a_bits_mask_nbit; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_acc_1 = _x1_a_bits_mask_T | x1_a_bits_mask_size & x1_a_bits_mask_bit; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_size_1 = x1_a_bits_mask_sizeOH[3]; // @[Misc.scala 208:26]
  wire  x1_a_bits_mask_bit_1 = auto_in_a_bits_address[3]; // @[Misc.scala 209:26]
  wire  x1_a_bits_mask_nbit_1 = ~x1_a_bits_mask_bit_1; // @[Misc.scala 210:20]
  wire  x1_a_bits_mask_eq_2 = x1_a_bits_mask_nbit & x1_a_bits_mask_nbit_1; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_2 = x1_a_bits_mask_acc | x1_a_bits_mask_size_1 & x1_a_bits_mask_eq_2; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_3 = x1_a_bits_mask_nbit & x1_a_bits_mask_bit_1; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_3 = x1_a_bits_mask_acc | x1_a_bits_mask_size_1 & x1_a_bits_mask_eq_3; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_4 = x1_a_bits_mask_bit & x1_a_bits_mask_nbit_1; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_4 = x1_a_bits_mask_acc_1 | x1_a_bits_mask_size_1 & x1_a_bits_mask_eq_4; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_5 = x1_a_bits_mask_bit & x1_a_bits_mask_bit_1; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_5 = x1_a_bits_mask_acc_1 | x1_a_bits_mask_size_1 & x1_a_bits_mask_eq_5; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_size_2 = x1_a_bits_mask_sizeOH[2]; // @[Misc.scala 208:26]
  wire  x1_a_bits_mask_bit_2 = auto_in_a_bits_address[2]; // @[Misc.scala 209:26]
  wire  x1_a_bits_mask_nbit_2 = ~x1_a_bits_mask_bit_2; // @[Misc.scala 210:20]
  wire  x1_a_bits_mask_eq_6 = x1_a_bits_mask_eq_2 & x1_a_bits_mask_nbit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_6 = x1_a_bits_mask_acc_2 | x1_a_bits_mask_size_2 & x1_a_bits_mask_eq_6; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_7 = x1_a_bits_mask_eq_2 & x1_a_bits_mask_bit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_7 = x1_a_bits_mask_acc_2 | x1_a_bits_mask_size_2 & x1_a_bits_mask_eq_7; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_8 = x1_a_bits_mask_eq_3 & x1_a_bits_mask_nbit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_8 = x1_a_bits_mask_acc_3 | x1_a_bits_mask_size_2 & x1_a_bits_mask_eq_8; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_9 = x1_a_bits_mask_eq_3 & x1_a_bits_mask_bit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_9 = x1_a_bits_mask_acc_3 | x1_a_bits_mask_size_2 & x1_a_bits_mask_eq_9; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_10 = x1_a_bits_mask_eq_4 & x1_a_bits_mask_nbit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_10 = x1_a_bits_mask_acc_4 | x1_a_bits_mask_size_2 & x1_a_bits_mask_eq_10; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_11 = x1_a_bits_mask_eq_4 & x1_a_bits_mask_bit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_11 = x1_a_bits_mask_acc_4 | x1_a_bits_mask_size_2 & x1_a_bits_mask_eq_11; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_12 = x1_a_bits_mask_eq_5 & x1_a_bits_mask_nbit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_12 = x1_a_bits_mask_acc_5 | x1_a_bits_mask_size_2 & x1_a_bits_mask_eq_12; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_13 = x1_a_bits_mask_eq_5 & x1_a_bits_mask_bit_2; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_13 = x1_a_bits_mask_acc_5 | x1_a_bits_mask_size_2 & x1_a_bits_mask_eq_13; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_size_3 = x1_a_bits_mask_sizeOH[1]; // @[Misc.scala 208:26]
  wire  x1_a_bits_mask_bit_3 = auto_in_a_bits_address[1]; // @[Misc.scala 209:26]
  wire  x1_a_bits_mask_nbit_3 = ~x1_a_bits_mask_bit_3; // @[Misc.scala 210:20]
  wire  x1_a_bits_mask_eq_14 = x1_a_bits_mask_eq_6 & x1_a_bits_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_14 = x1_a_bits_mask_acc_6 | x1_a_bits_mask_size_3 & x1_a_bits_mask_eq_14; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_15 = x1_a_bits_mask_eq_6 & x1_a_bits_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_15 = x1_a_bits_mask_acc_6 | x1_a_bits_mask_size_3 & x1_a_bits_mask_eq_15; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_16 = x1_a_bits_mask_eq_7 & x1_a_bits_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_16 = x1_a_bits_mask_acc_7 | x1_a_bits_mask_size_3 & x1_a_bits_mask_eq_16; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_17 = x1_a_bits_mask_eq_7 & x1_a_bits_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_17 = x1_a_bits_mask_acc_7 | x1_a_bits_mask_size_3 & x1_a_bits_mask_eq_17; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_18 = x1_a_bits_mask_eq_8 & x1_a_bits_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_18 = x1_a_bits_mask_acc_8 | x1_a_bits_mask_size_3 & x1_a_bits_mask_eq_18; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_19 = x1_a_bits_mask_eq_8 & x1_a_bits_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_19 = x1_a_bits_mask_acc_8 | x1_a_bits_mask_size_3 & x1_a_bits_mask_eq_19; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_20 = x1_a_bits_mask_eq_9 & x1_a_bits_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_20 = x1_a_bits_mask_acc_9 | x1_a_bits_mask_size_3 & x1_a_bits_mask_eq_20; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_21 = x1_a_bits_mask_eq_9 & x1_a_bits_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_21 = x1_a_bits_mask_acc_9 | x1_a_bits_mask_size_3 & x1_a_bits_mask_eq_21; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_22 = x1_a_bits_mask_eq_10 & x1_a_bits_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_22 = x1_a_bits_mask_acc_10 | x1_a_bits_mask_size_3 & x1_a_bits_mask_eq_22; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_23 = x1_a_bits_mask_eq_10 & x1_a_bits_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_23 = x1_a_bits_mask_acc_10 | x1_a_bits_mask_size_3 & x1_a_bits_mask_eq_23; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_24 = x1_a_bits_mask_eq_11 & x1_a_bits_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_24 = x1_a_bits_mask_acc_11 | x1_a_bits_mask_size_3 & x1_a_bits_mask_eq_24; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_25 = x1_a_bits_mask_eq_11 & x1_a_bits_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_25 = x1_a_bits_mask_acc_11 | x1_a_bits_mask_size_3 & x1_a_bits_mask_eq_25; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_26 = x1_a_bits_mask_eq_12 & x1_a_bits_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_26 = x1_a_bits_mask_acc_12 | x1_a_bits_mask_size_3 & x1_a_bits_mask_eq_26; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_27 = x1_a_bits_mask_eq_12 & x1_a_bits_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_27 = x1_a_bits_mask_acc_12 | x1_a_bits_mask_size_3 & x1_a_bits_mask_eq_27; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_28 = x1_a_bits_mask_eq_13 & x1_a_bits_mask_nbit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_28 = x1_a_bits_mask_acc_13 | x1_a_bits_mask_size_3 & x1_a_bits_mask_eq_28; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_29 = x1_a_bits_mask_eq_13 & x1_a_bits_mask_bit_3; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_29 = x1_a_bits_mask_acc_13 | x1_a_bits_mask_size_3 & x1_a_bits_mask_eq_29; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_size_4 = x1_a_bits_mask_sizeOH[0]; // @[Misc.scala 208:26]
  wire  x1_a_bits_mask_bit_4 = auto_in_a_bits_address[0]; // @[Misc.scala 209:26]
  wire  x1_a_bits_mask_nbit_4 = ~x1_a_bits_mask_bit_4; // @[Misc.scala 210:20]
  wire  x1_a_bits_mask_eq_30 = x1_a_bits_mask_eq_14 & x1_a_bits_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_30 = x1_a_bits_mask_acc_14 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_30; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_31 = x1_a_bits_mask_eq_14 & x1_a_bits_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_31 = x1_a_bits_mask_acc_14 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_31; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_32 = x1_a_bits_mask_eq_15 & x1_a_bits_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_32 = x1_a_bits_mask_acc_15 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_32; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_33 = x1_a_bits_mask_eq_15 & x1_a_bits_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_33 = x1_a_bits_mask_acc_15 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_33; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_34 = x1_a_bits_mask_eq_16 & x1_a_bits_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_34 = x1_a_bits_mask_acc_16 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_34; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_35 = x1_a_bits_mask_eq_16 & x1_a_bits_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_35 = x1_a_bits_mask_acc_16 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_35; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_36 = x1_a_bits_mask_eq_17 & x1_a_bits_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_36 = x1_a_bits_mask_acc_17 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_36; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_37 = x1_a_bits_mask_eq_17 & x1_a_bits_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_37 = x1_a_bits_mask_acc_17 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_37; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_38 = x1_a_bits_mask_eq_18 & x1_a_bits_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_38 = x1_a_bits_mask_acc_18 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_38; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_39 = x1_a_bits_mask_eq_18 & x1_a_bits_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_39 = x1_a_bits_mask_acc_18 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_39; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_40 = x1_a_bits_mask_eq_19 & x1_a_bits_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_40 = x1_a_bits_mask_acc_19 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_40; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_41 = x1_a_bits_mask_eq_19 & x1_a_bits_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_41 = x1_a_bits_mask_acc_19 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_41; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_42 = x1_a_bits_mask_eq_20 & x1_a_bits_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_42 = x1_a_bits_mask_acc_20 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_42; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_43 = x1_a_bits_mask_eq_20 & x1_a_bits_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_43 = x1_a_bits_mask_acc_20 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_43; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_44 = x1_a_bits_mask_eq_21 & x1_a_bits_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_44 = x1_a_bits_mask_acc_21 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_44; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_45 = x1_a_bits_mask_eq_21 & x1_a_bits_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_45 = x1_a_bits_mask_acc_21 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_45; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_46 = x1_a_bits_mask_eq_22 & x1_a_bits_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_46 = x1_a_bits_mask_acc_22 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_46; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_47 = x1_a_bits_mask_eq_22 & x1_a_bits_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_47 = x1_a_bits_mask_acc_22 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_47; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_48 = x1_a_bits_mask_eq_23 & x1_a_bits_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_48 = x1_a_bits_mask_acc_23 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_48; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_49 = x1_a_bits_mask_eq_23 & x1_a_bits_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_49 = x1_a_bits_mask_acc_23 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_49; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_50 = x1_a_bits_mask_eq_24 & x1_a_bits_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_50 = x1_a_bits_mask_acc_24 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_50; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_51 = x1_a_bits_mask_eq_24 & x1_a_bits_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_51 = x1_a_bits_mask_acc_24 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_51; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_52 = x1_a_bits_mask_eq_25 & x1_a_bits_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_52 = x1_a_bits_mask_acc_25 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_52; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_53 = x1_a_bits_mask_eq_25 & x1_a_bits_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_53 = x1_a_bits_mask_acc_25 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_53; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_54 = x1_a_bits_mask_eq_26 & x1_a_bits_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_54 = x1_a_bits_mask_acc_26 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_54; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_55 = x1_a_bits_mask_eq_26 & x1_a_bits_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_55 = x1_a_bits_mask_acc_26 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_55; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_56 = x1_a_bits_mask_eq_27 & x1_a_bits_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_56 = x1_a_bits_mask_acc_27 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_56; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_57 = x1_a_bits_mask_eq_27 & x1_a_bits_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_57 = x1_a_bits_mask_acc_27 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_57; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_58 = x1_a_bits_mask_eq_28 & x1_a_bits_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_58 = x1_a_bits_mask_acc_28 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_58; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_59 = x1_a_bits_mask_eq_28 & x1_a_bits_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_59 = x1_a_bits_mask_acc_28 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_59; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_60 = x1_a_bits_mask_eq_29 & x1_a_bits_mask_nbit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_60 = x1_a_bits_mask_acc_29 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_60; // @[Misc.scala 214:29]
  wire  x1_a_bits_mask_eq_61 = x1_a_bits_mask_eq_29 & x1_a_bits_mask_bit_4; // @[Misc.scala 213:27]
  wire  x1_a_bits_mask_acc_61 = x1_a_bits_mask_acc_29 | x1_a_bits_mask_size_4 & x1_a_bits_mask_eq_61; // @[Misc.scala 214:29]
  wire [7:0] x1_a_bits_mask_lo_lo = {x1_a_bits_mask_acc_37,x1_a_bits_mask_acc_36,x1_a_bits_mask_acc_35,
    x1_a_bits_mask_acc_34,x1_a_bits_mask_acc_33,x1_a_bits_mask_acc_32,x1_a_bits_mask_acc_31,x1_a_bits_mask_acc_30}; // @[Cat.scala 33:92]
  wire [15:0] x1_a_bits_mask_lo = {x1_a_bits_mask_acc_45,x1_a_bits_mask_acc_44,x1_a_bits_mask_acc_43,
    x1_a_bits_mask_acc_42,x1_a_bits_mask_acc_41,x1_a_bits_mask_acc_40,x1_a_bits_mask_acc_39,x1_a_bits_mask_acc_38,
    x1_a_bits_mask_lo_lo}; // @[Cat.scala 33:92]
  wire [7:0] x1_a_bits_mask_hi_lo = {x1_a_bits_mask_acc_53,x1_a_bits_mask_acc_52,x1_a_bits_mask_acc_51,
    x1_a_bits_mask_acc_50,x1_a_bits_mask_acc_49,x1_a_bits_mask_acc_48,x1_a_bits_mask_acc_47,x1_a_bits_mask_acc_46}; // @[Cat.scala 33:92]
  wire [31:0] _x1_a_bits_mask_T_1 = {x1_a_bits_mask_acc_61,x1_a_bits_mask_acc_60,x1_a_bits_mask_acc_59,
    x1_a_bits_mask_acc_58,x1_a_bits_mask_acc_57,x1_a_bits_mask_acc_56,x1_a_bits_mask_acc_55,x1_a_bits_mask_acc_54,
    x1_a_bits_mask_hi_lo,x1_a_bits_mask_lo}; // @[Cat.scala 33:92]
  reg  x1_a_bits_mask_rdata_written_once; // @[WidthWidget.scala 57:41]
  wire  x1_a_bits_mask_masked_enable_0 = enable_0 | ~x1_a_bits_mask_rdata_written_once; // @[WidthWidget.scala 58:42]
  wire  x1_a_bits_mask_masked_enable_1 = enable_1 | ~x1_a_bits_mask_rdata_written_once; // @[WidthWidget.scala 58:42]
  wire  x1_a_bits_mask_masked_enable_2 = enable_2 | ~x1_a_bits_mask_rdata_written_once; // @[WidthWidget.scala 58:42]
  reg [7:0] x1_a_bits_mask_rdata_0; // @[WidthWidget.scala 61:24]
  reg [7:0] x1_a_bits_mask_rdata_1; // @[WidthWidget.scala 61:24]
  reg [7:0] x1_a_bits_mask_rdata_2; // @[WidthWidget.scala 61:24]
  wire [7:0] x1_a_bits_mask_mdata_0 = x1_a_bits_mask_masked_enable_0 ? auto_in_a_bits_mask : x1_a_bits_mask_rdata_0; // @[WidthWidget.scala 63:88]
  wire [7:0] x1_a_bits_mask_mdata_1 = x1_a_bits_mask_masked_enable_1 ? auto_in_a_bits_mask : x1_a_bits_mask_rdata_1; // @[WidthWidget.scala 63:88]
  wire [7:0] x1_a_bits_mask_mdata_2 = x1_a_bits_mask_masked_enable_2 ? auto_in_a_bits_mask : x1_a_bits_mask_rdata_2; // @[WidthWidget.scala 63:88]
  wire  _GEN_8 = _T & _bundleIn_0_a_ready_T | x1_a_bits_mask_rdata_written_once; // @[WidthWidget.scala 64:35 65:30 57:41]
  wire [31:0] _x1_a_bits_mask_T_5 = {auto_in_a_bits_mask,x1_a_bits_mask_mdata_2,x1_a_bits_mask_mdata_1,
    x1_a_bits_mask_mdata_0}; // @[Cat.scala 33:92]
  wire [31:0] _x1_a_bits_mask_T_7 = hasData ? _x1_a_bits_mask_T_5 : 32'hffffffff; // @[WidthWidget.scala 80:93]
  wire [255:0] cated_bits_data = {repeated_repeater_io_deq_bits_data[255:64],auto_out_d_bits_data[63:0]}; // @[Cat.scala 33:92]
  wire [2:0] cated_bits_opcode = repeated_repeater_io_deq_bits_opcode; // @[WidthWidget.scala 156:25 157:15]
  wire  repeat_hasData = cated_bits_opcode[0]; // @[Edges.scala 105:36]
  wire [2:0] cated_bits_size = repeated_repeater_io_deq_bits_size; // @[WidthWidget.scala 156:25 157:15]
  wire [11:0] _repeat_limit_T_1 = 12'h1f << cated_bits_size; // @[package.scala 235:71]
  wire [4:0] _repeat_limit_T_3 = ~_repeat_limit_T_1[4:0]; // @[package.scala 235:46]
  wire [1:0] repeat_limit = _repeat_limit_T_3[4:3]; // @[WidthWidget.scala 98:47]
  reg [1:0] repeat_count; // @[WidthWidget.scala 100:26]
  wire  repeat_first = repeat_count == 2'h0; // @[WidthWidget.scala 101:25]
  wire  repeat_last = repeat_count == repeat_limit | ~repeat_hasData; // @[WidthWidget.scala 102:35]
  wire  cated_valid = repeated_repeater_io_deq_valid; // @[WidthWidget.scala 156:25 157:15]
  wire  _repeat_T = auto_in_d_ready & cated_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _repeat_count_T_1 = repeat_count + 2'h1; // @[WidthWidget.scala 105:24]
  reg [1:0] repeat_sel_sel_sources_0; // @[WidthWidget.scala 181:27]
  reg [1:0] repeat_sel_sel_sources_1; // @[WidthWidget.scala 181:27]
  reg [1:0] repeat_sel_sel_sources_2; // @[WidthWidget.scala 181:27]
  reg [1:0] repeat_sel_sel_sources_3; // @[WidthWidget.scala 181:27]
  wire [1:0] repeat_sel_sel_a_sel = auto_in_a_bits_address[4:3]; // @[WidthWidget.scala 182:38]
  wire [1:0] cated_bits_source = repeated_repeater_io_deq_bits_source; // @[WidthWidget.scala 156:25 157:15]
  wire  repeat_sel_sel_bypass = auto_in_a_valid & auto_in_a_bits_source == cated_bits_source; // @[WidthWidget.scala 190:33]
  wire [1:0] _GEN_23 = 2'h1 == cated_bits_source ? repeat_sel_sel_sources_1 : repeat_sel_sel_sources_0; // @[WidthWidget.scala 192:{17,17}]
  wire [1:0] _GEN_24 = 2'h2 == cated_bits_source ? repeat_sel_sel_sources_2 : _GEN_23; // @[WidthWidget.scala 192:{17,17}]
  wire [1:0] _GEN_25 = 2'h3 == cated_bits_source ? repeat_sel_sel_sources_3 : _GEN_24; // @[WidthWidget.scala 192:{17,17}]
  wire [1:0] repeat_sel_sel = repeat_sel_sel_bypass ? repeat_sel_sel_a_sel : _GEN_25; // @[WidthWidget.scala 192:17]
  reg [1:0] repeat_sel_hold_r; // @[Reg.scala 19:16]
  wire [1:0] _GEN_26 = repeat_first ? repeat_sel_sel : repeat_sel_hold_r; // @[Reg.scala 19:16 20:{18,22}]
  wire [1:0] _repeat_sel_T = ~repeat_limit; // @[WidthWidget.scala 117:18]
  wire [1:0] repeat_sel = _GEN_26 & _repeat_sel_T; // @[WidthWidget.scala 117:16]
  wire [1:0] repeat_index = repeat_sel | repeat_count; // @[WidthWidget.scala 121:24]
  wire [63:0] repeat_bundleIn_0_d_bits_data_mux_0 = cated_bits_data[63:0]; // @[WidthWidget.scala 123:55]
  wire [63:0] repeat_bundleIn_0_d_bits_data_mux_1 = cated_bits_data[127:64]; // @[WidthWidget.scala 123:55]
  wire [63:0] repeat_bundleIn_0_d_bits_data_mux_2 = cated_bits_data[191:128]; // @[WidthWidget.scala 123:55]
  wire [63:0] repeat_bundleIn_0_d_bits_data_mux_3 = cated_bits_data[255:192]; // @[WidthWidget.scala 123:55]
  wire [63:0] _GEN_28 = 2'h1 == repeat_index ? repeat_bundleIn_0_d_bits_data_mux_1 : repeat_bundleIn_0_d_bits_data_mux_0
    ; // @[WidthWidget.scala 132:{30,30}]
  wire [63:0] _GEN_29 = 2'h2 == repeat_index ? repeat_bundleIn_0_d_bits_data_mux_2 : _GEN_28; // @[WidthWidget.scala 132:{30,30}]
  Repeater repeated_repeater ( // @[Repeater.scala 35:26]
    .clock(repeated_repeater_clock),
    .reset(repeated_repeater_reset),
    .io_repeat(repeated_repeater_io_repeat),
    .io_enq_ready(repeated_repeater_io_enq_ready),
    .io_enq_valid(repeated_repeater_io_enq_valid),
    .io_enq_bits_opcode(repeated_repeater_io_enq_bits_opcode),
    .io_enq_bits_size(repeated_repeater_io_enq_bits_size),
    .io_enq_bits_source(repeated_repeater_io_enq_bits_source),
    .io_enq_bits_data(repeated_repeater_io_enq_bits_data),
    .io_deq_ready(repeated_repeater_io_deq_ready),
    .io_deq_valid(repeated_repeater_io_deq_valid),
    .io_deq_bits_opcode(repeated_repeater_io_deq_bits_opcode),
    .io_deq_bits_size(repeated_repeater_io_deq_bits_size),
    .io_deq_bits_source(repeated_repeater_io_deq_bits_source),
    .io_deq_bits_data(repeated_repeater_io_deq_bits_data)
  );
  assign auto_in_a_ready = auto_out_a_ready | ~last; // @[WidthWidget.scala 71:29]
  assign auto_in_d_valid = repeated_repeater_io_deq_valid; // @[WidthWidget.scala 156:25 157:15]
  assign auto_in_d_bits_data = 2'h3 == repeat_index ? repeat_bundleIn_0_d_bits_data_mux_3 : _GEN_29; // @[WidthWidget.scala 132:{30,30}]
  assign auto_out_a_valid = auto_in_a_valid & last; // @[WidthWidget.scala 72:29]
  assign auto_out_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign auto_out_a_bits_mask = _x1_a_bits_mask_T_1 & _x1_a_bits_mask_T_7; // @[WidthWidget.scala 80:88]
  assign auto_out_a_bits_data = {x1_a_bits_data_hi,x1_a_bits_data_lo}; // @[Cat.scala 33:92]
  assign auto_out_d_ready = repeated_repeater_io_enq_ready; // @[Nodes.scala 1212:84 Repeater.scala 37:21]
  assign repeated_repeater_clock = clock;
  assign repeated_repeater_reset = reset;
  assign repeated_repeater_io_repeat = ~repeat_last; // @[WidthWidget.scala 143:7]
  assign repeated_repeater_io_enq_valid = auto_out_d_valid; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign repeated_repeater_io_enq_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign repeated_repeater_io_enq_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign repeated_repeater_io_enq_bits_source = auto_out_d_bits_source; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign repeated_repeater_io_enq_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign repeated_repeater_io_deq_ready = auto_in_d_ready; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  always @(posedge clock) begin
    if (reset) begin // @[WidthWidget.scala 35:27]
      count <= 2'h0; // @[WidthWidget.scala 35:27]
    end else if (_T) begin // @[WidthWidget.scala 44:24]
      if (last) begin // @[WidthWidget.scala 47:21]
        count <= 2'h0; // @[WidthWidget.scala 48:17]
      end else begin
        count <= _count_T_1; // @[WidthWidget.scala 45:15]
      end
    end
    if (reset) begin // @[WidthWidget.scala 57:41]
      x1_a_bits_data_rdata_written_once <= 1'h0; // @[WidthWidget.scala 57:41]
    end else begin
      x1_a_bits_data_rdata_written_once <= _GEN_4;
    end
    if (_T & _bundleIn_0_a_ready_T) begin // @[WidthWidget.scala 64:35]
      if (x1_a_bits_data_masked_enable_0) begin // @[WidthWidget.scala 63:88]
        x1_a_bits_data_rdata_0 <= auto_in_a_bits_data;
      end
    end
    if (_T & _bundleIn_0_a_ready_T) begin // @[WidthWidget.scala 64:35]
      if (x1_a_bits_data_masked_enable_1) begin // @[WidthWidget.scala 63:88]
        x1_a_bits_data_rdata_1 <= auto_in_a_bits_data;
      end
    end
    if (_T & _bundleIn_0_a_ready_T) begin // @[WidthWidget.scala 64:35]
      if (x1_a_bits_data_masked_enable_2) begin // @[WidthWidget.scala 63:88]
        x1_a_bits_data_rdata_2 <= auto_in_a_bits_data;
      end
    end
    if (reset) begin // @[WidthWidget.scala 57:41]
      x1_a_bits_mask_rdata_written_once <= 1'h0; // @[WidthWidget.scala 57:41]
    end else begin
      x1_a_bits_mask_rdata_written_once <= _GEN_8;
    end
    if (_T & _bundleIn_0_a_ready_T) begin // @[WidthWidget.scala 64:35]
      if (x1_a_bits_mask_masked_enable_0) begin // @[WidthWidget.scala 63:88]
        x1_a_bits_mask_rdata_0 <= auto_in_a_bits_mask;
      end
    end
    if (_T & _bundleIn_0_a_ready_T) begin // @[WidthWidget.scala 64:35]
      if (x1_a_bits_mask_masked_enable_1) begin // @[WidthWidget.scala 63:88]
        x1_a_bits_mask_rdata_1 <= auto_in_a_bits_mask;
      end
    end
    if (_T & _bundleIn_0_a_ready_T) begin // @[WidthWidget.scala 64:35]
      if (x1_a_bits_mask_masked_enable_2) begin // @[WidthWidget.scala 63:88]
        x1_a_bits_mask_rdata_2 <= auto_in_a_bits_mask;
      end
    end
    if (reset) begin // @[WidthWidget.scala 100:26]
      repeat_count <= 2'h0; // @[WidthWidget.scala 100:26]
    end else if (_repeat_T) begin // @[WidthWidget.scala 104:25]
      if (repeat_last) begin // @[WidthWidget.scala 106:21]
        repeat_count <= 2'h0; // @[WidthWidget.scala 106:29]
      end else begin
        repeat_count <= _repeat_count_T_1; // @[WidthWidget.scala 105:15]
      end
    end
    if (_T) begin // @[WidthWidget.scala 183:28]
      if (2'h0 == auto_in_a_bits_source) begin // @[WidthWidget.scala 184:37]
        repeat_sel_sel_sources_0 <= repeat_sel_sel_a_sel; // @[WidthWidget.scala 184:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 183:28]
      if (2'h1 == auto_in_a_bits_source) begin // @[WidthWidget.scala 184:37]
        repeat_sel_sel_sources_1 <= repeat_sel_sel_a_sel; // @[WidthWidget.scala 184:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 183:28]
      if (2'h2 == auto_in_a_bits_source) begin // @[WidthWidget.scala 184:37]
        repeat_sel_sel_sources_2 <= repeat_sel_sel_a_sel; // @[WidthWidget.scala 184:37]
      end
    end
    if (_T) begin // @[WidthWidget.scala 183:28]
      if (2'h3 == auto_in_a_bits_source) begin // @[WidthWidget.scala 184:37]
        repeat_sel_sel_sources_3 <= repeat_sel_sel_a_sel; // @[WidthWidget.scala 184:37]
      end
    end
    if (repeat_first) begin // @[Reg.scala 20:18]
      if (repeat_sel_sel_bypass) begin // @[WidthWidget.scala 192:17]
        repeat_sel_hold_r <= repeat_sel_sel_a_sel;
      end else if (2'h3 == cated_bits_source) begin // @[WidthWidget.scala 192:17]
        repeat_sel_hold_r <= repeat_sel_sel_sources_3; // @[WidthWidget.scala 192:17]
      end else if (2'h2 == cated_bits_source) begin // @[WidthWidget.scala 192:17]
        repeat_sel_hold_r <= repeat_sel_sel_sources_2; // @[WidthWidget.scala 192:17]
      end else begin
        repeat_sel_hold_r <= _GEN_23;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  x1_a_bits_data_rdata_written_once = _RAND_1[0:0];
  _RAND_2 = {2{`RANDOM}};
  x1_a_bits_data_rdata_0 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  x1_a_bits_data_rdata_1 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  x1_a_bits_data_rdata_2 = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  x1_a_bits_mask_rdata_written_once = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  x1_a_bits_mask_rdata_0 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  x1_a_bits_mask_rdata_1 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  x1_a_bits_mask_rdata_2 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  repeat_count = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  repeat_sel_sel_sources_0 = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  repeat_sel_sel_sources_1 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  repeat_sel_sel_sources_2 = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  repeat_sel_sel_sources_3 = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  repeat_sel_hold_r = _RAND_14[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MaxPeriodFibonacciLFSR(
  input   clock,
  input   reset,
  output  io_out_0,
  output  io_out_1,
  output  io_out_2,
  output  io_out_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg  state_0; // @[PRNG.scala 55:49]
  reg  state_1; // @[PRNG.scala 55:49]
  reg  state_2; // @[PRNG.scala 55:49]
  reg  state_3; // @[PRNG.scala 55:49]
  wire  _T = state_3 ^ state_2; // @[LFSR.scala 15:41]
  assign io_out_0 = state_0; // @[PRNG.scala 78:10]
  assign io_out_1 = state_1; // @[PRNG.scala 78:10]
  assign io_out_2 = state_2; // @[PRNG.scala 78:10]
  assign io_out_3 = state_3; // @[PRNG.scala 78:10]
  always @(posedge clock) begin
    state_0 <= reset | _T; // @[PRNG.scala 55:{49,49}]
    if (reset) begin // @[PRNG.scala 55:49]
      state_1 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_1 <= state_0;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_2 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_2 <= state_1;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_3 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_3 <= state_2;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  state_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  state_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  state_3 = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BPU(
  input         clock,
  input         reset,
  input  [63:0] io_pc,
  input  [63:0] io_jmp_packet_target,
  input         io_jmp_packet_bp_update,
  input         io_jmp_packet_bp_taken,
  input  [63:0] io_jmp_packet_bp_pc,
  output [63:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [63:0] _RAND_513;
  reg [63:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [63:0] _RAND_516;
  reg [63:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [63:0] _RAND_519;
  reg [63:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [63:0] _RAND_522;
  reg [63:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [63:0] _RAND_525;
  reg [63:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [63:0] _RAND_528;
  reg [63:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [63:0] _RAND_531;
  reg [63:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [63:0] _RAND_534;
  reg [63:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [63:0] _RAND_537;
  reg [63:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [63:0] _RAND_540;
  reg [63:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [63:0] _RAND_543;
  reg [63:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [63:0] _RAND_546;
  reg [63:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [63:0] _RAND_549;
  reg [63:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [63:0] _RAND_552;
  reg [63:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [63:0] _RAND_555;
  reg [63:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [63:0] _RAND_558;
  reg [63:0] _RAND_559;
  reg [31:0] _RAND_560;
`endif // RANDOMIZE_REG_INIT
  wire  btb_replace_idx_prng_clock; // @[PRNG.scala 91:22]
  wire  btb_replace_idx_prng_reset; // @[PRNG.scala 91:22]
  wire  btb_replace_idx_prng_io_out_0; // @[PRNG.scala 91:22]
  wire  btb_replace_idx_prng_io_out_1; // @[PRNG.scala 91:22]
  wire  btb_replace_idx_prng_io_out_2; // @[PRNG.scala 91:22]
  wire  btb_replace_idx_prng_io_out_3; // @[PRNG.scala 91:22]
  reg [8:0] ghr; // @[BPU.scala 26:20]
  reg [1:0] pht_0; // @[BPU.scala 27:20]
  reg [1:0] pht_1; // @[BPU.scala 27:20]
  reg [1:0] pht_2; // @[BPU.scala 27:20]
  reg [1:0] pht_3; // @[BPU.scala 27:20]
  reg [1:0] pht_4; // @[BPU.scala 27:20]
  reg [1:0] pht_5; // @[BPU.scala 27:20]
  reg [1:0] pht_6; // @[BPU.scala 27:20]
  reg [1:0] pht_7; // @[BPU.scala 27:20]
  reg [1:0] pht_8; // @[BPU.scala 27:20]
  reg [1:0] pht_9; // @[BPU.scala 27:20]
  reg [1:0] pht_10; // @[BPU.scala 27:20]
  reg [1:0] pht_11; // @[BPU.scala 27:20]
  reg [1:0] pht_12; // @[BPU.scala 27:20]
  reg [1:0] pht_13; // @[BPU.scala 27:20]
  reg [1:0] pht_14; // @[BPU.scala 27:20]
  reg [1:0] pht_15; // @[BPU.scala 27:20]
  reg [1:0] pht_16; // @[BPU.scala 27:20]
  reg [1:0] pht_17; // @[BPU.scala 27:20]
  reg [1:0] pht_18; // @[BPU.scala 27:20]
  reg [1:0] pht_19; // @[BPU.scala 27:20]
  reg [1:0] pht_20; // @[BPU.scala 27:20]
  reg [1:0] pht_21; // @[BPU.scala 27:20]
  reg [1:0] pht_22; // @[BPU.scala 27:20]
  reg [1:0] pht_23; // @[BPU.scala 27:20]
  reg [1:0] pht_24; // @[BPU.scala 27:20]
  reg [1:0] pht_25; // @[BPU.scala 27:20]
  reg [1:0] pht_26; // @[BPU.scala 27:20]
  reg [1:0] pht_27; // @[BPU.scala 27:20]
  reg [1:0] pht_28; // @[BPU.scala 27:20]
  reg [1:0] pht_29; // @[BPU.scala 27:20]
  reg [1:0] pht_30; // @[BPU.scala 27:20]
  reg [1:0] pht_31; // @[BPU.scala 27:20]
  reg [1:0] pht_32; // @[BPU.scala 27:20]
  reg [1:0] pht_33; // @[BPU.scala 27:20]
  reg [1:0] pht_34; // @[BPU.scala 27:20]
  reg [1:0] pht_35; // @[BPU.scala 27:20]
  reg [1:0] pht_36; // @[BPU.scala 27:20]
  reg [1:0] pht_37; // @[BPU.scala 27:20]
  reg [1:0] pht_38; // @[BPU.scala 27:20]
  reg [1:0] pht_39; // @[BPU.scala 27:20]
  reg [1:0] pht_40; // @[BPU.scala 27:20]
  reg [1:0] pht_41; // @[BPU.scala 27:20]
  reg [1:0] pht_42; // @[BPU.scala 27:20]
  reg [1:0] pht_43; // @[BPU.scala 27:20]
  reg [1:0] pht_44; // @[BPU.scala 27:20]
  reg [1:0] pht_45; // @[BPU.scala 27:20]
  reg [1:0] pht_46; // @[BPU.scala 27:20]
  reg [1:0] pht_47; // @[BPU.scala 27:20]
  reg [1:0] pht_48; // @[BPU.scala 27:20]
  reg [1:0] pht_49; // @[BPU.scala 27:20]
  reg [1:0] pht_50; // @[BPU.scala 27:20]
  reg [1:0] pht_51; // @[BPU.scala 27:20]
  reg [1:0] pht_52; // @[BPU.scala 27:20]
  reg [1:0] pht_53; // @[BPU.scala 27:20]
  reg [1:0] pht_54; // @[BPU.scala 27:20]
  reg [1:0] pht_55; // @[BPU.scala 27:20]
  reg [1:0] pht_56; // @[BPU.scala 27:20]
  reg [1:0] pht_57; // @[BPU.scala 27:20]
  reg [1:0] pht_58; // @[BPU.scala 27:20]
  reg [1:0] pht_59; // @[BPU.scala 27:20]
  reg [1:0] pht_60; // @[BPU.scala 27:20]
  reg [1:0] pht_61; // @[BPU.scala 27:20]
  reg [1:0] pht_62; // @[BPU.scala 27:20]
  reg [1:0] pht_63; // @[BPU.scala 27:20]
  reg [1:0] pht_64; // @[BPU.scala 27:20]
  reg [1:0] pht_65; // @[BPU.scala 27:20]
  reg [1:0] pht_66; // @[BPU.scala 27:20]
  reg [1:0] pht_67; // @[BPU.scala 27:20]
  reg [1:0] pht_68; // @[BPU.scala 27:20]
  reg [1:0] pht_69; // @[BPU.scala 27:20]
  reg [1:0] pht_70; // @[BPU.scala 27:20]
  reg [1:0] pht_71; // @[BPU.scala 27:20]
  reg [1:0] pht_72; // @[BPU.scala 27:20]
  reg [1:0] pht_73; // @[BPU.scala 27:20]
  reg [1:0] pht_74; // @[BPU.scala 27:20]
  reg [1:0] pht_75; // @[BPU.scala 27:20]
  reg [1:0] pht_76; // @[BPU.scala 27:20]
  reg [1:0] pht_77; // @[BPU.scala 27:20]
  reg [1:0] pht_78; // @[BPU.scala 27:20]
  reg [1:0] pht_79; // @[BPU.scala 27:20]
  reg [1:0] pht_80; // @[BPU.scala 27:20]
  reg [1:0] pht_81; // @[BPU.scala 27:20]
  reg [1:0] pht_82; // @[BPU.scala 27:20]
  reg [1:0] pht_83; // @[BPU.scala 27:20]
  reg [1:0] pht_84; // @[BPU.scala 27:20]
  reg [1:0] pht_85; // @[BPU.scala 27:20]
  reg [1:0] pht_86; // @[BPU.scala 27:20]
  reg [1:0] pht_87; // @[BPU.scala 27:20]
  reg [1:0] pht_88; // @[BPU.scala 27:20]
  reg [1:0] pht_89; // @[BPU.scala 27:20]
  reg [1:0] pht_90; // @[BPU.scala 27:20]
  reg [1:0] pht_91; // @[BPU.scala 27:20]
  reg [1:0] pht_92; // @[BPU.scala 27:20]
  reg [1:0] pht_93; // @[BPU.scala 27:20]
  reg [1:0] pht_94; // @[BPU.scala 27:20]
  reg [1:0] pht_95; // @[BPU.scala 27:20]
  reg [1:0] pht_96; // @[BPU.scala 27:20]
  reg [1:0] pht_97; // @[BPU.scala 27:20]
  reg [1:0] pht_98; // @[BPU.scala 27:20]
  reg [1:0] pht_99; // @[BPU.scala 27:20]
  reg [1:0] pht_100; // @[BPU.scala 27:20]
  reg [1:0] pht_101; // @[BPU.scala 27:20]
  reg [1:0] pht_102; // @[BPU.scala 27:20]
  reg [1:0] pht_103; // @[BPU.scala 27:20]
  reg [1:0] pht_104; // @[BPU.scala 27:20]
  reg [1:0] pht_105; // @[BPU.scala 27:20]
  reg [1:0] pht_106; // @[BPU.scala 27:20]
  reg [1:0] pht_107; // @[BPU.scala 27:20]
  reg [1:0] pht_108; // @[BPU.scala 27:20]
  reg [1:0] pht_109; // @[BPU.scala 27:20]
  reg [1:0] pht_110; // @[BPU.scala 27:20]
  reg [1:0] pht_111; // @[BPU.scala 27:20]
  reg [1:0] pht_112; // @[BPU.scala 27:20]
  reg [1:0] pht_113; // @[BPU.scala 27:20]
  reg [1:0] pht_114; // @[BPU.scala 27:20]
  reg [1:0] pht_115; // @[BPU.scala 27:20]
  reg [1:0] pht_116; // @[BPU.scala 27:20]
  reg [1:0] pht_117; // @[BPU.scala 27:20]
  reg [1:0] pht_118; // @[BPU.scala 27:20]
  reg [1:0] pht_119; // @[BPU.scala 27:20]
  reg [1:0] pht_120; // @[BPU.scala 27:20]
  reg [1:0] pht_121; // @[BPU.scala 27:20]
  reg [1:0] pht_122; // @[BPU.scala 27:20]
  reg [1:0] pht_123; // @[BPU.scala 27:20]
  reg [1:0] pht_124; // @[BPU.scala 27:20]
  reg [1:0] pht_125; // @[BPU.scala 27:20]
  reg [1:0] pht_126; // @[BPU.scala 27:20]
  reg [1:0] pht_127; // @[BPU.scala 27:20]
  reg [1:0] pht_128; // @[BPU.scala 27:20]
  reg [1:0] pht_129; // @[BPU.scala 27:20]
  reg [1:0] pht_130; // @[BPU.scala 27:20]
  reg [1:0] pht_131; // @[BPU.scala 27:20]
  reg [1:0] pht_132; // @[BPU.scala 27:20]
  reg [1:0] pht_133; // @[BPU.scala 27:20]
  reg [1:0] pht_134; // @[BPU.scala 27:20]
  reg [1:0] pht_135; // @[BPU.scala 27:20]
  reg [1:0] pht_136; // @[BPU.scala 27:20]
  reg [1:0] pht_137; // @[BPU.scala 27:20]
  reg [1:0] pht_138; // @[BPU.scala 27:20]
  reg [1:0] pht_139; // @[BPU.scala 27:20]
  reg [1:0] pht_140; // @[BPU.scala 27:20]
  reg [1:0] pht_141; // @[BPU.scala 27:20]
  reg [1:0] pht_142; // @[BPU.scala 27:20]
  reg [1:0] pht_143; // @[BPU.scala 27:20]
  reg [1:0] pht_144; // @[BPU.scala 27:20]
  reg [1:0] pht_145; // @[BPU.scala 27:20]
  reg [1:0] pht_146; // @[BPU.scala 27:20]
  reg [1:0] pht_147; // @[BPU.scala 27:20]
  reg [1:0] pht_148; // @[BPU.scala 27:20]
  reg [1:0] pht_149; // @[BPU.scala 27:20]
  reg [1:0] pht_150; // @[BPU.scala 27:20]
  reg [1:0] pht_151; // @[BPU.scala 27:20]
  reg [1:0] pht_152; // @[BPU.scala 27:20]
  reg [1:0] pht_153; // @[BPU.scala 27:20]
  reg [1:0] pht_154; // @[BPU.scala 27:20]
  reg [1:0] pht_155; // @[BPU.scala 27:20]
  reg [1:0] pht_156; // @[BPU.scala 27:20]
  reg [1:0] pht_157; // @[BPU.scala 27:20]
  reg [1:0] pht_158; // @[BPU.scala 27:20]
  reg [1:0] pht_159; // @[BPU.scala 27:20]
  reg [1:0] pht_160; // @[BPU.scala 27:20]
  reg [1:0] pht_161; // @[BPU.scala 27:20]
  reg [1:0] pht_162; // @[BPU.scala 27:20]
  reg [1:0] pht_163; // @[BPU.scala 27:20]
  reg [1:0] pht_164; // @[BPU.scala 27:20]
  reg [1:0] pht_165; // @[BPU.scala 27:20]
  reg [1:0] pht_166; // @[BPU.scala 27:20]
  reg [1:0] pht_167; // @[BPU.scala 27:20]
  reg [1:0] pht_168; // @[BPU.scala 27:20]
  reg [1:0] pht_169; // @[BPU.scala 27:20]
  reg [1:0] pht_170; // @[BPU.scala 27:20]
  reg [1:0] pht_171; // @[BPU.scala 27:20]
  reg [1:0] pht_172; // @[BPU.scala 27:20]
  reg [1:0] pht_173; // @[BPU.scala 27:20]
  reg [1:0] pht_174; // @[BPU.scala 27:20]
  reg [1:0] pht_175; // @[BPU.scala 27:20]
  reg [1:0] pht_176; // @[BPU.scala 27:20]
  reg [1:0] pht_177; // @[BPU.scala 27:20]
  reg [1:0] pht_178; // @[BPU.scala 27:20]
  reg [1:0] pht_179; // @[BPU.scala 27:20]
  reg [1:0] pht_180; // @[BPU.scala 27:20]
  reg [1:0] pht_181; // @[BPU.scala 27:20]
  reg [1:0] pht_182; // @[BPU.scala 27:20]
  reg [1:0] pht_183; // @[BPU.scala 27:20]
  reg [1:0] pht_184; // @[BPU.scala 27:20]
  reg [1:0] pht_185; // @[BPU.scala 27:20]
  reg [1:0] pht_186; // @[BPU.scala 27:20]
  reg [1:0] pht_187; // @[BPU.scala 27:20]
  reg [1:0] pht_188; // @[BPU.scala 27:20]
  reg [1:0] pht_189; // @[BPU.scala 27:20]
  reg [1:0] pht_190; // @[BPU.scala 27:20]
  reg [1:0] pht_191; // @[BPU.scala 27:20]
  reg [1:0] pht_192; // @[BPU.scala 27:20]
  reg [1:0] pht_193; // @[BPU.scala 27:20]
  reg [1:0] pht_194; // @[BPU.scala 27:20]
  reg [1:0] pht_195; // @[BPU.scala 27:20]
  reg [1:0] pht_196; // @[BPU.scala 27:20]
  reg [1:0] pht_197; // @[BPU.scala 27:20]
  reg [1:0] pht_198; // @[BPU.scala 27:20]
  reg [1:0] pht_199; // @[BPU.scala 27:20]
  reg [1:0] pht_200; // @[BPU.scala 27:20]
  reg [1:0] pht_201; // @[BPU.scala 27:20]
  reg [1:0] pht_202; // @[BPU.scala 27:20]
  reg [1:0] pht_203; // @[BPU.scala 27:20]
  reg [1:0] pht_204; // @[BPU.scala 27:20]
  reg [1:0] pht_205; // @[BPU.scala 27:20]
  reg [1:0] pht_206; // @[BPU.scala 27:20]
  reg [1:0] pht_207; // @[BPU.scala 27:20]
  reg [1:0] pht_208; // @[BPU.scala 27:20]
  reg [1:0] pht_209; // @[BPU.scala 27:20]
  reg [1:0] pht_210; // @[BPU.scala 27:20]
  reg [1:0] pht_211; // @[BPU.scala 27:20]
  reg [1:0] pht_212; // @[BPU.scala 27:20]
  reg [1:0] pht_213; // @[BPU.scala 27:20]
  reg [1:0] pht_214; // @[BPU.scala 27:20]
  reg [1:0] pht_215; // @[BPU.scala 27:20]
  reg [1:0] pht_216; // @[BPU.scala 27:20]
  reg [1:0] pht_217; // @[BPU.scala 27:20]
  reg [1:0] pht_218; // @[BPU.scala 27:20]
  reg [1:0] pht_219; // @[BPU.scala 27:20]
  reg [1:0] pht_220; // @[BPU.scala 27:20]
  reg [1:0] pht_221; // @[BPU.scala 27:20]
  reg [1:0] pht_222; // @[BPU.scala 27:20]
  reg [1:0] pht_223; // @[BPU.scala 27:20]
  reg [1:0] pht_224; // @[BPU.scala 27:20]
  reg [1:0] pht_225; // @[BPU.scala 27:20]
  reg [1:0] pht_226; // @[BPU.scala 27:20]
  reg [1:0] pht_227; // @[BPU.scala 27:20]
  reg [1:0] pht_228; // @[BPU.scala 27:20]
  reg [1:0] pht_229; // @[BPU.scala 27:20]
  reg [1:0] pht_230; // @[BPU.scala 27:20]
  reg [1:0] pht_231; // @[BPU.scala 27:20]
  reg [1:0] pht_232; // @[BPU.scala 27:20]
  reg [1:0] pht_233; // @[BPU.scala 27:20]
  reg [1:0] pht_234; // @[BPU.scala 27:20]
  reg [1:0] pht_235; // @[BPU.scala 27:20]
  reg [1:0] pht_236; // @[BPU.scala 27:20]
  reg [1:0] pht_237; // @[BPU.scala 27:20]
  reg [1:0] pht_238; // @[BPU.scala 27:20]
  reg [1:0] pht_239; // @[BPU.scala 27:20]
  reg [1:0] pht_240; // @[BPU.scala 27:20]
  reg [1:0] pht_241; // @[BPU.scala 27:20]
  reg [1:0] pht_242; // @[BPU.scala 27:20]
  reg [1:0] pht_243; // @[BPU.scala 27:20]
  reg [1:0] pht_244; // @[BPU.scala 27:20]
  reg [1:0] pht_245; // @[BPU.scala 27:20]
  reg [1:0] pht_246; // @[BPU.scala 27:20]
  reg [1:0] pht_247; // @[BPU.scala 27:20]
  reg [1:0] pht_248; // @[BPU.scala 27:20]
  reg [1:0] pht_249; // @[BPU.scala 27:20]
  reg [1:0] pht_250; // @[BPU.scala 27:20]
  reg [1:0] pht_251; // @[BPU.scala 27:20]
  reg [1:0] pht_252; // @[BPU.scala 27:20]
  reg [1:0] pht_253; // @[BPU.scala 27:20]
  reg [1:0] pht_254; // @[BPU.scala 27:20]
  reg [1:0] pht_255; // @[BPU.scala 27:20]
  reg [1:0] pht_256; // @[BPU.scala 27:20]
  reg [1:0] pht_257; // @[BPU.scala 27:20]
  reg [1:0] pht_258; // @[BPU.scala 27:20]
  reg [1:0] pht_259; // @[BPU.scala 27:20]
  reg [1:0] pht_260; // @[BPU.scala 27:20]
  reg [1:0] pht_261; // @[BPU.scala 27:20]
  reg [1:0] pht_262; // @[BPU.scala 27:20]
  reg [1:0] pht_263; // @[BPU.scala 27:20]
  reg [1:0] pht_264; // @[BPU.scala 27:20]
  reg [1:0] pht_265; // @[BPU.scala 27:20]
  reg [1:0] pht_266; // @[BPU.scala 27:20]
  reg [1:0] pht_267; // @[BPU.scala 27:20]
  reg [1:0] pht_268; // @[BPU.scala 27:20]
  reg [1:0] pht_269; // @[BPU.scala 27:20]
  reg [1:0] pht_270; // @[BPU.scala 27:20]
  reg [1:0] pht_271; // @[BPU.scala 27:20]
  reg [1:0] pht_272; // @[BPU.scala 27:20]
  reg [1:0] pht_273; // @[BPU.scala 27:20]
  reg [1:0] pht_274; // @[BPU.scala 27:20]
  reg [1:0] pht_275; // @[BPU.scala 27:20]
  reg [1:0] pht_276; // @[BPU.scala 27:20]
  reg [1:0] pht_277; // @[BPU.scala 27:20]
  reg [1:0] pht_278; // @[BPU.scala 27:20]
  reg [1:0] pht_279; // @[BPU.scala 27:20]
  reg [1:0] pht_280; // @[BPU.scala 27:20]
  reg [1:0] pht_281; // @[BPU.scala 27:20]
  reg [1:0] pht_282; // @[BPU.scala 27:20]
  reg [1:0] pht_283; // @[BPU.scala 27:20]
  reg [1:0] pht_284; // @[BPU.scala 27:20]
  reg [1:0] pht_285; // @[BPU.scala 27:20]
  reg [1:0] pht_286; // @[BPU.scala 27:20]
  reg [1:0] pht_287; // @[BPU.scala 27:20]
  reg [1:0] pht_288; // @[BPU.scala 27:20]
  reg [1:0] pht_289; // @[BPU.scala 27:20]
  reg [1:0] pht_290; // @[BPU.scala 27:20]
  reg [1:0] pht_291; // @[BPU.scala 27:20]
  reg [1:0] pht_292; // @[BPU.scala 27:20]
  reg [1:0] pht_293; // @[BPU.scala 27:20]
  reg [1:0] pht_294; // @[BPU.scala 27:20]
  reg [1:0] pht_295; // @[BPU.scala 27:20]
  reg [1:0] pht_296; // @[BPU.scala 27:20]
  reg [1:0] pht_297; // @[BPU.scala 27:20]
  reg [1:0] pht_298; // @[BPU.scala 27:20]
  reg [1:0] pht_299; // @[BPU.scala 27:20]
  reg [1:0] pht_300; // @[BPU.scala 27:20]
  reg [1:0] pht_301; // @[BPU.scala 27:20]
  reg [1:0] pht_302; // @[BPU.scala 27:20]
  reg [1:0] pht_303; // @[BPU.scala 27:20]
  reg [1:0] pht_304; // @[BPU.scala 27:20]
  reg [1:0] pht_305; // @[BPU.scala 27:20]
  reg [1:0] pht_306; // @[BPU.scala 27:20]
  reg [1:0] pht_307; // @[BPU.scala 27:20]
  reg [1:0] pht_308; // @[BPU.scala 27:20]
  reg [1:0] pht_309; // @[BPU.scala 27:20]
  reg [1:0] pht_310; // @[BPU.scala 27:20]
  reg [1:0] pht_311; // @[BPU.scala 27:20]
  reg [1:0] pht_312; // @[BPU.scala 27:20]
  reg [1:0] pht_313; // @[BPU.scala 27:20]
  reg [1:0] pht_314; // @[BPU.scala 27:20]
  reg [1:0] pht_315; // @[BPU.scala 27:20]
  reg [1:0] pht_316; // @[BPU.scala 27:20]
  reg [1:0] pht_317; // @[BPU.scala 27:20]
  reg [1:0] pht_318; // @[BPU.scala 27:20]
  reg [1:0] pht_319; // @[BPU.scala 27:20]
  reg [1:0] pht_320; // @[BPU.scala 27:20]
  reg [1:0] pht_321; // @[BPU.scala 27:20]
  reg [1:0] pht_322; // @[BPU.scala 27:20]
  reg [1:0] pht_323; // @[BPU.scala 27:20]
  reg [1:0] pht_324; // @[BPU.scala 27:20]
  reg [1:0] pht_325; // @[BPU.scala 27:20]
  reg [1:0] pht_326; // @[BPU.scala 27:20]
  reg [1:0] pht_327; // @[BPU.scala 27:20]
  reg [1:0] pht_328; // @[BPU.scala 27:20]
  reg [1:0] pht_329; // @[BPU.scala 27:20]
  reg [1:0] pht_330; // @[BPU.scala 27:20]
  reg [1:0] pht_331; // @[BPU.scala 27:20]
  reg [1:0] pht_332; // @[BPU.scala 27:20]
  reg [1:0] pht_333; // @[BPU.scala 27:20]
  reg [1:0] pht_334; // @[BPU.scala 27:20]
  reg [1:0] pht_335; // @[BPU.scala 27:20]
  reg [1:0] pht_336; // @[BPU.scala 27:20]
  reg [1:0] pht_337; // @[BPU.scala 27:20]
  reg [1:0] pht_338; // @[BPU.scala 27:20]
  reg [1:0] pht_339; // @[BPU.scala 27:20]
  reg [1:0] pht_340; // @[BPU.scala 27:20]
  reg [1:0] pht_341; // @[BPU.scala 27:20]
  reg [1:0] pht_342; // @[BPU.scala 27:20]
  reg [1:0] pht_343; // @[BPU.scala 27:20]
  reg [1:0] pht_344; // @[BPU.scala 27:20]
  reg [1:0] pht_345; // @[BPU.scala 27:20]
  reg [1:0] pht_346; // @[BPU.scala 27:20]
  reg [1:0] pht_347; // @[BPU.scala 27:20]
  reg [1:0] pht_348; // @[BPU.scala 27:20]
  reg [1:0] pht_349; // @[BPU.scala 27:20]
  reg [1:0] pht_350; // @[BPU.scala 27:20]
  reg [1:0] pht_351; // @[BPU.scala 27:20]
  reg [1:0] pht_352; // @[BPU.scala 27:20]
  reg [1:0] pht_353; // @[BPU.scala 27:20]
  reg [1:0] pht_354; // @[BPU.scala 27:20]
  reg [1:0] pht_355; // @[BPU.scala 27:20]
  reg [1:0] pht_356; // @[BPU.scala 27:20]
  reg [1:0] pht_357; // @[BPU.scala 27:20]
  reg [1:0] pht_358; // @[BPU.scala 27:20]
  reg [1:0] pht_359; // @[BPU.scala 27:20]
  reg [1:0] pht_360; // @[BPU.scala 27:20]
  reg [1:0] pht_361; // @[BPU.scala 27:20]
  reg [1:0] pht_362; // @[BPU.scala 27:20]
  reg [1:0] pht_363; // @[BPU.scala 27:20]
  reg [1:0] pht_364; // @[BPU.scala 27:20]
  reg [1:0] pht_365; // @[BPU.scala 27:20]
  reg [1:0] pht_366; // @[BPU.scala 27:20]
  reg [1:0] pht_367; // @[BPU.scala 27:20]
  reg [1:0] pht_368; // @[BPU.scala 27:20]
  reg [1:0] pht_369; // @[BPU.scala 27:20]
  reg [1:0] pht_370; // @[BPU.scala 27:20]
  reg [1:0] pht_371; // @[BPU.scala 27:20]
  reg [1:0] pht_372; // @[BPU.scala 27:20]
  reg [1:0] pht_373; // @[BPU.scala 27:20]
  reg [1:0] pht_374; // @[BPU.scala 27:20]
  reg [1:0] pht_375; // @[BPU.scala 27:20]
  reg [1:0] pht_376; // @[BPU.scala 27:20]
  reg [1:0] pht_377; // @[BPU.scala 27:20]
  reg [1:0] pht_378; // @[BPU.scala 27:20]
  reg [1:0] pht_379; // @[BPU.scala 27:20]
  reg [1:0] pht_380; // @[BPU.scala 27:20]
  reg [1:0] pht_381; // @[BPU.scala 27:20]
  reg [1:0] pht_382; // @[BPU.scala 27:20]
  reg [1:0] pht_383; // @[BPU.scala 27:20]
  reg [1:0] pht_384; // @[BPU.scala 27:20]
  reg [1:0] pht_385; // @[BPU.scala 27:20]
  reg [1:0] pht_386; // @[BPU.scala 27:20]
  reg [1:0] pht_387; // @[BPU.scala 27:20]
  reg [1:0] pht_388; // @[BPU.scala 27:20]
  reg [1:0] pht_389; // @[BPU.scala 27:20]
  reg [1:0] pht_390; // @[BPU.scala 27:20]
  reg [1:0] pht_391; // @[BPU.scala 27:20]
  reg [1:0] pht_392; // @[BPU.scala 27:20]
  reg [1:0] pht_393; // @[BPU.scala 27:20]
  reg [1:0] pht_394; // @[BPU.scala 27:20]
  reg [1:0] pht_395; // @[BPU.scala 27:20]
  reg [1:0] pht_396; // @[BPU.scala 27:20]
  reg [1:0] pht_397; // @[BPU.scala 27:20]
  reg [1:0] pht_398; // @[BPU.scala 27:20]
  reg [1:0] pht_399; // @[BPU.scala 27:20]
  reg [1:0] pht_400; // @[BPU.scala 27:20]
  reg [1:0] pht_401; // @[BPU.scala 27:20]
  reg [1:0] pht_402; // @[BPU.scala 27:20]
  reg [1:0] pht_403; // @[BPU.scala 27:20]
  reg [1:0] pht_404; // @[BPU.scala 27:20]
  reg [1:0] pht_405; // @[BPU.scala 27:20]
  reg [1:0] pht_406; // @[BPU.scala 27:20]
  reg [1:0] pht_407; // @[BPU.scala 27:20]
  reg [1:0] pht_408; // @[BPU.scala 27:20]
  reg [1:0] pht_409; // @[BPU.scala 27:20]
  reg [1:0] pht_410; // @[BPU.scala 27:20]
  reg [1:0] pht_411; // @[BPU.scala 27:20]
  reg [1:0] pht_412; // @[BPU.scala 27:20]
  reg [1:0] pht_413; // @[BPU.scala 27:20]
  reg [1:0] pht_414; // @[BPU.scala 27:20]
  reg [1:0] pht_415; // @[BPU.scala 27:20]
  reg [1:0] pht_416; // @[BPU.scala 27:20]
  reg [1:0] pht_417; // @[BPU.scala 27:20]
  reg [1:0] pht_418; // @[BPU.scala 27:20]
  reg [1:0] pht_419; // @[BPU.scala 27:20]
  reg [1:0] pht_420; // @[BPU.scala 27:20]
  reg [1:0] pht_421; // @[BPU.scala 27:20]
  reg [1:0] pht_422; // @[BPU.scala 27:20]
  reg [1:0] pht_423; // @[BPU.scala 27:20]
  reg [1:0] pht_424; // @[BPU.scala 27:20]
  reg [1:0] pht_425; // @[BPU.scala 27:20]
  reg [1:0] pht_426; // @[BPU.scala 27:20]
  reg [1:0] pht_427; // @[BPU.scala 27:20]
  reg [1:0] pht_428; // @[BPU.scala 27:20]
  reg [1:0] pht_429; // @[BPU.scala 27:20]
  reg [1:0] pht_430; // @[BPU.scala 27:20]
  reg [1:0] pht_431; // @[BPU.scala 27:20]
  reg [1:0] pht_432; // @[BPU.scala 27:20]
  reg [1:0] pht_433; // @[BPU.scala 27:20]
  reg [1:0] pht_434; // @[BPU.scala 27:20]
  reg [1:0] pht_435; // @[BPU.scala 27:20]
  reg [1:0] pht_436; // @[BPU.scala 27:20]
  reg [1:0] pht_437; // @[BPU.scala 27:20]
  reg [1:0] pht_438; // @[BPU.scala 27:20]
  reg [1:0] pht_439; // @[BPU.scala 27:20]
  reg [1:0] pht_440; // @[BPU.scala 27:20]
  reg [1:0] pht_441; // @[BPU.scala 27:20]
  reg [1:0] pht_442; // @[BPU.scala 27:20]
  reg [1:0] pht_443; // @[BPU.scala 27:20]
  reg [1:0] pht_444; // @[BPU.scala 27:20]
  reg [1:0] pht_445; // @[BPU.scala 27:20]
  reg [1:0] pht_446; // @[BPU.scala 27:20]
  reg [1:0] pht_447; // @[BPU.scala 27:20]
  reg [1:0] pht_448; // @[BPU.scala 27:20]
  reg [1:0] pht_449; // @[BPU.scala 27:20]
  reg [1:0] pht_450; // @[BPU.scala 27:20]
  reg [1:0] pht_451; // @[BPU.scala 27:20]
  reg [1:0] pht_452; // @[BPU.scala 27:20]
  reg [1:0] pht_453; // @[BPU.scala 27:20]
  reg [1:0] pht_454; // @[BPU.scala 27:20]
  reg [1:0] pht_455; // @[BPU.scala 27:20]
  reg [1:0] pht_456; // @[BPU.scala 27:20]
  reg [1:0] pht_457; // @[BPU.scala 27:20]
  reg [1:0] pht_458; // @[BPU.scala 27:20]
  reg [1:0] pht_459; // @[BPU.scala 27:20]
  reg [1:0] pht_460; // @[BPU.scala 27:20]
  reg [1:0] pht_461; // @[BPU.scala 27:20]
  reg [1:0] pht_462; // @[BPU.scala 27:20]
  reg [1:0] pht_463; // @[BPU.scala 27:20]
  reg [1:0] pht_464; // @[BPU.scala 27:20]
  reg [1:0] pht_465; // @[BPU.scala 27:20]
  reg [1:0] pht_466; // @[BPU.scala 27:20]
  reg [1:0] pht_467; // @[BPU.scala 27:20]
  reg [1:0] pht_468; // @[BPU.scala 27:20]
  reg [1:0] pht_469; // @[BPU.scala 27:20]
  reg [1:0] pht_470; // @[BPU.scala 27:20]
  reg [1:0] pht_471; // @[BPU.scala 27:20]
  reg [1:0] pht_472; // @[BPU.scala 27:20]
  reg [1:0] pht_473; // @[BPU.scala 27:20]
  reg [1:0] pht_474; // @[BPU.scala 27:20]
  reg [1:0] pht_475; // @[BPU.scala 27:20]
  reg [1:0] pht_476; // @[BPU.scala 27:20]
  reg [1:0] pht_477; // @[BPU.scala 27:20]
  reg [1:0] pht_478; // @[BPU.scala 27:20]
  reg [1:0] pht_479; // @[BPU.scala 27:20]
  reg [1:0] pht_480; // @[BPU.scala 27:20]
  reg [1:0] pht_481; // @[BPU.scala 27:20]
  reg [1:0] pht_482; // @[BPU.scala 27:20]
  reg [1:0] pht_483; // @[BPU.scala 27:20]
  reg [1:0] pht_484; // @[BPU.scala 27:20]
  reg [1:0] pht_485; // @[BPU.scala 27:20]
  reg [1:0] pht_486; // @[BPU.scala 27:20]
  reg [1:0] pht_487; // @[BPU.scala 27:20]
  reg [1:0] pht_488; // @[BPU.scala 27:20]
  reg [1:0] pht_489; // @[BPU.scala 27:20]
  reg [1:0] pht_490; // @[BPU.scala 27:20]
  reg [1:0] pht_491; // @[BPU.scala 27:20]
  reg [1:0] pht_492; // @[BPU.scala 27:20]
  reg [1:0] pht_493; // @[BPU.scala 27:20]
  reg [1:0] pht_494; // @[BPU.scala 27:20]
  reg [1:0] pht_495; // @[BPU.scala 27:20]
  reg [1:0] pht_496; // @[BPU.scala 27:20]
  reg [1:0] pht_497; // @[BPU.scala 27:20]
  reg [1:0] pht_498; // @[BPU.scala 27:20]
  reg [1:0] pht_499; // @[BPU.scala 27:20]
  reg [1:0] pht_500; // @[BPU.scala 27:20]
  reg [1:0] pht_501; // @[BPU.scala 27:20]
  reg [1:0] pht_502; // @[BPU.scala 27:20]
  reg [1:0] pht_503; // @[BPU.scala 27:20]
  reg [1:0] pht_504; // @[BPU.scala 27:20]
  reg [1:0] pht_505; // @[BPU.scala 27:20]
  reg [1:0] pht_506; // @[BPU.scala 27:20]
  reg [1:0] pht_507; // @[BPU.scala 27:20]
  reg [1:0] pht_508; // @[BPU.scala 27:20]
  reg [1:0] pht_509; // @[BPU.scala 27:20]
  reg [1:0] pht_510; // @[BPU.scala 27:20]
  reg [1:0] pht_511; // @[BPU.scala 27:20]
  reg [36:0] btb_0_tag; // @[BPU.scala 28:20]
  reg [36:0] btb_0_target; // @[BPU.scala 28:20]
  reg  btb_0_valid; // @[BPU.scala 28:20]
  reg [36:0] btb_1_tag; // @[BPU.scala 28:20]
  reg [36:0] btb_1_target; // @[BPU.scala 28:20]
  reg  btb_1_valid; // @[BPU.scala 28:20]
  reg [36:0] btb_2_tag; // @[BPU.scala 28:20]
  reg [36:0] btb_2_target; // @[BPU.scala 28:20]
  reg  btb_2_valid; // @[BPU.scala 28:20]
  reg [36:0] btb_3_tag; // @[BPU.scala 28:20]
  reg [36:0] btb_3_target; // @[BPU.scala 28:20]
  reg  btb_3_valid; // @[BPU.scala 28:20]
  reg [36:0] btb_4_tag; // @[BPU.scala 28:20]
  reg [36:0] btb_4_target; // @[BPU.scala 28:20]
  reg  btb_4_valid; // @[BPU.scala 28:20]
  reg [36:0] btb_5_tag; // @[BPU.scala 28:20]
  reg [36:0] btb_5_target; // @[BPU.scala 28:20]
  reg  btb_5_valid; // @[BPU.scala 28:20]
  reg [36:0] btb_6_tag; // @[BPU.scala 28:20]
  reg [36:0] btb_6_target; // @[BPU.scala 28:20]
  reg  btb_6_valid; // @[BPU.scala 28:20]
  reg [36:0] btb_7_tag; // @[BPU.scala 28:20]
  reg [36:0] btb_7_target; // @[BPU.scala 28:20]
  reg  btb_7_valid; // @[BPU.scala 28:20]
  reg [36:0] btb_8_tag; // @[BPU.scala 28:20]
  reg [36:0] btb_8_target; // @[BPU.scala 28:20]
  reg  btb_8_valid; // @[BPU.scala 28:20]
  reg [36:0] btb_9_tag; // @[BPU.scala 28:20]
  reg [36:0] btb_9_target; // @[BPU.scala 28:20]
  reg  btb_9_valid; // @[BPU.scala 28:20]
  reg [36:0] btb_10_tag; // @[BPU.scala 28:20]
  reg [36:0] btb_10_target; // @[BPU.scala 28:20]
  reg  btb_10_valid; // @[BPU.scala 28:20]
  reg [36:0] btb_11_tag; // @[BPU.scala 28:20]
  reg [36:0] btb_11_target; // @[BPU.scala 28:20]
  reg  btb_11_valid; // @[BPU.scala 28:20]
  reg [36:0] btb_12_tag; // @[BPU.scala 28:20]
  reg [36:0] btb_12_target; // @[BPU.scala 28:20]
  reg  btb_12_valid; // @[BPU.scala 28:20]
  reg [36:0] btb_13_tag; // @[BPU.scala 28:20]
  reg [36:0] btb_13_target; // @[BPU.scala 28:20]
  reg  btb_13_valid; // @[BPU.scala 28:20]
  reg [36:0] btb_14_tag; // @[BPU.scala 28:20]
  reg [36:0] btb_14_target; // @[BPU.scala 28:20]
  reg  btb_14_valid; // @[BPU.scala 28:20]
  reg [36:0] btb_15_tag; // @[BPU.scala 28:20]
  reg [36:0] btb_15_target; // @[BPU.scala 28:20]
  reg  btb_15_valid; // @[BPU.scala 28:20]
  wire [8:0] pht_ridx = io_pc[10:2] ^ ghr; // @[BPU.scala 31:40]
  wire [1:0] _GEN_1 = 9'h1 == pht_ridx ? pht_1 : pht_0; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_2 = 9'h2 == pht_ridx ? pht_2 : _GEN_1; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_3 = 9'h3 == pht_ridx ? pht_3 : _GEN_2; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_4 = 9'h4 == pht_ridx ? pht_4 : _GEN_3; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_5 = 9'h5 == pht_ridx ? pht_5 : _GEN_4; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_6 = 9'h6 == pht_ridx ? pht_6 : _GEN_5; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_7 = 9'h7 == pht_ridx ? pht_7 : _GEN_6; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_8 = 9'h8 == pht_ridx ? pht_8 : _GEN_7; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_9 = 9'h9 == pht_ridx ? pht_9 : _GEN_8; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_10 = 9'ha == pht_ridx ? pht_10 : _GEN_9; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_11 = 9'hb == pht_ridx ? pht_11 : _GEN_10; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_12 = 9'hc == pht_ridx ? pht_12 : _GEN_11; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_13 = 9'hd == pht_ridx ? pht_13 : _GEN_12; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_14 = 9'he == pht_ridx ? pht_14 : _GEN_13; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_15 = 9'hf == pht_ridx ? pht_15 : _GEN_14; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_16 = 9'h10 == pht_ridx ? pht_16 : _GEN_15; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_17 = 9'h11 == pht_ridx ? pht_17 : _GEN_16; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_18 = 9'h12 == pht_ridx ? pht_18 : _GEN_17; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_19 = 9'h13 == pht_ridx ? pht_19 : _GEN_18; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_20 = 9'h14 == pht_ridx ? pht_20 : _GEN_19; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_21 = 9'h15 == pht_ridx ? pht_21 : _GEN_20; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_22 = 9'h16 == pht_ridx ? pht_22 : _GEN_21; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_23 = 9'h17 == pht_ridx ? pht_23 : _GEN_22; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_24 = 9'h18 == pht_ridx ? pht_24 : _GEN_23; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_25 = 9'h19 == pht_ridx ? pht_25 : _GEN_24; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_26 = 9'h1a == pht_ridx ? pht_26 : _GEN_25; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_27 = 9'h1b == pht_ridx ? pht_27 : _GEN_26; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_28 = 9'h1c == pht_ridx ? pht_28 : _GEN_27; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_29 = 9'h1d == pht_ridx ? pht_29 : _GEN_28; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_30 = 9'h1e == pht_ridx ? pht_30 : _GEN_29; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_31 = 9'h1f == pht_ridx ? pht_31 : _GEN_30; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_32 = 9'h20 == pht_ridx ? pht_32 : _GEN_31; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_33 = 9'h21 == pht_ridx ? pht_33 : _GEN_32; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_34 = 9'h22 == pht_ridx ? pht_34 : _GEN_33; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_35 = 9'h23 == pht_ridx ? pht_35 : _GEN_34; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_36 = 9'h24 == pht_ridx ? pht_36 : _GEN_35; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_37 = 9'h25 == pht_ridx ? pht_37 : _GEN_36; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_38 = 9'h26 == pht_ridx ? pht_38 : _GEN_37; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_39 = 9'h27 == pht_ridx ? pht_39 : _GEN_38; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_40 = 9'h28 == pht_ridx ? pht_40 : _GEN_39; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_41 = 9'h29 == pht_ridx ? pht_41 : _GEN_40; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_42 = 9'h2a == pht_ridx ? pht_42 : _GEN_41; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_43 = 9'h2b == pht_ridx ? pht_43 : _GEN_42; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_44 = 9'h2c == pht_ridx ? pht_44 : _GEN_43; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_45 = 9'h2d == pht_ridx ? pht_45 : _GEN_44; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_46 = 9'h2e == pht_ridx ? pht_46 : _GEN_45; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_47 = 9'h2f == pht_ridx ? pht_47 : _GEN_46; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_48 = 9'h30 == pht_ridx ? pht_48 : _GEN_47; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_49 = 9'h31 == pht_ridx ? pht_49 : _GEN_48; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_50 = 9'h32 == pht_ridx ? pht_50 : _GEN_49; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_51 = 9'h33 == pht_ridx ? pht_51 : _GEN_50; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_52 = 9'h34 == pht_ridx ? pht_52 : _GEN_51; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_53 = 9'h35 == pht_ridx ? pht_53 : _GEN_52; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_54 = 9'h36 == pht_ridx ? pht_54 : _GEN_53; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_55 = 9'h37 == pht_ridx ? pht_55 : _GEN_54; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_56 = 9'h38 == pht_ridx ? pht_56 : _GEN_55; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_57 = 9'h39 == pht_ridx ? pht_57 : _GEN_56; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_58 = 9'h3a == pht_ridx ? pht_58 : _GEN_57; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_59 = 9'h3b == pht_ridx ? pht_59 : _GEN_58; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_60 = 9'h3c == pht_ridx ? pht_60 : _GEN_59; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_61 = 9'h3d == pht_ridx ? pht_61 : _GEN_60; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_62 = 9'h3e == pht_ridx ? pht_62 : _GEN_61; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_63 = 9'h3f == pht_ridx ? pht_63 : _GEN_62; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_64 = 9'h40 == pht_ridx ? pht_64 : _GEN_63; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_65 = 9'h41 == pht_ridx ? pht_65 : _GEN_64; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_66 = 9'h42 == pht_ridx ? pht_66 : _GEN_65; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_67 = 9'h43 == pht_ridx ? pht_67 : _GEN_66; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_68 = 9'h44 == pht_ridx ? pht_68 : _GEN_67; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_69 = 9'h45 == pht_ridx ? pht_69 : _GEN_68; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_70 = 9'h46 == pht_ridx ? pht_70 : _GEN_69; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_71 = 9'h47 == pht_ridx ? pht_71 : _GEN_70; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_72 = 9'h48 == pht_ridx ? pht_72 : _GEN_71; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_73 = 9'h49 == pht_ridx ? pht_73 : _GEN_72; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_74 = 9'h4a == pht_ridx ? pht_74 : _GEN_73; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_75 = 9'h4b == pht_ridx ? pht_75 : _GEN_74; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_76 = 9'h4c == pht_ridx ? pht_76 : _GEN_75; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_77 = 9'h4d == pht_ridx ? pht_77 : _GEN_76; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_78 = 9'h4e == pht_ridx ? pht_78 : _GEN_77; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_79 = 9'h4f == pht_ridx ? pht_79 : _GEN_78; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_80 = 9'h50 == pht_ridx ? pht_80 : _GEN_79; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_81 = 9'h51 == pht_ridx ? pht_81 : _GEN_80; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_82 = 9'h52 == pht_ridx ? pht_82 : _GEN_81; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_83 = 9'h53 == pht_ridx ? pht_83 : _GEN_82; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_84 = 9'h54 == pht_ridx ? pht_84 : _GEN_83; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_85 = 9'h55 == pht_ridx ? pht_85 : _GEN_84; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_86 = 9'h56 == pht_ridx ? pht_86 : _GEN_85; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_87 = 9'h57 == pht_ridx ? pht_87 : _GEN_86; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_88 = 9'h58 == pht_ridx ? pht_88 : _GEN_87; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_89 = 9'h59 == pht_ridx ? pht_89 : _GEN_88; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_90 = 9'h5a == pht_ridx ? pht_90 : _GEN_89; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_91 = 9'h5b == pht_ridx ? pht_91 : _GEN_90; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_92 = 9'h5c == pht_ridx ? pht_92 : _GEN_91; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_93 = 9'h5d == pht_ridx ? pht_93 : _GEN_92; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_94 = 9'h5e == pht_ridx ? pht_94 : _GEN_93; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_95 = 9'h5f == pht_ridx ? pht_95 : _GEN_94; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_96 = 9'h60 == pht_ridx ? pht_96 : _GEN_95; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_97 = 9'h61 == pht_ridx ? pht_97 : _GEN_96; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_98 = 9'h62 == pht_ridx ? pht_98 : _GEN_97; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_99 = 9'h63 == pht_ridx ? pht_99 : _GEN_98; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_100 = 9'h64 == pht_ridx ? pht_100 : _GEN_99; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_101 = 9'h65 == pht_ridx ? pht_101 : _GEN_100; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_102 = 9'h66 == pht_ridx ? pht_102 : _GEN_101; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_103 = 9'h67 == pht_ridx ? pht_103 : _GEN_102; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_104 = 9'h68 == pht_ridx ? pht_104 : _GEN_103; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_105 = 9'h69 == pht_ridx ? pht_105 : _GEN_104; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_106 = 9'h6a == pht_ridx ? pht_106 : _GEN_105; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_107 = 9'h6b == pht_ridx ? pht_107 : _GEN_106; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_108 = 9'h6c == pht_ridx ? pht_108 : _GEN_107; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_109 = 9'h6d == pht_ridx ? pht_109 : _GEN_108; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_110 = 9'h6e == pht_ridx ? pht_110 : _GEN_109; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_111 = 9'h6f == pht_ridx ? pht_111 : _GEN_110; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_112 = 9'h70 == pht_ridx ? pht_112 : _GEN_111; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_113 = 9'h71 == pht_ridx ? pht_113 : _GEN_112; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_114 = 9'h72 == pht_ridx ? pht_114 : _GEN_113; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_115 = 9'h73 == pht_ridx ? pht_115 : _GEN_114; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_116 = 9'h74 == pht_ridx ? pht_116 : _GEN_115; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_117 = 9'h75 == pht_ridx ? pht_117 : _GEN_116; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_118 = 9'h76 == pht_ridx ? pht_118 : _GEN_117; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_119 = 9'h77 == pht_ridx ? pht_119 : _GEN_118; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_120 = 9'h78 == pht_ridx ? pht_120 : _GEN_119; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_121 = 9'h79 == pht_ridx ? pht_121 : _GEN_120; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_122 = 9'h7a == pht_ridx ? pht_122 : _GEN_121; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_123 = 9'h7b == pht_ridx ? pht_123 : _GEN_122; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_124 = 9'h7c == pht_ridx ? pht_124 : _GEN_123; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_125 = 9'h7d == pht_ridx ? pht_125 : _GEN_124; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_126 = 9'h7e == pht_ridx ? pht_126 : _GEN_125; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_127 = 9'h7f == pht_ridx ? pht_127 : _GEN_126; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_128 = 9'h80 == pht_ridx ? pht_128 : _GEN_127; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_129 = 9'h81 == pht_ridx ? pht_129 : _GEN_128; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_130 = 9'h82 == pht_ridx ? pht_130 : _GEN_129; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_131 = 9'h83 == pht_ridx ? pht_131 : _GEN_130; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_132 = 9'h84 == pht_ridx ? pht_132 : _GEN_131; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_133 = 9'h85 == pht_ridx ? pht_133 : _GEN_132; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_134 = 9'h86 == pht_ridx ? pht_134 : _GEN_133; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_135 = 9'h87 == pht_ridx ? pht_135 : _GEN_134; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_136 = 9'h88 == pht_ridx ? pht_136 : _GEN_135; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_137 = 9'h89 == pht_ridx ? pht_137 : _GEN_136; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_138 = 9'h8a == pht_ridx ? pht_138 : _GEN_137; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_139 = 9'h8b == pht_ridx ? pht_139 : _GEN_138; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_140 = 9'h8c == pht_ridx ? pht_140 : _GEN_139; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_141 = 9'h8d == pht_ridx ? pht_141 : _GEN_140; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_142 = 9'h8e == pht_ridx ? pht_142 : _GEN_141; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_143 = 9'h8f == pht_ridx ? pht_143 : _GEN_142; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_144 = 9'h90 == pht_ridx ? pht_144 : _GEN_143; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_145 = 9'h91 == pht_ridx ? pht_145 : _GEN_144; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_146 = 9'h92 == pht_ridx ? pht_146 : _GEN_145; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_147 = 9'h93 == pht_ridx ? pht_147 : _GEN_146; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_148 = 9'h94 == pht_ridx ? pht_148 : _GEN_147; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_149 = 9'h95 == pht_ridx ? pht_149 : _GEN_148; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_150 = 9'h96 == pht_ridx ? pht_150 : _GEN_149; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_151 = 9'h97 == pht_ridx ? pht_151 : _GEN_150; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_152 = 9'h98 == pht_ridx ? pht_152 : _GEN_151; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_153 = 9'h99 == pht_ridx ? pht_153 : _GEN_152; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_154 = 9'h9a == pht_ridx ? pht_154 : _GEN_153; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_155 = 9'h9b == pht_ridx ? pht_155 : _GEN_154; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_156 = 9'h9c == pht_ridx ? pht_156 : _GEN_155; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_157 = 9'h9d == pht_ridx ? pht_157 : _GEN_156; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_158 = 9'h9e == pht_ridx ? pht_158 : _GEN_157; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_159 = 9'h9f == pht_ridx ? pht_159 : _GEN_158; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_160 = 9'ha0 == pht_ridx ? pht_160 : _GEN_159; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_161 = 9'ha1 == pht_ridx ? pht_161 : _GEN_160; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_162 = 9'ha2 == pht_ridx ? pht_162 : _GEN_161; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_163 = 9'ha3 == pht_ridx ? pht_163 : _GEN_162; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_164 = 9'ha4 == pht_ridx ? pht_164 : _GEN_163; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_165 = 9'ha5 == pht_ridx ? pht_165 : _GEN_164; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_166 = 9'ha6 == pht_ridx ? pht_166 : _GEN_165; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_167 = 9'ha7 == pht_ridx ? pht_167 : _GEN_166; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_168 = 9'ha8 == pht_ridx ? pht_168 : _GEN_167; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_169 = 9'ha9 == pht_ridx ? pht_169 : _GEN_168; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_170 = 9'haa == pht_ridx ? pht_170 : _GEN_169; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_171 = 9'hab == pht_ridx ? pht_171 : _GEN_170; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_172 = 9'hac == pht_ridx ? pht_172 : _GEN_171; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_173 = 9'had == pht_ridx ? pht_173 : _GEN_172; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_174 = 9'hae == pht_ridx ? pht_174 : _GEN_173; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_175 = 9'haf == pht_ridx ? pht_175 : _GEN_174; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_176 = 9'hb0 == pht_ridx ? pht_176 : _GEN_175; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_177 = 9'hb1 == pht_ridx ? pht_177 : _GEN_176; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_178 = 9'hb2 == pht_ridx ? pht_178 : _GEN_177; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_179 = 9'hb3 == pht_ridx ? pht_179 : _GEN_178; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_180 = 9'hb4 == pht_ridx ? pht_180 : _GEN_179; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_181 = 9'hb5 == pht_ridx ? pht_181 : _GEN_180; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_182 = 9'hb6 == pht_ridx ? pht_182 : _GEN_181; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_183 = 9'hb7 == pht_ridx ? pht_183 : _GEN_182; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_184 = 9'hb8 == pht_ridx ? pht_184 : _GEN_183; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_185 = 9'hb9 == pht_ridx ? pht_185 : _GEN_184; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_186 = 9'hba == pht_ridx ? pht_186 : _GEN_185; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_187 = 9'hbb == pht_ridx ? pht_187 : _GEN_186; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_188 = 9'hbc == pht_ridx ? pht_188 : _GEN_187; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_189 = 9'hbd == pht_ridx ? pht_189 : _GEN_188; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_190 = 9'hbe == pht_ridx ? pht_190 : _GEN_189; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_191 = 9'hbf == pht_ridx ? pht_191 : _GEN_190; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_192 = 9'hc0 == pht_ridx ? pht_192 : _GEN_191; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_193 = 9'hc1 == pht_ridx ? pht_193 : _GEN_192; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_194 = 9'hc2 == pht_ridx ? pht_194 : _GEN_193; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_195 = 9'hc3 == pht_ridx ? pht_195 : _GEN_194; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_196 = 9'hc4 == pht_ridx ? pht_196 : _GEN_195; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_197 = 9'hc5 == pht_ridx ? pht_197 : _GEN_196; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_198 = 9'hc6 == pht_ridx ? pht_198 : _GEN_197; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_199 = 9'hc7 == pht_ridx ? pht_199 : _GEN_198; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_200 = 9'hc8 == pht_ridx ? pht_200 : _GEN_199; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_201 = 9'hc9 == pht_ridx ? pht_201 : _GEN_200; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_202 = 9'hca == pht_ridx ? pht_202 : _GEN_201; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_203 = 9'hcb == pht_ridx ? pht_203 : _GEN_202; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_204 = 9'hcc == pht_ridx ? pht_204 : _GEN_203; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_205 = 9'hcd == pht_ridx ? pht_205 : _GEN_204; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_206 = 9'hce == pht_ridx ? pht_206 : _GEN_205; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_207 = 9'hcf == pht_ridx ? pht_207 : _GEN_206; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_208 = 9'hd0 == pht_ridx ? pht_208 : _GEN_207; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_209 = 9'hd1 == pht_ridx ? pht_209 : _GEN_208; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_210 = 9'hd2 == pht_ridx ? pht_210 : _GEN_209; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_211 = 9'hd3 == pht_ridx ? pht_211 : _GEN_210; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_212 = 9'hd4 == pht_ridx ? pht_212 : _GEN_211; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_213 = 9'hd5 == pht_ridx ? pht_213 : _GEN_212; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_214 = 9'hd6 == pht_ridx ? pht_214 : _GEN_213; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_215 = 9'hd7 == pht_ridx ? pht_215 : _GEN_214; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_216 = 9'hd8 == pht_ridx ? pht_216 : _GEN_215; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_217 = 9'hd9 == pht_ridx ? pht_217 : _GEN_216; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_218 = 9'hda == pht_ridx ? pht_218 : _GEN_217; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_219 = 9'hdb == pht_ridx ? pht_219 : _GEN_218; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_220 = 9'hdc == pht_ridx ? pht_220 : _GEN_219; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_221 = 9'hdd == pht_ridx ? pht_221 : _GEN_220; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_222 = 9'hde == pht_ridx ? pht_222 : _GEN_221; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_223 = 9'hdf == pht_ridx ? pht_223 : _GEN_222; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_224 = 9'he0 == pht_ridx ? pht_224 : _GEN_223; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_225 = 9'he1 == pht_ridx ? pht_225 : _GEN_224; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_226 = 9'he2 == pht_ridx ? pht_226 : _GEN_225; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_227 = 9'he3 == pht_ridx ? pht_227 : _GEN_226; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_228 = 9'he4 == pht_ridx ? pht_228 : _GEN_227; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_229 = 9'he5 == pht_ridx ? pht_229 : _GEN_228; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_230 = 9'he6 == pht_ridx ? pht_230 : _GEN_229; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_231 = 9'he7 == pht_ridx ? pht_231 : _GEN_230; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_232 = 9'he8 == pht_ridx ? pht_232 : _GEN_231; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_233 = 9'he9 == pht_ridx ? pht_233 : _GEN_232; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_234 = 9'hea == pht_ridx ? pht_234 : _GEN_233; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_235 = 9'heb == pht_ridx ? pht_235 : _GEN_234; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_236 = 9'hec == pht_ridx ? pht_236 : _GEN_235; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_237 = 9'hed == pht_ridx ? pht_237 : _GEN_236; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_238 = 9'hee == pht_ridx ? pht_238 : _GEN_237; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_239 = 9'hef == pht_ridx ? pht_239 : _GEN_238; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_240 = 9'hf0 == pht_ridx ? pht_240 : _GEN_239; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_241 = 9'hf1 == pht_ridx ? pht_241 : _GEN_240; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_242 = 9'hf2 == pht_ridx ? pht_242 : _GEN_241; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_243 = 9'hf3 == pht_ridx ? pht_243 : _GEN_242; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_244 = 9'hf4 == pht_ridx ? pht_244 : _GEN_243; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_245 = 9'hf5 == pht_ridx ? pht_245 : _GEN_244; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_246 = 9'hf6 == pht_ridx ? pht_246 : _GEN_245; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_247 = 9'hf7 == pht_ridx ? pht_247 : _GEN_246; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_248 = 9'hf8 == pht_ridx ? pht_248 : _GEN_247; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_249 = 9'hf9 == pht_ridx ? pht_249 : _GEN_248; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_250 = 9'hfa == pht_ridx ? pht_250 : _GEN_249; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_251 = 9'hfb == pht_ridx ? pht_251 : _GEN_250; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_252 = 9'hfc == pht_ridx ? pht_252 : _GEN_251; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_253 = 9'hfd == pht_ridx ? pht_253 : _GEN_252; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_254 = 9'hfe == pht_ridx ? pht_254 : _GEN_253; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_255 = 9'hff == pht_ridx ? pht_255 : _GEN_254; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_256 = 9'h100 == pht_ridx ? pht_256 : _GEN_255; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_257 = 9'h101 == pht_ridx ? pht_257 : _GEN_256; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_258 = 9'h102 == pht_ridx ? pht_258 : _GEN_257; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_259 = 9'h103 == pht_ridx ? pht_259 : _GEN_258; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_260 = 9'h104 == pht_ridx ? pht_260 : _GEN_259; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_261 = 9'h105 == pht_ridx ? pht_261 : _GEN_260; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_262 = 9'h106 == pht_ridx ? pht_262 : _GEN_261; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_263 = 9'h107 == pht_ridx ? pht_263 : _GEN_262; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_264 = 9'h108 == pht_ridx ? pht_264 : _GEN_263; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_265 = 9'h109 == pht_ridx ? pht_265 : _GEN_264; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_266 = 9'h10a == pht_ridx ? pht_266 : _GEN_265; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_267 = 9'h10b == pht_ridx ? pht_267 : _GEN_266; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_268 = 9'h10c == pht_ridx ? pht_268 : _GEN_267; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_269 = 9'h10d == pht_ridx ? pht_269 : _GEN_268; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_270 = 9'h10e == pht_ridx ? pht_270 : _GEN_269; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_271 = 9'h10f == pht_ridx ? pht_271 : _GEN_270; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_272 = 9'h110 == pht_ridx ? pht_272 : _GEN_271; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_273 = 9'h111 == pht_ridx ? pht_273 : _GEN_272; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_274 = 9'h112 == pht_ridx ? pht_274 : _GEN_273; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_275 = 9'h113 == pht_ridx ? pht_275 : _GEN_274; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_276 = 9'h114 == pht_ridx ? pht_276 : _GEN_275; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_277 = 9'h115 == pht_ridx ? pht_277 : _GEN_276; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_278 = 9'h116 == pht_ridx ? pht_278 : _GEN_277; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_279 = 9'h117 == pht_ridx ? pht_279 : _GEN_278; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_280 = 9'h118 == pht_ridx ? pht_280 : _GEN_279; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_281 = 9'h119 == pht_ridx ? pht_281 : _GEN_280; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_282 = 9'h11a == pht_ridx ? pht_282 : _GEN_281; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_283 = 9'h11b == pht_ridx ? pht_283 : _GEN_282; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_284 = 9'h11c == pht_ridx ? pht_284 : _GEN_283; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_285 = 9'h11d == pht_ridx ? pht_285 : _GEN_284; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_286 = 9'h11e == pht_ridx ? pht_286 : _GEN_285; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_287 = 9'h11f == pht_ridx ? pht_287 : _GEN_286; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_288 = 9'h120 == pht_ridx ? pht_288 : _GEN_287; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_289 = 9'h121 == pht_ridx ? pht_289 : _GEN_288; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_290 = 9'h122 == pht_ridx ? pht_290 : _GEN_289; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_291 = 9'h123 == pht_ridx ? pht_291 : _GEN_290; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_292 = 9'h124 == pht_ridx ? pht_292 : _GEN_291; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_293 = 9'h125 == pht_ridx ? pht_293 : _GEN_292; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_294 = 9'h126 == pht_ridx ? pht_294 : _GEN_293; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_295 = 9'h127 == pht_ridx ? pht_295 : _GEN_294; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_296 = 9'h128 == pht_ridx ? pht_296 : _GEN_295; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_297 = 9'h129 == pht_ridx ? pht_297 : _GEN_296; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_298 = 9'h12a == pht_ridx ? pht_298 : _GEN_297; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_299 = 9'h12b == pht_ridx ? pht_299 : _GEN_298; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_300 = 9'h12c == pht_ridx ? pht_300 : _GEN_299; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_301 = 9'h12d == pht_ridx ? pht_301 : _GEN_300; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_302 = 9'h12e == pht_ridx ? pht_302 : _GEN_301; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_303 = 9'h12f == pht_ridx ? pht_303 : _GEN_302; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_304 = 9'h130 == pht_ridx ? pht_304 : _GEN_303; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_305 = 9'h131 == pht_ridx ? pht_305 : _GEN_304; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_306 = 9'h132 == pht_ridx ? pht_306 : _GEN_305; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_307 = 9'h133 == pht_ridx ? pht_307 : _GEN_306; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_308 = 9'h134 == pht_ridx ? pht_308 : _GEN_307; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_309 = 9'h135 == pht_ridx ? pht_309 : _GEN_308; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_310 = 9'h136 == pht_ridx ? pht_310 : _GEN_309; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_311 = 9'h137 == pht_ridx ? pht_311 : _GEN_310; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_312 = 9'h138 == pht_ridx ? pht_312 : _GEN_311; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_313 = 9'h139 == pht_ridx ? pht_313 : _GEN_312; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_314 = 9'h13a == pht_ridx ? pht_314 : _GEN_313; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_315 = 9'h13b == pht_ridx ? pht_315 : _GEN_314; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_316 = 9'h13c == pht_ridx ? pht_316 : _GEN_315; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_317 = 9'h13d == pht_ridx ? pht_317 : _GEN_316; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_318 = 9'h13e == pht_ridx ? pht_318 : _GEN_317; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_319 = 9'h13f == pht_ridx ? pht_319 : _GEN_318; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_320 = 9'h140 == pht_ridx ? pht_320 : _GEN_319; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_321 = 9'h141 == pht_ridx ? pht_321 : _GEN_320; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_322 = 9'h142 == pht_ridx ? pht_322 : _GEN_321; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_323 = 9'h143 == pht_ridx ? pht_323 : _GEN_322; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_324 = 9'h144 == pht_ridx ? pht_324 : _GEN_323; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_325 = 9'h145 == pht_ridx ? pht_325 : _GEN_324; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_326 = 9'h146 == pht_ridx ? pht_326 : _GEN_325; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_327 = 9'h147 == pht_ridx ? pht_327 : _GEN_326; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_328 = 9'h148 == pht_ridx ? pht_328 : _GEN_327; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_329 = 9'h149 == pht_ridx ? pht_329 : _GEN_328; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_330 = 9'h14a == pht_ridx ? pht_330 : _GEN_329; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_331 = 9'h14b == pht_ridx ? pht_331 : _GEN_330; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_332 = 9'h14c == pht_ridx ? pht_332 : _GEN_331; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_333 = 9'h14d == pht_ridx ? pht_333 : _GEN_332; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_334 = 9'h14e == pht_ridx ? pht_334 : _GEN_333; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_335 = 9'h14f == pht_ridx ? pht_335 : _GEN_334; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_336 = 9'h150 == pht_ridx ? pht_336 : _GEN_335; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_337 = 9'h151 == pht_ridx ? pht_337 : _GEN_336; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_338 = 9'h152 == pht_ridx ? pht_338 : _GEN_337; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_339 = 9'h153 == pht_ridx ? pht_339 : _GEN_338; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_340 = 9'h154 == pht_ridx ? pht_340 : _GEN_339; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_341 = 9'h155 == pht_ridx ? pht_341 : _GEN_340; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_342 = 9'h156 == pht_ridx ? pht_342 : _GEN_341; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_343 = 9'h157 == pht_ridx ? pht_343 : _GEN_342; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_344 = 9'h158 == pht_ridx ? pht_344 : _GEN_343; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_345 = 9'h159 == pht_ridx ? pht_345 : _GEN_344; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_346 = 9'h15a == pht_ridx ? pht_346 : _GEN_345; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_347 = 9'h15b == pht_ridx ? pht_347 : _GEN_346; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_348 = 9'h15c == pht_ridx ? pht_348 : _GEN_347; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_349 = 9'h15d == pht_ridx ? pht_349 : _GEN_348; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_350 = 9'h15e == pht_ridx ? pht_350 : _GEN_349; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_351 = 9'h15f == pht_ridx ? pht_351 : _GEN_350; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_352 = 9'h160 == pht_ridx ? pht_352 : _GEN_351; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_353 = 9'h161 == pht_ridx ? pht_353 : _GEN_352; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_354 = 9'h162 == pht_ridx ? pht_354 : _GEN_353; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_355 = 9'h163 == pht_ridx ? pht_355 : _GEN_354; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_356 = 9'h164 == pht_ridx ? pht_356 : _GEN_355; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_357 = 9'h165 == pht_ridx ? pht_357 : _GEN_356; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_358 = 9'h166 == pht_ridx ? pht_358 : _GEN_357; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_359 = 9'h167 == pht_ridx ? pht_359 : _GEN_358; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_360 = 9'h168 == pht_ridx ? pht_360 : _GEN_359; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_361 = 9'h169 == pht_ridx ? pht_361 : _GEN_360; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_362 = 9'h16a == pht_ridx ? pht_362 : _GEN_361; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_363 = 9'h16b == pht_ridx ? pht_363 : _GEN_362; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_364 = 9'h16c == pht_ridx ? pht_364 : _GEN_363; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_365 = 9'h16d == pht_ridx ? pht_365 : _GEN_364; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_366 = 9'h16e == pht_ridx ? pht_366 : _GEN_365; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_367 = 9'h16f == pht_ridx ? pht_367 : _GEN_366; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_368 = 9'h170 == pht_ridx ? pht_368 : _GEN_367; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_369 = 9'h171 == pht_ridx ? pht_369 : _GEN_368; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_370 = 9'h172 == pht_ridx ? pht_370 : _GEN_369; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_371 = 9'h173 == pht_ridx ? pht_371 : _GEN_370; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_372 = 9'h174 == pht_ridx ? pht_372 : _GEN_371; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_373 = 9'h175 == pht_ridx ? pht_373 : _GEN_372; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_374 = 9'h176 == pht_ridx ? pht_374 : _GEN_373; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_375 = 9'h177 == pht_ridx ? pht_375 : _GEN_374; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_376 = 9'h178 == pht_ridx ? pht_376 : _GEN_375; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_377 = 9'h179 == pht_ridx ? pht_377 : _GEN_376; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_378 = 9'h17a == pht_ridx ? pht_378 : _GEN_377; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_379 = 9'h17b == pht_ridx ? pht_379 : _GEN_378; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_380 = 9'h17c == pht_ridx ? pht_380 : _GEN_379; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_381 = 9'h17d == pht_ridx ? pht_381 : _GEN_380; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_382 = 9'h17e == pht_ridx ? pht_382 : _GEN_381; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_383 = 9'h17f == pht_ridx ? pht_383 : _GEN_382; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_384 = 9'h180 == pht_ridx ? pht_384 : _GEN_383; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_385 = 9'h181 == pht_ridx ? pht_385 : _GEN_384; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_386 = 9'h182 == pht_ridx ? pht_386 : _GEN_385; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_387 = 9'h183 == pht_ridx ? pht_387 : _GEN_386; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_388 = 9'h184 == pht_ridx ? pht_388 : _GEN_387; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_389 = 9'h185 == pht_ridx ? pht_389 : _GEN_388; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_390 = 9'h186 == pht_ridx ? pht_390 : _GEN_389; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_391 = 9'h187 == pht_ridx ? pht_391 : _GEN_390; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_392 = 9'h188 == pht_ridx ? pht_392 : _GEN_391; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_393 = 9'h189 == pht_ridx ? pht_393 : _GEN_392; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_394 = 9'h18a == pht_ridx ? pht_394 : _GEN_393; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_395 = 9'h18b == pht_ridx ? pht_395 : _GEN_394; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_396 = 9'h18c == pht_ridx ? pht_396 : _GEN_395; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_397 = 9'h18d == pht_ridx ? pht_397 : _GEN_396; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_398 = 9'h18e == pht_ridx ? pht_398 : _GEN_397; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_399 = 9'h18f == pht_ridx ? pht_399 : _GEN_398; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_400 = 9'h190 == pht_ridx ? pht_400 : _GEN_399; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_401 = 9'h191 == pht_ridx ? pht_401 : _GEN_400; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_402 = 9'h192 == pht_ridx ? pht_402 : _GEN_401; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_403 = 9'h193 == pht_ridx ? pht_403 : _GEN_402; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_404 = 9'h194 == pht_ridx ? pht_404 : _GEN_403; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_405 = 9'h195 == pht_ridx ? pht_405 : _GEN_404; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_406 = 9'h196 == pht_ridx ? pht_406 : _GEN_405; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_407 = 9'h197 == pht_ridx ? pht_407 : _GEN_406; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_408 = 9'h198 == pht_ridx ? pht_408 : _GEN_407; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_409 = 9'h199 == pht_ridx ? pht_409 : _GEN_408; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_410 = 9'h19a == pht_ridx ? pht_410 : _GEN_409; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_411 = 9'h19b == pht_ridx ? pht_411 : _GEN_410; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_412 = 9'h19c == pht_ridx ? pht_412 : _GEN_411; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_413 = 9'h19d == pht_ridx ? pht_413 : _GEN_412; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_414 = 9'h19e == pht_ridx ? pht_414 : _GEN_413; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_415 = 9'h19f == pht_ridx ? pht_415 : _GEN_414; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_416 = 9'h1a0 == pht_ridx ? pht_416 : _GEN_415; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_417 = 9'h1a1 == pht_ridx ? pht_417 : _GEN_416; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_418 = 9'h1a2 == pht_ridx ? pht_418 : _GEN_417; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_419 = 9'h1a3 == pht_ridx ? pht_419 : _GEN_418; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_420 = 9'h1a4 == pht_ridx ? pht_420 : _GEN_419; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_421 = 9'h1a5 == pht_ridx ? pht_421 : _GEN_420; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_422 = 9'h1a6 == pht_ridx ? pht_422 : _GEN_421; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_423 = 9'h1a7 == pht_ridx ? pht_423 : _GEN_422; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_424 = 9'h1a8 == pht_ridx ? pht_424 : _GEN_423; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_425 = 9'h1a9 == pht_ridx ? pht_425 : _GEN_424; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_426 = 9'h1aa == pht_ridx ? pht_426 : _GEN_425; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_427 = 9'h1ab == pht_ridx ? pht_427 : _GEN_426; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_428 = 9'h1ac == pht_ridx ? pht_428 : _GEN_427; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_429 = 9'h1ad == pht_ridx ? pht_429 : _GEN_428; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_430 = 9'h1ae == pht_ridx ? pht_430 : _GEN_429; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_431 = 9'h1af == pht_ridx ? pht_431 : _GEN_430; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_432 = 9'h1b0 == pht_ridx ? pht_432 : _GEN_431; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_433 = 9'h1b1 == pht_ridx ? pht_433 : _GEN_432; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_434 = 9'h1b2 == pht_ridx ? pht_434 : _GEN_433; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_435 = 9'h1b3 == pht_ridx ? pht_435 : _GEN_434; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_436 = 9'h1b4 == pht_ridx ? pht_436 : _GEN_435; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_437 = 9'h1b5 == pht_ridx ? pht_437 : _GEN_436; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_438 = 9'h1b6 == pht_ridx ? pht_438 : _GEN_437; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_439 = 9'h1b7 == pht_ridx ? pht_439 : _GEN_438; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_440 = 9'h1b8 == pht_ridx ? pht_440 : _GEN_439; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_441 = 9'h1b9 == pht_ridx ? pht_441 : _GEN_440; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_442 = 9'h1ba == pht_ridx ? pht_442 : _GEN_441; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_443 = 9'h1bb == pht_ridx ? pht_443 : _GEN_442; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_444 = 9'h1bc == pht_ridx ? pht_444 : _GEN_443; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_445 = 9'h1bd == pht_ridx ? pht_445 : _GEN_444; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_446 = 9'h1be == pht_ridx ? pht_446 : _GEN_445; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_447 = 9'h1bf == pht_ridx ? pht_447 : _GEN_446; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_448 = 9'h1c0 == pht_ridx ? pht_448 : _GEN_447; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_449 = 9'h1c1 == pht_ridx ? pht_449 : _GEN_448; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_450 = 9'h1c2 == pht_ridx ? pht_450 : _GEN_449; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_451 = 9'h1c3 == pht_ridx ? pht_451 : _GEN_450; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_452 = 9'h1c4 == pht_ridx ? pht_452 : _GEN_451; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_453 = 9'h1c5 == pht_ridx ? pht_453 : _GEN_452; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_454 = 9'h1c6 == pht_ridx ? pht_454 : _GEN_453; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_455 = 9'h1c7 == pht_ridx ? pht_455 : _GEN_454; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_456 = 9'h1c8 == pht_ridx ? pht_456 : _GEN_455; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_457 = 9'h1c9 == pht_ridx ? pht_457 : _GEN_456; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_458 = 9'h1ca == pht_ridx ? pht_458 : _GEN_457; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_459 = 9'h1cb == pht_ridx ? pht_459 : _GEN_458; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_460 = 9'h1cc == pht_ridx ? pht_460 : _GEN_459; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_461 = 9'h1cd == pht_ridx ? pht_461 : _GEN_460; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_462 = 9'h1ce == pht_ridx ? pht_462 : _GEN_461; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_463 = 9'h1cf == pht_ridx ? pht_463 : _GEN_462; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_464 = 9'h1d0 == pht_ridx ? pht_464 : _GEN_463; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_465 = 9'h1d1 == pht_ridx ? pht_465 : _GEN_464; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_466 = 9'h1d2 == pht_ridx ? pht_466 : _GEN_465; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_467 = 9'h1d3 == pht_ridx ? pht_467 : _GEN_466; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_468 = 9'h1d4 == pht_ridx ? pht_468 : _GEN_467; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_469 = 9'h1d5 == pht_ridx ? pht_469 : _GEN_468; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_470 = 9'h1d6 == pht_ridx ? pht_470 : _GEN_469; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_471 = 9'h1d7 == pht_ridx ? pht_471 : _GEN_470; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_472 = 9'h1d8 == pht_ridx ? pht_472 : _GEN_471; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_473 = 9'h1d9 == pht_ridx ? pht_473 : _GEN_472; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_474 = 9'h1da == pht_ridx ? pht_474 : _GEN_473; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_475 = 9'h1db == pht_ridx ? pht_475 : _GEN_474; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_476 = 9'h1dc == pht_ridx ? pht_476 : _GEN_475; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_477 = 9'h1dd == pht_ridx ? pht_477 : _GEN_476; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_478 = 9'h1de == pht_ridx ? pht_478 : _GEN_477; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_479 = 9'h1df == pht_ridx ? pht_479 : _GEN_478; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_480 = 9'h1e0 == pht_ridx ? pht_480 : _GEN_479; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_481 = 9'h1e1 == pht_ridx ? pht_481 : _GEN_480; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_482 = 9'h1e2 == pht_ridx ? pht_482 : _GEN_481; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_483 = 9'h1e3 == pht_ridx ? pht_483 : _GEN_482; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_484 = 9'h1e4 == pht_ridx ? pht_484 : _GEN_483; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_485 = 9'h1e5 == pht_ridx ? pht_485 : _GEN_484; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_486 = 9'h1e6 == pht_ridx ? pht_486 : _GEN_485; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_487 = 9'h1e7 == pht_ridx ? pht_487 : _GEN_486; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_488 = 9'h1e8 == pht_ridx ? pht_488 : _GEN_487; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_489 = 9'h1e9 == pht_ridx ? pht_489 : _GEN_488; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_490 = 9'h1ea == pht_ridx ? pht_490 : _GEN_489; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_491 = 9'h1eb == pht_ridx ? pht_491 : _GEN_490; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_492 = 9'h1ec == pht_ridx ? pht_492 : _GEN_491; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_493 = 9'h1ed == pht_ridx ? pht_493 : _GEN_492; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_494 = 9'h1ee == pht_ridx ? pht_494 : _GEN_493; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_495 = 9'h1ef == pht_ridx ? pht_495 : _GEN_494; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_496 = 9'h1f0 == pht_ridx ? pht_496 : _GEN_495; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_497 = 9'h1f1 == pht_ridx ? pht_497 : _GEN_496; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_498 = 9'h1f2 == pht_ridx ? pht_498 : _GEN_497; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_499 = 9'h1f3 == pht_ridx ? pht_499 : _GEN_498; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_500 = 9'h1f4 == pht_ridx ? pht_500 : _GEN_499; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_501 = 9'h1f5 == pht_ridx ? pht_501 : _GEN_500; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_502 = 9'h1f6 == pht_ridx ? pht_502 : _GEN_501; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_503 = 9'h1f7 == pht_ridx ? pht_503 : _GEN_502; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_504 = 9'h1f8 == pht_ridx ? pht_504 : _GEN_503; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_505 = 9'h1f9 == pht_ridx ? pht_505 : _GEN_504; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_506 = 9'h1fa == pht_ridx ? pht_506 : _GEN_505; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_507 = 9'h1fb == pht_ridx ? pht_507 : _GEN_506; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_508 = 9'h1fc == pht_ridx ? pht_508 : _GEN_507; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_509 = 9'h1fd == pht_ridx ? pht_509 : _GEN_508; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_510 = 9'h1fe == pht_ridx ? pht_510 : _GEN_509; // @[BPU.scala 33:{30,30}]
  wire [1:0] _GEN_511 = 9'h1ff == pht_ridx ? pht_511 : _GEN_510; // @[BPU.scala 33:{30,30}]
  wire  pht_taken = _GEN_511 >= 2'h2; // @[BPU.scala 33:30]
  wire [36:0] _GEN_513 = btb_0_valid & btb_0_tag == io_pc[38:2] ? btb_0_target : 37'h0; // @[BPU.scala 39:67 41:17 37:30]
  wire [36:0] _GEN_515 = btb_1_valid & btb_1_tag == io_pc[38:2] ? btb_1_target : _GEN_513; // @[BPU.scala 39:67 41:17]
  wire [36:0] _GEN_517 = btb_2_valid & btb_2_tag == io_pc[38:2] ? btb_2_target : _GEN_515; // @[BPU.scala 39:67 41:17]
  wire [36:0] _GEN_519 = btb_3_valid & btb_3_tag == io_pc[38:2] ? btb_3_target : _GEN_517; // @[BPU.scala 39:67 41:17]
  wire [36:0] _GEN_521 = btb_4_valid & btb_4_tag == io_pc[38:2] ? btb_4_target : _GEN_519; // @[BPU.scala 39:67 41:17]
  wire [36:0] _GEN_523 = btb_5_valid & btb_5_tag == io_pc[38:2] ? btb_5_target : _GEN_521; // @[BPU.scala 39:67 41:17]
  wire [36:0] _GEN_525 = btb_6_valid & btb_6_tag == io_pc[38:2] ? btb_6_target : _GEN_523; // @[BPU.scala 39:67 41:17]
  wire [36:0] _GEN_527 = btb_7_valid & btb_7_tag == io_pc[38:2] ? btb_7_target : _GEN_525; // @[BPU.scala 39:67 41:17]
  wire [36:0] _GEN_529 = btb_8_valid & btb_8_tag == io_pc[38:2] ? btb_8_target : _GEN_527; // @[BPU.scala 39:67 41:17]
  wire  _GEN_530 = btb_9_valid & btb_9_tag == io_pc[38:2] | (btb_8_valid & btb_8_tag == io_pc[38:2] | (btb_7_valid &
    btb_7_tag == io_pc[38:2] | (btb_6_valid & btb_6_tag == io_pc[38:2] | (btb_5_valid & btb_5_tag == io_pc[38:2] | (
    btb_4_valid & btb_4_tag == io_pc[38:2] | (btb_3_valid & btb_3_tag == io_pc[38:2] | (btb_2_valid & btb_2_tag == io_pc
    [38:2] | (btb_1_valid & btb_1_tag == io_pc[38:2] | btb_0_valid & btb_0_tag == io_pc[38:2])))))))); // @[BPU.scala 39:67 40:17]
  wire [36:0] _GEN_531 = btb_9_valid & btb_9_tag == io_pc[38:2] ? btb_9_target : _GEN_529; // @[BPU.scala 39:67 41:17]
  wire [36:0] _GEN_533 = btb_10_valid & btb_10_tag == io_pc[38:2] ? btb_10_target : _GEN_531; // @[BPU.scala 39:67 41:17]
  wire [36:0] _GEN_535 = btb_11_valid & btb_11_tag == io_pc[38:2] ? btb_11_target : _GEN_533; // @[BPU.scala 39:67 41:17]
  wire [36:0] _GEN_537 = btb_12_valid & btb_12_tag == io_pc[38:2] ? btb_12_target : _GEN_535; // @[BPU.scala 39:67 41:17]
  wire [36:0] _GEN_539 = btb_13_valid & btb_13_tag == io_pc[38:2] ? btb_13_target : _GEN_537; // @[BPU.scala 39:67 41:17]
  wire [36:0] _GEN_541 = btb_14_valid & btb_14_tag == io_pc[38:2] ? btb_14_target : _GEN_539; // @[BPU.scala 39:67 41:17]
  wire  btb_rhit = btb_15_valid & btb_15_tag == io_pc[38:2] | (btb_14_valid & btb_14_tag == io_pc[38:2] | (btb_13_valid
     & btb_13_tag == io_pc[38:2] | (btb_12_valid & btb_12_tag == io_pc[38:2] | (btb_11_valid & btb_11_tag == io_pc[38:2]
     | (btb_10_valid & btb_10_tag == io_pc[38:2] | _GEN_530))))); // @[BPU.scala 39:67 40:17]
  wire [36:0] btb_rdata = btb_15_valid & btb_15_tag == io_pc[38:2] ? btb_15_target : _GEN_541; // @[BPU.scala 39:67 41:17]
  wire [63:0] _io_out_T_1 = io_pc + 64'h4; // @[BPU.scala 46:19]
  wire [38:0] _io_out_T_2 = {btb_rdata,2'h0}; // @[Cat.scala 33:92]
  wire [24:0] _io_out_T_5 = _io_out_T_2[38] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _io_out_T_6 = {_io_out_T_5,btb_rdata,2'h0}; // @[Cat.scala 33:92]
  wire [8:0] pht_widx = io_jmp_packet_bp_pc[10:2] ^ ghr; // @[BPU.scala 52:53]
  wire [7:0] _ghr_T_1 = {ghr[7:1],io_jmp_packet_bp_taken}; // @[Cat.scala 33:92]
  wire [1:0] _pht_T_1 = io_jmp_packet_bp_taken ? 2'h2 : 2'h0; // @[BPU.scala 60:19]
  wire [1:0] _pht_T_2 = io_jmp_packet_bp_taken ? 2'h3 : 2'h1; // @[BPU.scala 61:19]
  wire [1:0] _pht_T_3 = io_jmp_packet_bp_taken ? 2'h3 : 2'h2; // @[BPU.scala 62:19]
  wire [1:0] _GEN_546 = 9'h1 == pht_widx ? pht_1 : pht_0; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_547 = 9'h2 == pht_widx ? pht_2 : _GEN_546; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_548 = 9'h3 == pht_widx ? pht_3 : _GEN_547; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_549 = 9'h4 == pht_widx ? pht_4 : _GEN_548; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_550 = 9'h5 == pht_widx ? pht_5 : _GEN_549; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_551 = 9'h6 == pht_widx ? pht_6 : _GEN_550; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_552 = 9'h7 == pht_widx ? pht_7 : _GEN_551; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_553 = 9'h8 == pht_widx ? pht_8 : _GEN_552; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_554 = 9'h9 == pht_widx ? pht_9 : _GEN_553; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_555 = 9'ha == pht_widx ? pht_10 : _GEN_554; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_556 = 9'hb == pht_widx ? pht_11 : _GEN_555; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_557 = 9'hc == pht_widx ? pht_12 : _GEN_556; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_558 = 9'hd == pht_widx ? pht_13 : _GEN_557; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_559 = 9'he == pht_widx ? pht_14 : _GEN_558; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_560 = 9'hf == pht_widx ? pht_15 : _GEN_559; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_561 = 9'h10 == pht_widx ? pht_16 : _GEN_560; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_562 = 9'h11 == pht_widx ? pht_17 : _GEN_561; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_563 = 9'h12 == pht_widx ? pht_18 : _GEN_562; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_564 = 9'h13 == pht_widx ? pht_19 : _GEN_563; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_565 = 9'h14 == pht_widx ? pht_20 : _GEN_564; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_566 = 9'h15 == pht_widx ? pht_21 : _GEN_565; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_567 = 9'h16 == pht_widx ? pht_22 : _GEN_566; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_568 = 9'h17 == pht_widx ? pht_23 : _GEN_567; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_569 = 9'h18 == pht_widx ? pht_24 : _GEN_568; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_570 = 9'h19 == pht_widx ? pht_25 : _GEN_569; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_571 = 9'h1a == pht_widx ? pht_26 : _GEN_570; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_572 = 9'h1b == pht_widx ? pht_27 : _GEN_571; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_573 = 9'h1c == pht_widx ? pht_28 : _GEN_572; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_574 = 9'h1d == pht_widx ? pht_29 : _GEN_573; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_575 = 9'h1e == pht_widx ? pht_30 : _GEN_574; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_576 = 9'h1f == pht_widx ? pht_31 : _GEN_575; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_577 = 9'h20 == pht_widx ? pht_32 : _GEN_576; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_578 = 9'h21 == pht_widx ? pht_33 : _GEN_577; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_579 = 9'h22 == pht_widx ? pht_34 : _GEN_578; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_580 = 9'h23 == pht_widx ? pht_35 : _GEN_579; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_581 = 9'h24 == pht_widx ? pht_36 : _GEN_580; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_582 = 9'h25 == pht_widx ? pht_37 : _GEN_581; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_583 = 9'h26 == pht_widx ? pht_38 : _GEN_582; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_584 = 9'h27 == pht_widx ? pht_39 : _GEN_583; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_585 = 9'h28 == pht_widx ? pht_40 : _GEN_584; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_586 = 9'h29 == pht_widx ? pht_41 : _GEN_585; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_587 = 9'h2a == pht_widx ? pht_42 : _GEN_586; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_588 = 9'h2b == pht_widx ? pht_43 : _GEN_587; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_589 = 9'h2c == pht_widx ? pht_44 : _GEN_588; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_590 = 9'h2d == pht_widx ? pht_45 : _GEN_589; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_591 = 9'h2e == pht_widx ? pht_46 : _GEN_590; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_592 = 9'h2f == pht_widx ? pht_47 : _GEN_591; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_593 = 9'h30 == pht_widx ? pht_48 : _GEN_592; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_594 = 9'h31 == pht_widx ? pht_49 : _GEN_593; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_595 = 9'h32 == pht_widx ? pht_50 : _GEN_594; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_596 = 9'h33 == pht_widx ? pht_51 : _GEN_595; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_597 = 9'h34 == pht_widx ? pht_52 : _GEN_596; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_598 = 9'h35 == pht_widx ? pht_53 : _GEN_597; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_599 = 9'h36 == pht_widx ? pht_54 : _GEN_598; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_600 = 9'h37 == pht_widx ? pht_55 : _GEN_599; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_601 = 9'h38 == pht_widx ? pht_56 : _GEN_600; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_602 = 9'h39 == pht_widx ? pht_57 : _GEN_601; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_603 = 9'h3a == pht_widx ? pht_58 : _GEN_602; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_604 = 9'h3b == pht_widx ? pht_59 : _GEN_603; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_605 = 9'h3c == pht_widx ? pht_60 : _GEN_604; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_606 = 9'h3d == pht_widx ? pht_61 : _GEN_605; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_607 = 9'h3e == pht_widx ? pht_62 : _GEN_606; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_608 = 9'h3f == pht_widx ? pht_63 : _GEN_607; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_609 = 9'h40 == pht_widx ? pht_64 : _GEN_608; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_610 = 9'h41 == pht_widx ? pht_65 : _GEN_609; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_611 = 9'h42 == pht_widx ? pht_66 : _GEN_610; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_612 = 9'h43 == pht_widx ? pht_67 : _GEN_611; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_613 = 9'h44 == pht_widx ? pht_68 : _GEN_612; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_614 = 9'h45 == pht_widx ? pht_69 : _GEN_613; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_615 = 9'h46 == pht_widx ? pht_70 : _GEN_614; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_616 = 9'h47 == pht_widx ? pht_71 : _GEN_615; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_617 = 9'h48 == pht_widx ? pht_72 : _GEN_616; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_618 = 9'h49 == pht_widx ? pht_73 : _GEN_617; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_619 = 9'h4a == pht_widx ? pht_74 : _GEN_618; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_620 = 9'h4b == pht_widx ? pht_75 : _GEN_619; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_621 = 9'h4c == pht_widx ? pht_76 : _GEN_620; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_622 = 9'h4d == pht_widx ? pht_77 : _GEN_621; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_623 = 9'h4e == pht_widx ? pht_78 : _GEN_622; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_624 = 9'h4f == pht_widx ? pht_79 : _GEN_623; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_625 = 9'h50 == pht_widx ? pht_80 : _GEN_624; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_626 = 9'h51 == pht_widx ? pht_81 : _GEN_625; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_627 = 9'h52 == pht_widx ? pht_82 : _GEN_626; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_628 = 9'h53 == pht_widx ? pht_83 : _GEN_627; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_629 = 9'h54 == pht_widx ? pht_84 : _GEN_628; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_630 = 9'h55 == pht_widx ? pht_85 : _GEN_629; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_631 = 9'h56 == pht_widx ? pht_86 : _GEN_630; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_632 = 9'h57 == pht_widx ? pht_87 : _GEN_631; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_633 = 9'h58 == pht_widx ? pht_88 : _GEN_632; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_634 = 9'h59 == pht_widx ? pht_89 : _GEN_633; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_635 = 9'h5a == pht_widx ? pht_90 : _GEN_634; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_636 = 9'h5b == pht_widx ? pht_91 : _GEN_635; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_637 = 9'h5c == pht_widx ? pht_92 : _GEN_636; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_638 = 9'h5d == pht_widx ? pht_93 : _GEN_637; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_639 = 9'h5e == pht_widx ? pht_94 : _GEN_638; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_640 = 9'h5f == pht_widx ? pht_95 : _GEN_639; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_641 = 9'h60 == pht_widx ? pht_96 : _GEN_640; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_642 = 9'h61 == pht_widx ? pht_97 : _GEN_641; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_643 = 9'h62 == pht_widx ? pht_98 : _GEN_642; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_644 = 9'h63 == pht_widx ? pht_99 : _GEN_643; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_645 = 9'h64 == pht_widx ? pht_100 : _GEN_644; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_646 = 9'h65 == pht_widx ? pht_101 : _GEN_645; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_647 = 9'h66 == pht_widx ? pht_102 : _GEN_646; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_648 = 9'h67 == pht_widx ? pht_103 : _GEN_647; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_649 = 9'h68 == pht_widx ? pht_104 : _GEN_648; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_650 = 9'h69 == pht_widx ? pht_105 : _GEN_649; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_651 = 9'h6a == pht_widx ? pht_106 : _GEN_650; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_652 = 9'h6b == pht_widx ? pht_107 : _GEN_651; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_653 = 9'h6c == pht_widx ? pht_108 : _GEN_652; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_654 = 9'h6d == pht_widx ? pht_109 : _GEN_653; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_655 = 9'h6e == pht_widx ? pht_110 : _GEN_654; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_656 = 9'h6f == pht_widx ? pht_111 : _GEN_655; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_657 = 9'h70 == pht_widx ? pht_112 : _GEN_656; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_658 = 9'h71 == pht_widx ? pht_113 : _GEN_657; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_659 = 9'h72 == pht_widx ? pht_114 : _GEN_658; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_660 = 9'h73 == pht_widx ? pht_115 : _GEN_659; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_661 = 9'h74 == pht_widx ? pht_116 : _GEN_660; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_662 = 9'h75 == pht_widx ? pht_117 : _GEN_661; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_663 = 9'h76 == pht_widx ? pht_118 : _GEN_662; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_664 = 9'h77 == pht_widx ? pht_119 : _GEN_663; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_665 = 9'h78 == pht_widx ? pht_120 : _GEN_664; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_666 = 9'h79 == pht_widx ? pht_121 : _GEN_665; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_667 = 9'h7a == pht_widx ? pht_122 : _GEN_666; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_668 = 9'h7b == pht_widx ? pht_123 : _GEN_667; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_669 = 9'h7c == pht_widx ? pht_124 : _GEN_668; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_670 = 9'h7d == pht_widx ? pht_125 : _GEN_669; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_671 = 9'h7e == pht_widx ? pht_126 : _GEN_670; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_672 = 9'h7f == pht_widx ? pht_127 : _GEN_671; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_673 = 9'h80 == pht_widx ? pht_128 : _GEN_672; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_674 = 9'h81 == pht_widx ? pht_129 : _GEN_673; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_675 = 9'h82 == pht_widx ? pht_130 : _GEN_674; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_676 = 9'h83 == pht_widx ? pht_131 : _GEN_675; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_677 = 9'h84 == pht_widx ? pht_132 : _GEN_676; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_678 = 9'h85 == pht_widx ? pht_133 : _GEN_677; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_679 = 9'h86 == pht_widx ? pht_134 : _GEN_678; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_680 = 9'h87 == pht_widx ? pht_135 : _GEN_679; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_681 = 9'h88 == pht_widx ? pht_136 : _GEN_680; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_682 = 9'h89 == pht_widx ? pht_137 : _GEN_681; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_683 = 9'h8a == pht_widx ? pht_138 : _GEN_682; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_684 = 9'h8b == pht_widx ? pht_139 : _GEN_683; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_685 = 9'h8c == pht_widx ? pht_140 : _GEN_684; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_686 = 9'h8d == pht_widx ? pht_141 : _GEN_685; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_687 = 9'h8e == pht_widx ? pht_142 : _GEN_686; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_688 = 9'h8f == pht_widx ? pht_143 : _GEN_687; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_689 = 9'h90 == pht_widx ? pht_144 : _GEN_688; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_690 = 9'h91 == pht_widx ? pht_145 : _GEN_689; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_691 = 9'h92 == pht_widx ? pht_146 : _GEN_690; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_692 = 9'h93 == pht_widx ? pht_147 : _GEN_691; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_693 = 9'h94 == pht_widx ? pht_148 : _GEN_692; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_694 = 9'h95 == pht_widx ? pht_149 : _GEN_693; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_695 = 9'h96 == pht_widx ? pht_150 : _GEN_694; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_696 = 9'h97 == pht_widx ? pht_151 : _GEN_695; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_697 = 9'h98 == pht_widx ? pht_152 : _GEN_696; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_698 = 9'h99 == pht_widx ? pht_153 : _GEN_697; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_699 = 9'h9a == pht_widx ? pht_154 : _GEN_698; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_700 = 9'h9b == pht_widx ? pht_155 : _GEN_699; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_701 = 9'h9c == pht_widx ? pht_156 : _GEN_700; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_702 = 9'h9d == pht_widx ? pht_157 : _GEN_701; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_703 = 9'h9e == pht_widx ? pht_158 : _GEN_702; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_704 = 9'h9f == pht_widx ? pht_159 : _GEN_703; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_705 = 9'ha0 == pht_widx ? pht_160 : _GEN_704; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_706 = 9'ha1 == pht_widx ? pht_161 : _GEN_705; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_707 = 9'ha2 == pht_widx ? pht_162 : _GEN_706; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_708 = 9'ha3 == pht_widx ? pht_163 : _GEN_707; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_709 = 9'ha4 == pht_widx ? pht_164 : _GEN_708; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_710 = 9'ha5 == pht_widx ? pht_165 : _GEN_709; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_711 = 9'ha6 == pht_widx ? pht_166 : _GEN_710; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_712 = 9'ha7 == pht_widx ? pht_167 : _GEN_711; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_713 = 9'ha8 == pht_widx ? pht_168 : _GEN_712; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_714 = 9'ha9 == pht_widx ? pht_169 : _GEN_713; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_715 = 9'haa == pht_widx ? pht_170 : _GEN_714; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_716 = 9'hab == pht_widx ? pht_171 : _GEN_715; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_717 = 9'hac == pht_widx ? pht_172 : _GEN_716; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_718 = 9'had == pht_widx ? pht_173 : _GEN_717; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_719 = 9'hae == pht_widx ? pht_174 : _GEN_718; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_720 = 9'haf == pht_widx ? pht_175 : _GEN_719; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_721 = 9'hb0 == pht_widx ? pht_176 : _GEN_720; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_722 = 9'hb1 == pht_widx ? pht_177 : _GEN_721; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_723 = 9'hb2 == pht_widx ? pht_178 : _GEN_722; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_724 = 9'hb3 == pht_widx ? pht_179 : _GEN_723; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_725 = 9'hb4 == pht_widx ? pht_180 : _GEN_724; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_726 = 9'hb5 == pht_widx ? pht_181 : _GEN_725; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_727 = 9'hb6 == pht_widx ? pht_182 : _GEN_726; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_728 = 9'hb7 == pht_widx ? pht_183 : _GEN_727; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_729 = 9'hb8 == pht_widx ? pht_184 : _GEN_728; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_730 = 9'hb9 == pht_widx ? pht_185 : _GEN_729; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_731 = 9'hba == pht_widx ? pht_186 : _GEN_730; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_732 = 9'hbb == pht_widx ? pht_187 : _GEN_731; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_733 = 9'hbc == pht_widx ? pht_188 : _GEN_732; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_734 = 9'hbd == pht_widx ? pht_189 : _GEN_733; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_735 = 9'hbe == pht_widx ? pht_190 : _GEN_734; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_736 = 9'hbf == pht_widx ? pht_191 : _GEN_735; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_737 = 9'hc0 == pht_widx ? pht_192 : _GEN_736; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_738 = 9'hc1 == pht_widx ? pht_193 : _GEN_737; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_739 = 9'hc2 == pht_widx ? pht_194 : _GEN_738; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_740 = 9'hc3 == pht_widx ? pht_195 : _GEN_739; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_741 = 9'hc4 == pht_widx ? pht_196 : _GEN_740; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_742 = 9'hc5 == pht_widx ? pht_197 : _GEN_741; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_743 = 9'hc6 == pht_widx ? pht_198 : _GEN_742; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_744 = 9'hc7 == pht_widx ? pht_199 : _GEN_743; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_745 = 9'hc8 == pht_widx ? pht_200 : _GEN_744; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_746 = 9'hc9 == pht_widx ? pht_201 : _GEN_745; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_747 = 9'hca == pht_widx ? pht_202 : _GEN_746; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_748 = 9'hcb == pht_widx ? pht_203 : _GEN_747; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_749 = 9'hcc == pht_widx ? pht_204 : _GEN_748; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_750 = 9'hcd == pht_widx ? pht_205 : _GEN_749; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_751 = 9'hce == pht_widx ? pht_206 : _GEN_750; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_752 = 9'hcf == pht_widx ? pht_207 : _GEN_751; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_753 = 9'hd0 == pht_widx ? pht_208 : _GEN_752; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_754 = 9'hd1 == pht_widx ? pht_209 : _GEN_753; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_755 = 9'hd2 == pht_widx ? pht_210 : _GEN_754; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_756 = 9'hd3 == pht_widx ? pht_211 : _GEN_755; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_757 = 9'hd4 == pht_widx ? pht_212 : _GEN_756; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_758 = 9'hd5 == pht_widx ? pht_213 : _GEN_757; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_759 = 9'hd6 == pht_widx ? pht_214 : _GEN_758; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_760 = 9'hd7 == pht_widx ? pht_215 : _GEN_759; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_761 = 9'hd8 == pht_widx ? pht_216 : _GEN_760; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_762 = 9'hd9 == pht_widx ? pht_217 : _GEN_761; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_763 = 9'hda == pht_widx ? pht_218 : _GEN_762; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_764 = 9'hdb == pht_widx ? pht_219 : _GEN_763; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_765 = 9'hdc == pht_widx ? pht_220 : _GEN_764; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_766 = 9'hdd == pht_widx ? pht_221 : _GEN_765; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_767 = 9'hde == pht_widx ? pht_222 : _GEN_766; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_768 = 9'hdf == pht_widx ? pht_223 : _GEN_767; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_769 = 9'he0 == pht_widx ? pht_224 : _GEN_768; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_770 = 9'he1 == pht_widx ? pht_225 : _GEN_769; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_771 = 9'he2 == pht_widx ? pht_226 : _GEN_770; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_772 = 9'he3 == pht_widx ? pht_227 : _GEN_771; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_773 = 9'he4 == pht_widx ? pht_228 : _GEN_772; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_774 = 9'he5 == pht_widx ? pht_229 : _GEN_773; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_775 = 9'he6 == pht_widx ? pht_230 : _GEN_774; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_776 = 9'he7 == pht_widx ? pht_231 : _GEN_775; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_777 = 9'he8 == pht_widx ? pht_232 : _GEN_776; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_778 = 9'he9 == pht_widx ? pht_233 : _GEN_777; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_779 = 9'hea == pht_widx ? pht_234 : _GEN_778; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_780 = 9'heb == pht_widx ? pht_235 : _GEN_779; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_781 = 9'hec == pht_widx ? pht_236 : _GEN_780; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_782 = 9'hed == pht_widx ? pht_237 : _GEN_781; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_783 = 9'hee == pht_widx ? pht_238 : _GEN_782; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_784 = 9'hef == pht_widx ? pht_239 : _GEN_783; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_785 = 9'hf0 == pht_widx ? pht_240 : _GEN_784; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_786 = 9'hf1 == pht_widx ? pht_241 : _GEN_785; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_787 = 9'hf2 == pht_widx ? pht_242 : _GEN_786; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_788 = 9'hf3 == pht_widx ? pht_243 : _GEN_787; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_789 = 9'hf4 == pht_widx ? pht_244 : _GEN_788; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_790 = 9'hf5 == pht_widx ? pht_245 : _GEN_789; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_791 = 9'hf6 == pht_widx ? pht_246 : _GEN_790; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_792 = 9'hf7 == pht_widx ? pht_247 : _GEN_791; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_793 = 9'hf8 == pht_widx ? pht_248 : _GEN_792; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_794 = 9'hf9 == pht_widx ? pht_249 : _GEN_793; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_795 = 9'hfa == pht_widx ? pht_250 : _GEN_794; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_796 = 9'hfb == pht_widx ? pht_251 : _GEN_795; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_797 = 9'hfc == pht_widx ? pht_252 : _GEN_796; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_798 = 9'hfd == pht_widx ? pht_253 : _GEN_797; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_799 = 9'hfe == pht_widx ? pht_254 : _GEN_798; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_800 = 9'hff == pht_widx ? pht_255 : _GEN_799; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_801 = 9'h100 == pht_widx ? pht_256 : _GEN_800; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_802 = 9'h101 == pht_widx ? pht_257 : _GEN_801; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_803 = 9'h102 == pht_widx ? pht_258 : _GEN_802; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_804 = 9'h103 == pht_widx ? pht_259 : _GEN_803; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_805 = 9'h104 == pht_widx ? pht_260 : _GEN_804; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_806 = 9'h105 == pht_widx ? pht_261 : _GEN_805; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_807 = 9'h106 == pht_widx ? pht_262 : _GEN_806; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_808 = 9'h107 == pht_widx ? pht_263 : _GEN_807; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_809 = 9'h108 == pht_widx ? pht_264 : _GEN_808; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_810 = 9'h109 == pht_widx ? pht_265 : _GEN_809; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_811 = 9'h10a == pht_widx ? pht_266 : _GEN_810; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_812 = 9'h10b == pht_widx ? pht_267 : _GEN_811; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_813 = 9'h10c == pht_widx ? pht_268 : _GEN_812; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_814 = 9'h10d == pht_widx ? pht_269 : _GEN_813; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_815 = 9'h10e == pht_widx ? pht_270 : _GEN_814; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_816 = 9'h10f == pht_widx ? pht_271 : _GEN_815; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_817 = 9'h110 == pht_widx ? pht_272 : _GEN_816; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_818 = 9'h111 == pht_widx ? pht_273 : _GEN_817; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_819 = 9'h112 == pht_widx ? pht_274 : _GEN_818; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_820 = 9'h113 == pht_widx ? pht_275 : _GEN_819; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_821 = 9'h114 == pht_widx ? pht_276 : _GEN_820; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_822 = 9'h115 == pht_widx ? pht_277 : _GEN_821; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_823 = 9'h116 == pht_widx ? pht_278 : _GEN_822; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_824 = 9'h117 == pht_widx ? pht_279 : _GEN_823; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_825 = 9'h118 == pht_widx ? pht_280 : _GEN_824; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_826 = 9'h119 == pht_widx ? pht_281 : _GEN_825; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_827 = 9'h11a == pht_widx ? pht_282 : _GEN_826; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_828 = 9'h11b == pht_widx ? pht_283 : _GEN_827; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_829 = 9'h11c == pht_widx ? pht_284 : _GEN_828; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_830 = 9'h11d == pht_widx ? pht_285 : _GEN_829; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_831 = 9'h11e == pht_widx ? pht_286 : _GEN_830; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_832 = 9'h11f == pht_widx ? pht_287 : _GEN_831; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_833 = 9'h120 == pht_widx ? pht_288 : _GEN_832; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_834 = 9'h121 == pht_widx ? pht_289 : _GEN_833; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_835 = 9'h122 == pht_widx ? pht_290 : _GEN_834; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_836 = 9'h123 == pht_widx ? pht_291 : _GEN_835; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_837 = 9'h124 == pht_widx ? pht_292 : _GEN_836; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_838 = 9'h125 == pht_widx ? pht_293 : _GEN_837; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_839 = 9'h126 == pht_widx ? pht_294 : _GEN_838; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_840 = 9'h127 == pht_widx ? pht_295 : _GEN_839; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_841 = 9'h128 == pht_widx ? pht_296 : _GEN_840; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_842 = 9'h129 == pht_widx ? pht_297 : _GEN_841; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_843 = 9'h12a == pht_widx ? pht_298 : _GEN_842; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_844 = 9'h12b == pht_widx ? pht_299 : _GEN_843; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_845 = 9'h12c == pht_widx ? pht_300 : _GEN_844; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_846 = 9'h12d == pht_widx ? pht_301 : _GEN_845; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_847 = 9'h12e == pht_widx ? pht_302 : _GEN_846; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_848 = 9'h12f == pht_widx ? pht_303 : _GEN_847; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_849 = 9'h130 == pht_widx ? pht_304 : _GEN_848; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_850 = 9'h131 == pht_widx ? pht_305 : _GEN_849; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_851 = 9'h132 == pht_widx ? pht_306 : _GEN_850; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_852 = 9'h133 == pht_widx ? pht_307 : _GEN_851; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_853 = 9'h134 == pht_widx ? pht_308 : _GEN_852; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_854 = 9'h135 == pht_widx ? pht_309 : _GEN_853; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_855 = 9'h136 == pht_widx ? pht_310 : _GEN_854; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_856 = 9'h137 == pht_widx ? pht_311 : _GEN_855; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_857 = 9'h138 == pht_widx ? pht_312 : _GEN_856; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_858 = 9'h139 == pht_widx ? pht_313 : _GEN_857; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_859 = 9'h13a == pht_widx ? pht_314 : _GEN_858; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_860 = 9'h13b == pht_widx ? pht_315 : _GEN_859; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_861 = 9'h13c == pht_widx ? pht_316 : _GEN_860; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_862 = 9'h13d == pht_widx ? pht_317 : _GEN_861; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_863 = 9'h13e == pht_widx ? pht_318 : _GEN_862; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_864 = 9'h13f == pht_widx ? pht_319 : _GEN_863; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_865 = 9'h140 == pht_widx ? pht_320 : _GEN_864; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_866 = 9'h141 == pht_widx ? pht_321 : _GEN_865; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_867 = 9'h142 == pht_widx ? pht_322 : _GEN_866; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_868 = 9'h143 == pht_widx ? pht_323 : _GEN_867; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_869 = 9'h144 == pht_widx ? pht_324 : _GEN_868; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_870 = 9'h145 == pht_widx ? pht_325 : _GEN_869; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_871 = 9'h146 == pht_widx ? pht_326 : _GEN_870; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_872 = 9'h147 == pht_widx ? pht_327 : _GEN_871; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_873 = 9'h148 == pht_widx ? pht_328 : _GEN_872; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_874 = 9'h149 == pht_widx ? pht_329 : _GEN_873; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_875 = 9'h14a == pht_widx ? pht_330 : _GEN_874; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_876 = 9'h14b == pht_widx ? pht_331 : _GEN_875; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_877 = 9'h14c == pht_widx ? pht_332 : _GEN_876; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_878 = 9'h14d == pht_widx ? pht_333 : _GEN_877; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_879 = 9'h14e == pht_widx ? pht_334 : _GEN_878; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_880 = 9'h14f == pht_widx ? pht_335 : _GEN_879; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_881 = 9'h150 == pht_widx ? pht_336 : _GEN_880; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_882 = 9'h151 == pht_widx ? pht_337 : _GEN_881; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_883 = 9'h152 == pht_widx ? pht_338 : _GEN_882; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_884 = 9'h153 == pht_widx ? pht_339 : _GEN_883; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_885 = 9'h154 == pht_widx ? pht_340 : _GEN_884; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_886 = 9'h155 == pht_widx ? pht_341 : _GEN_885; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_887 = 9'h156 == pht_widx ? pht_342 : _GEN_886; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_888 = 9'h157 == pht_widx ? pht_343 : _GEN_887; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_889 = 9'h158 == pht_widx ? pht_344 : _GEN_888; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_890 = 9'h159 == pht_widx ? pht_345 : _GEN_889; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_891 = 9'h15a == pht_widx ? pht_346 : _GEN_890; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_892 = 9'h15b == pht_widx ? pht_347 : _GEN_891; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_893 = 9'h15c == pht_widx ? pht_348 : _GEN_892; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_894 = 9'h15d == pht_widx ? pht_349 : _GEN_893; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_895 = 9'h15e == pht_widx ? pht_350 : _GEN_894; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_896 = 9'h15f == pht_widx ? pht_351 : _GEN_895; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_897 = 9'h160 == pht_widx ? pht_352 : _GEN_896; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_898 = 9'h161 == pht_widx ? pht_353 : _GEN_897; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_899 = 9'h162 == pht_widx ? pht_354 : _GEN_898; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_900 = 9'h163 == pht_widx ? pht_355 : _GEN_899; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_901 = 9'h164 == pht_widx ? pht_356 : _GEN_900; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_902 = 9'h165 == pht_widx ? pht_357 : _GEN_901; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_903 = 9'h166 == pht_widx ? pht_358 : _GEN_902; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_904 = 9'h167 == pht_widx ? pht_359 : _GEN_903; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_905 = 9'h168 == pht_widx ? pht_360 : _GEN_904; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_906 = 9'h169 == pht_widx ? pht_361 : _GEN_905; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_907 = 9'h16a == pht_widx ? pht_362 : _GEN_906; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_908 = 9'h16b == pht_widx ? pht_363 : _GEN_907; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_909 = 9'h16c == pht_widx ? pht_364 : _GEN_908; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_910 = 9'h16d == pht_widx ? pht_365 : _GEN_909; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_911 = 9'h16e == pht_widx ? pht_366 : _GEN_910; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_912 = 9'h16f == pht_widx ? pht_367 : _GEN_911; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_913 = 9'h170 == pht_widx ? pht_368 : _GEN_912; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_914 = 9'h171 == pht_widx ? pht_369 : _GEN_913; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_915 = 9'h172 == pht_widx ? pht_370 : _GEN_914; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_916 = 9'h173 == pht_widx ? pht_371 : _GEN_915; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_917 = 9'h174 == pht_widx ? pht_372 : _GEN_916; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_918 = 9'h175 == pht_widx ? pht_373 : _GEN_917; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_919 = 9'h176 == pht_widx ? pht_374 : _GEN_918; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_920 = 9'h177 == pht_widx ? pht_375 : _GEN_919; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_921 = 9'h178 == pht_widx ? pht_376 : _GEN_920; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_922 = 9'h179 == pht_widx ? pht_377 : _GEN_921; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_923 = 9'h17a == pht_widx ? pht_378 : _GEN_922; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_924 = 9'h17b == pht_widx ? pht_379 : _GEN_923; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_925 = 9'h17c == pht_widx ? pht_380 : _GEN_924; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_926 = 9'h17d == pht_widx ? pht_381 : _GEN_925; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_927 = 9'h17e == pht_widx ? pht_382 : _GEN_926; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_928 = 9'h17f == pht_widx ? pht_383 : _GEN_927; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_929 = 9'h180 == pht_widx ? pht_384 : _GEN_928; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_930 = 9'h181 == pht_widx ? pht_385 : _GEN_929; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_931 = 9'h182 == pht_widx ? pht_386 : _GEN_930; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_932 = 9'h183 == pht_widx ? pht_387 : _GEN_931; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_933 = 9'h184 == pht_widx ? pht_388 : _GEN_932; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_934 = 9'h185 == pht_widx ? pht_389 : _GEN_933; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_935 = 9'h186 == pht_widx ? pht_390 : _GEN_934; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_936 = 9'h187 == pht_widx ? pht_391 : _GEN_935; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_937 = 9'h188 == pht_widx ? pht_392 : _GEN_936; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_938 = 9'h189 == pht_widx ? pht_393 : _GEN_937; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_939 = 9'h18a == pht_widx ? pht_394 : _GEN_938; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_940 = 9'h18b == pht_widx ? pht_395 : _GEN_939; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_941 = 9'h18c == pht_widx ? pht_396 : _GEN_940; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_942 = 9'h18d == pht_widx ? pht_397 : _GEN_941; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_943 = 9'h18e == pht_widx ? pht_398 : _GEN_942; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_944 = 9'h18f == pht_widx ? pht_399 : _GEN_943; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_945 = 9'h190 == pht_widx ? pht_400 : _GEN_944; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_946 = 9'h191 == pht_widx ? pht_401 : _GEN_945; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_947 = 9'h192 == pht_widx ? pht_402 : _GEN_946; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_948 = 9'h193 == pht_widx ? pht_403 : _GEN_947; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_949 = 9'h194 == pht_widx ? pht_404 : _GEN_948; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_950 = 9'h195 == pht_widx ? pht_405 : _GEN_949; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_951 = 9'h196 == pht_widx ? pht_406 : _GEN_950; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_952 = 9'h197 == pht_widx ? pht_407 : _GEN_951; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_953 = 9'h198 == pht_widx ? pht_408 : _GEN_952; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_954 = 9'h199 == pht_widx ? pht_409 : _GEN_953; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_955 = 9'h19a == pht_widx ? pht_410 : _GEN_954; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_956 = 9'h19b == pht_widx ? pht_411 : _GEN_955; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_957 = 9'h19c == pht_widx ? pht_412 : _GEN_956; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_958 = 9'h19d == pht_widx ? pht_413 : _GEN_957; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_959 = 9'h19e == pht_widx ? pht_414 : _GEN_958; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_960 = 9'h19f == pht_widx ? pht_415 : _GEN_959; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_961 = 9'h1a0 == pht_widx ? pht_416 : _GEN_960; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_962 = 9'h1a1 == pht_widx ? pht_417 : _GEN_961; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_963 = 9'h1a2 == pht_widx ? pht_418 : _GEN_962; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_964 = 9'h1a3 == pht_widx ? pht_419 : _GEN_963; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_965 = 9'h1a4 == pht_widx ? pht_420 : _GEN_964; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_966 = 9'h1a5 == pht_widx ? pht_421 : _GEN_965; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_967 = 9'h1a6 == pht_widx ? pht_422 : _GEN_966; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_968 = 9'h1a7 == pht_widx ? pht_423 : _GEN_967; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_969 = 9'h1a8 == pht_widx ? pht_424 : _GEN_968; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_970 = 9'h1a9 == pht_widx ? pht_425 : _GEN_969; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_971 = 9'h1aa == pht_widx ? pht_426 : _GEN_970; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_972 = 9'h1ab == pht_widx ? pht_427 : _GEN_971; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_973 = 9'h1ac == pht_widx ? pht_428 : _GEN_972; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_974 = 9'h1ad == pht_widx ? pht_429 : _GEN_973; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_975 = 9'h1ae == pht_widx ? pht_430 : _GEN_974; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_976 = 9'h1af == pht_widx ? pht_431 : _GEN_975; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_977 = 9'h1b0 == pht_widx ? pht_432 : _GEN_976; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_978 = 9'h1b1 == pht_widx ? pht_433 : _GEN_977; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_979 = 9'h1b2 == pht_widx ? pht_434 : _GEN_978; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_980 = 9'h1b3 == pht_widx ? pht_435 : _GEN_979; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_981 = 9'h1b4 == pht_widx ? pht_436 : _GEN_980; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_982 = 9'h1b5 == pht_widx ? pht_437 : _GEN_981; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_983 = 9'h1b6 == pht_widx ? pht_438 : _GEN_982; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_984 = 9'h1b7 == pht_widx ? pht_439 : _GEN_983; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_985 = 9'h1b8 == pht_widx ? pht_440 : _GEN_984; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_986 = 9'h1b9 == pht_widx ? pht_441 : _GEN_985; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_987 = 9'h1ba == pht_widx ? pht_442 : _GEN_986; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_988 = 9'h1bb == pht_widx ? pht_443 : _GEN_987; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_989 = 9'h1bc == pht_widx ? pht_444 : _GEN_988; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_990 = 9'h1bd == pht_widx ? pht_445 : _GEN_989; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_991 = 9'h1be == pht_widx ? pht_446 : _GEN_990; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_992 = 9'h1bf == pht_widx ? pht_447 : _GEN_991; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_993 = 9'h1c0 == pht_widx ? pht_448 : _GEN_992; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_994 = 9'h1c1 == pht_widx ? pht_449 : _GEN_993; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_995 = 9'h1c2 == pht_widx ? pht_450 : _GEN_994; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_996 = 9'h1c3 == pht_widx ? pht_451 : _GEN_995; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_997 = 9'h1c4 == pht_widx ? pht_452 : _GEN_996; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_998 = 9'h1c5 == pht_widx ? pht_453 : _GEN_997; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_999 = 9'h1c6 == pht_widx ? pht_454 : _GEN_998; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1000 = 9'h1c7 == pht_widx ? pht_455 : _GEN_999; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1001 = 9'h1c8 == pht_widx ? pht_456 : _GEN_1000; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1002 = 9'h1c9 == pht_widx ? pht_457 : _GEN_1001; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1003 = 9'h1ca == pht_widx ? pht_458 : _GEN_1002; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1004 = 9'h1cb == pht_widx ? pht_459 : _GEN_1003; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1005 = 9'h1cc == pht_widx ? pht_460 : _GEN_1004; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1006 = 9'h1cd == pht_widx ? pht_461 : _GEN_1005; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1007 = 9'h1ce == pht_widx ? pht_462 : _GEN_1006; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1008 = 9'h1cf == pht_widx ? pht_463 : _GEN_1007; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1009 = 9'h1d0 == pht_widx ? pht_464 : _GEN_1008; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1010 = 9'h1d1 == pht_widx ? pht_465 : _GEN_1009; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1011 = 9'h1d2 == pht_widx ? pht_466 : _GEN_1010; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1012 = 9'h1d3 == pht_widx ? pht_467 : _GEN_1011; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1013 = 9'h1d4 == pht_widx ? pht_468 : _GEN_1012; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1014 = 9'h1d5 == pht_widx ? pht_469 : _GEN_1013; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1015 = 9'h1d6 == pht_widx ? pht_470 : _GEN_1014; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1016 = 9'h1d7 == pht_widx ? pht_471 : _GEN_1015; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1017 = 9'h1d8 == pht_widx ? pht_472 : _GEN_1016; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1018 = 9'h1d9 == pht_widx ? pht_473 : _GEN_1017; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1019 = 9'h1da == pht_widx ? pht_474 : _GEN_1018; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1020 = 9'h1db == pht_widx ? pht_475 : _GEN_1019; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1021 = 9'h1dc == pht_widx ? pht_476 : _GEN_1020; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1022 = 9'h1dd == pht_widx ? pht_477 : _GEN_1021; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1023 = 9'h1de == pht_widx ? pht_478 : _GEN_1022; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1024 = 9'h1df == pht_widx ? pht_479 : _GEN_1023; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1025 = 9'h1e0 == pht_widx ? pht_480 : _GEN_1024; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1026 = 9'h1e1 == pht_widx ? pht_481 : _GEN_1025; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1027 = 9'h1e2 == pht_widx ? pht_482 : _GEN_1026; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1028 = 9'h1e3 == pht_widx ? pht_483 : _GEN_1027; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1029 = 9'h1e4 == pht_widx ? pht_484 : _GEN_1028; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1030 = 9'h1e5 == pht_widx ? pht_485 : _GEN_1029; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1031 = 9'h1e6 == pht_widx ? pht_486 : _GEN_1030; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1032 = 9'h1e7 == pht_widx ? pht_487 : _GEN_1031; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1033 = 9'h1e8 == pht_widx ? pht_488 : _GEN_1032; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1034 = 9'h1e9 == pht_widx ? pht_489 : _GEN_1033; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1035 = 9'h1ea == pht_widx ? pht_490 : _GEN_1034; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1036 = 9'h1eb == pht_widx ? pht_491 : _GEN_1035; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1037 = 9'h1ec == pht_widx ? pht_492 : _GEN_1036; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1038 = 9'h1ed == pht_widx ? pht_493 : _GEN_1037; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1039 = 9'h1ee == pht_widx ? pht_494 : _GEN_1038; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1040 = 9'h1ef == pht_widx ? pht_495 : _GEN_1039; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1041 = 9'h1f0 == pht_widx ? pht_496 : _GEN_1040; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1042 = 9'h1f1 == pht_widx ? pht_497 : _GEN_1041; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1043 = 9'h1f2 == pht_widx ? pht_498 : _GEN_1042; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1044 = 9'h1f3 == pht_widx ? pht_499 : _GEN_1043; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1045 = 9'h1f4 == pht_widx ? pht_500 : _GEN_1044; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1046 = 9'h1f5 == pht_widx ? pht_501 : _GEN_1045; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1047 = 9'h1f6 == pht_widx ? pht_502 : _GEN_1046; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1048 = 9'h1f7 == pht_widx ? pht_503 : _GEN_1047; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1049 = 9'h1f8 == pht_widx ? pht_504 : _GEN_1048; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1050 = 9'h1f9 == pht_widx ? pht_505 : _GEN_1049; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1051 = 9'h1fa == pht_widx ? pht_506 : _GEN_1050; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1052 = 9'h1fb == pht_widx ? pht_507 : _GEN_1051; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1053 = 9'h1fc == pht_widx ? pht_508 : _GEN_1052; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1054 = 9'h1fd == pht_widx ? pht_509 : _GEN_1053; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1055 = 9'h1fe == pht_widx ? pht_510 : _GEN_1054; // @[Mux.scala 81:{61,61}]
  wire [1:0] _GEN_1056 = 9'h1ff == pht_widx ? pht_511 : _GEN_1055; // @[Mux.scala 81:{61,61}]
  wire [1:0] _pht_T_5 = 2'h1 == _GEN_1056 ? _pht_T_1 : {{1'd0}, io_jmp_packet_bp_taken}; // @[Mux.scala 81:58]
  wire [1:0] _pht_T_7 = 2'h2 == _GEN_1056 ? _pht_T_2 : _pht_T_5; // @[Mux.scala 81:58]
  wire [3:0] _GEN_2085 = btb_1_valid & btb_1_tag == io_jmp_packet_bp_pc[38:2] ? 4'h1 : 4'h0; // @[BPU.scala 71:81 73:20]
  wire [3:0] _GEN_2087 = btb_2_valid & btb_2_tag == io_jmp_packet_bp_pc[38:2] ? 4'h2 : _GEN_2085; // @[BPU.scala 71:81 73:20]
  wire [3:0] _GEN_2089 = btb_3_valid & btb_3_tag == io_jmp_packet_bp_pc[38:2] ? 4'h3 : _GEN_2087; // @[BPU.scala 71:81 73:20]
  wire [3:0] _GEN_2091 = btb_4_valid & btb_4_tag == io_jmp_packet_bp_pc[38:2] ? 4'h4 : _GEN_2089; // @[BPU.scala 71:81 73:20]
  wire [3:0] _GEN_2093 = btb_5_valid & btb_5_tag == io_jmp_packet_bp_pc[38:2] ? 4'h5 : _GEN_2091; // @[BPU.scala 71:81 73:20]
  wire [3:0] _GEN_2095 = btb_6_valid & btb_6_tag == io_jmp_packet_bp_pc[38:2] ? 4'h6 : _GEN_2093; // @[BPU.scala 71:81 73:20]
  wire [3:0] _GEN_2097 = btb_7_valid & btb_7_tag == io_jmp_packet_bp_pc[38:2] ? 4'h7 : _GEN_2095; // @[BPU.scala 71:81 73:20]
  wire [3:0] _GEN_2099 = btb_8_valid & btb_8_tag == io_jmp_packet_bp_pc[38:2] ? 4'h8 : _GEN_2097; // @[BPU.scala 71:81 73:20]
  wire  _GEN_2100 = btb_9_valid & btb_9_tag == io_jmp_packet_bp_pc[38:2] | (btb_8_valid & btb_8_tag ==
    io_jmp_packet_bp_pc[38:2] | (btb_7_valid & btb_7_tag == io_jmp_packet_bp_pc[38:2] | (btb_6_valid & btb_6_tag ==
    io_jmp_packet_bp_pc[38:2] | (btb_5_valid & btb_5_tag == io_jmp_packet_bp_pc[38:2] | (btb_4_valid & btb_4_tag ==
    io_jmp_packet_bp_pc[38:2] | (btb_3_valid & btb_3_tag == io_jmp_packet_bp_pc[38:2] | (btb_2_valid & btb_2_tag ==
    io_jmp_packet_bp_pc[38:2] | (btb_1_valid & btb_1_tag == io_jmp_packet_bp_pc[38:2] | btb_0_valid & btb_0_tag ==
    io_jmp_packet_bp_pc[38:2])))))))); // @[BPU.scala 71:81 72:20]
  wire [3:0] _GEN_2101 = btb_9_valid & btb_9_tag == io_jmp_packet_bp_pc[38:2] ? 4'h9 : _GEN_2099; // @[BPU.scala 71:81 73:20]
  wire [3:0] _GEN_2103 = btb_10_valid & btb_10_tag == io_jmp_packet_bp_pc[38:2] ? 4'ha : _GEN_2101; // @[BPU.scala 71:81 73:20]
  wire [3:0] _GEN_2105 = btb_11_valid & btb_11_tag == io_jmp_packet_bp_pc[38:2] ? 4'hb : _GEN_2103; // @[BPU.scala 71:81 73:20]
  wire [3:0] _GEN_2107 = btb_12_valid & btb_12_tag == io_jmp_packet_bp_pc[38:2] ? 4'hc : _GEN_2105; // @[BPU.scala 71:81 73:20]
  wire [3:0] _GEN_2109 = btb_13_valid & btb_13_tag == io_jmp_packet_bp_pc[38:2] ? 4'hd : _GEN_2107; // @[BPU.scala 71:81 73:20]
  wire [3:0] _GEN_2111 = btb_14_valid & btb_14_tag == io_jmp_packet_bp_pc[38:2] ? 4'he : _GEN_2109; // @[BPU.scala 71:81 73:20]
  wire  btb_whit = btb_15_valid & btb_15_tag == io_jmp_packet_bp_pc[38:2] | (btb_14_valid & btb_14_tag ==
    io_jmp_packet_bp_pc[38:2] | (btb_13_valid & btb_13_tag == io_jmp_packet_bp_pc[38:2] | (btb_12_valid & btb_12_tag ==
    io_jmp_packet_bp_pc[38:2] | (btb_11_valid & btb_11_tag == io_jmp_packet_bp_pc[38:2] | (btb_10_valid & btb_10_tag ==
    io_jmp_packet_bp_pc[38:2] | _GEN_2100))))); // @[BPU.scala 71:81 72:20]
  wire [3:0] btb_whit_way = btb_15_valid & btb_15_tag == io_jmp_packet_bp_pc[38:2] ? 4'hf : _GEN_2111; // @[BPU.scala 71:81 73:20]
  wire [3:0] _btb_replace_idx_T = {btb_replace_idx_prng_io_out_3,btb_replace_idx_prng_io_out_2,
    btb_replace_idx_prng_io_out_1,btb_replace_idx_prng_io_out_0}; // @[PRNG.scala 95:17]
  wire [3:0] btb_replace_idx = btb_whit ? btb_whit_way : _btb_replace_idx_T; // @[BPU.scala 77:25]
  wire  _GEN_2114 = 4'h0 == btb_replace_idx | btb_0_valid; // @[BPU.scala 28:20 79:{33,33}]
  wire  _GEN_2115 = 4'h1 == btb_replace_idx | btb_1_valid; // @[BPU.scala 28:20 79:{33,33}]
  wire  _GEN_2116 = 4'h2 == btb_replace_idx | btb_2_valid; // @[BPU.scala 28:20 79:{33,33}]
  wire  _GEN_2117 = 4'h3 == btb_replace_idx | btb_3_valid; // @[BPU.scala 28:20 79:{33,33}]
  wire  _GEN_2118 = 4'h4 == btb_replace_idx | btb_4_valid; // @[BPU.scala 28:20 79:{33,33}]
  wire  _GEN_2119 = 4'h5 == btb_replace_idx | btb_5_valid; // @[BPU.scala 28:20 79:{33,33}]
  wire  _GEN_2120 = 4'h6 == btb_replace_idx | btb_6_valid; // @[BPU.scala 28:20 79:{33,33}]
  wire  _GEN_2121 = 4'h7 == btb_replace_idx | btb_7_valid; // @[BPU.scala 28:20 79:{33,33}]
  wire  _GEN_2122 = 4'h8 == btb_replace_idx | btb_8_valid; // @[BPU.scala 28:20 79:{33,33}]
  wire  _GEN_2123 = 4'h9 == btb_replace_idx | btb_9_valid; // @[BPU.scala 28:20 79:{33,33}]
  wire  _GEN_2124 = 4'ha == btb_replace_idx | btb_10_valid; // @[BPU.scala 28:20 79:{33,33}]
  wire  _GEN_2125 = 4'hb == btb_replace_idx | btb_11_valid; // @[BPU.scala 28:20 79:{33,33}]
  wire  _GEN_2126 = 4'hc == btb_replace_idx | btb_12_valid; // @[BPU.scala 28:20 79:{33,33}]
  wire  _GEN_2127 = 4'hd == btb_replace_idx | btb_13_valid; // @[BPU.scala 28:20 79:{33,33}]
  wire  _GEN_2128 = 4'he == btb_replace_idx | btb_14_valid; // @[BPU.scala 28:20 79:{33,33}]
  wire  _GEN_2129 = 4'hf == btb_replace_idx | btb_15_valid; // @[BPU.scala 28:20 79:{33,33}]
  MaxPeriodFibonacciLFSR btb_replace_idx_prng ( // @[PRNG.scala 91:22]
    .clock(btb_replace_idx_prng_clock),
    .reset(btb_replace_idx_prng_reset),
    .io_out_0(btb_replace_idx_prng_io_out_0),
    .io_out_1(btb_replace_idx_prng_io_out_1),
    .io_out_2(btb_replace_idx_prng_io_out_2),
    .io_out_3(btb_replace_idx_prng_io_out_3)
  );
  assign io_out = pht_taken & btb_rhit ? _io_out_T_6 : _io_out_T_1; // @[BPU.scala 46:10 47:31 48:12]
  assign btb_replace_idx_prng_clock = clock;
  assign btb_replace_idx_prng_reset = reset;
  always @(posedge clock) begin
    if (reset) begin // @[BPU.scala 26:20]
      ghr <= 9'h0; // @[BPU.scala 26:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      ghr <= {{1'd0}, _ghr_T_1}; // @[BPU.scala 54:9]
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_0 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h0 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_0 <= _pht_T_3;
        end else begin
          pht_0 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_1 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_1 <= _pht_T_3;
        end else begin
          pht_1 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_2 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h2 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_2 <= _pht_T_3;
        end else begin
          pht_2 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_3 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h3 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_3 <= _pht_T_3;
        end else begin
          pht_3 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_4 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h4 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_4 <= _pht_T_3;
        end else begin
          pht_4 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_5 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h5 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_5 <= _pht_T_3;
        end else begin
          pht_5 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_6 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h6 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_6 <= _pht_T_3;
        end else begin
          pht_6 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_7 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h7 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_7 <= _pht_T_3;
        end else begin
          pht_7 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_8 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h8 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_8 <= _pht_T_3;
        end else begin
          pht_8 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_9 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h9 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_9 <= _pht_T_3;
        end else begin
          pht_9 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_10 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'ha == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_10 <= _pht_T_3;
        end else begin
          pht_10 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_11 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hb == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_11 <= _pht_T_3;
        end else begin
          pht_11 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_12 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hc == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_12 <= _pht_T_3;
        end else begin
          pht_12 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_13 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hd == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_13 <= _pht_T_3;
        end else begin
          pht_13 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_14 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'he == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_14 <= _pht_T_3;
        end else begin
          pht_14 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_15 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hf == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_15 <= _pht_T_3;
        end else begin
          pht_15 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_16 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h10 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_16 <= _pht_T_3;
        end else begin
          pht_16 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_17 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h11 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_17 <= _pht_T_3;
        end else begin
          pht_17 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_18 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h12 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_18 <= _pht_T_3;
        end else begin
          pht_18 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_19 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h13 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_19 <= _pht_T_3;
        end else begin
          pht_19 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_20 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h14 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_20 <= _pht_T_3;
        end else begin
          pht_20 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_21 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h15 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_21 <= _pht_T_3;
        end else begin
          pht_21 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_22 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h16 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_22 <= _pht_T_3;
        end else begin
          pht_22 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_23 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h17 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_23 <= _pht_T_3;
        end else begin
          pht_23 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_24 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h18 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_24 <= _pht_T_3;
        end else begin
          pht_24 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_25 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h19 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_25 <= _pht_T_3;
        end else begin
          pht_25 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_26 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1a == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_26 <= _pht_T_3;
        end else begin
          pht_26 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_27 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1b == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_27 <= _pht_T_3;
        end else begin
          pht_27 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_28 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1c == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_28 <= _pht_T_3;
        end else begin
          pht_28 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_29 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1d == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_29 <= _pht_T_3;
        end else begin
          pht_29 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_30 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1e == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_30 <= _pht_T_3;
        end else begin
          pht_30 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_31 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1f == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_31 <= _pht_T_3;
        end else begin
          pht_31 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_32 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h20 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_32 <= _pht_T_3;
        end else begin
          pht_32 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_33 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h21 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_33 <= _pht_T_3;
        end else begin
          pht_33 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_34 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h22 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_34 <= _pht_T_3;
        end else begin
          pht_34 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_35 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h23 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_35 <= _pht_T_3;
        end else begin
          pht_35 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_36 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h24 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_36 <= _pht_T_3;
        end else begin
          pht_36 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_37 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h25 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_37 <= _pht_T_3;
        end else begin
          pht_37 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_38 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h26 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_38 <= _pht_T_3;
        end else begin
          pht_38 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_39 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h27 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_39 <= _pht_T_3;
        end else begin
          pht_39 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_40 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h28 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_40 <= _pht_T_3;
        end else begin
          pht_40 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_41 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h29 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_41 <= _pht_T_3;
        end else begin
          pht_41 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_42 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h2a == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_42 <= _pht_T_3;
        end else begin
          pht_42 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_43 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h2b == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_43 <= _pht_T_3;
        end else begin
          pht_43 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_44 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h2c == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_44 <= _pht_T_3;
        end else begin
          pht_44 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_45 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h2d == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_45 <= _pht_T_3;
        end else begin
          pht_45 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_46 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h2e == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_46 <= _pht_T_3;
        end else begin
          pht_46 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_47 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h2f == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_47 <= _pht_T_3;
        end else begin
          pht_47 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_48 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h30 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_48 <= _pht_T_3;
        end else begin
          pht_48 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_49 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h31 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_49 <= _pht_T_3;
        end else begin
          pht_49 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_50 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h32 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_50 <= _pht_T_3;
        end else begin
          pht_50 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_51 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h33 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_51 <= _pht_T_3;
        end else begin
          pht_51 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_52 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h34 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_52 <= _pht_T_3;
        end else begin
          pht_52 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_53 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h35 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_53 <= _pht_T_3;
        end else begin
          pht_53 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_54 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h36 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_54 <= _pht_T_3;
        end else begin
          pht_54 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_55 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h37 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_55 <= _pht_T_3;
        end else begin
          pht_55 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_56 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h38 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_56 <= _pht_T_3;
        end else begin
          pht_56 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_57 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h39 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_57 <= _pht_T_3;
        end else begin
          pht_57 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_58 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h3a == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_58 <= _pht_T_3;
        end else begin
          pht_58 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_59 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h3b == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_59 <= _pht_T_3;
        end else begin
          pht_59 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_60 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h3c == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_60 <= _pht_T_3;
        end else begin
          pht_60 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_61 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h3d == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_61 <= _pht_T_3;
        end else begin
          pht_61 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_62 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h3e == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_62 <= _pht_T_3;
        end else begin
          pht_62 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_63 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h3f == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_63 <= _pht_T_3;
        end else begin
          pht_63 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_64 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h40 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_64 <= _pht_T_3;
        end else begin
          pht_64 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_65 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h41 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_65 <= _pht_T_3;
        end else begin
          pht_65 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_66 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h42 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_66 <= _pht_T_3;
        end else begin
          pht_66 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_67 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h43 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_67 <= _pht_T_3;
        end else begin
          pht_67 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_68 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h44 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_68 <= _pht_T_3;
        end else begin
          pht_68 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_69 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h45 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_69 <= _pht_T_3;
        end else begin
          pht_69 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_70 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h46 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_70 <= _pht_T_3;
        end else begin
          pht_70 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_71 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h47 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_71 <= _pht_T_3;
        end else begin
          pht_71 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_72 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h48 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_72 <= _pht_T_3;
        end else begin
          pht_72 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_73 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h49 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_73 <= _pht_T_3;
        end else begin
          pht_73 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_74 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h4a == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_74 <= _pht_T_3;
        end else begin
          pht_74 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_75 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h4b == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_75 <= _pht_T_3;
        end else begin
          pht_75 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_76 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h4c == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_76 <= _pht_T_3;
        end else begin
          pht_76 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_77 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h4d == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_77 <= _pht_T_3;
        end else begin
          pht_77 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_78 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h4e == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_78 <= _pht_T_3;
        end else begin
          pht_78 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_79 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h4f == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_79 <= _pht_T_3;
        end else begin
          pht_79 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_80 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h50 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_80 <= _pht_T_3;
        end else begin
          pht_80 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_81 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h51 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_81 <= _pht_T_3;
        end else begin
          pht_81 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_82 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h52 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_82 <= _pht_T_3;
        end else begin
          pht_82 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_83 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h53 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_83 <= _pht_T_3;
        end else begin
          pht_83 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_84 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h54 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_84 <= _pht_T_3;
        end else begin
          pht_84 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_85 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h55 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_85 <= _pht_T_3;
        end else begin
          pht_85 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_86 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h56 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_86 <= _pht_T_3;
        end else begin
          pht_86 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_87 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h57 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_87 <= _pht_T_3;
        end else begin
          pht_87 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_88 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h58 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_88 <= _pht_T_3;
        end else begin
          pht_88 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_89 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h59 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_89 <= _pht_T_3;
        end else begin
          pht_89 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_90 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h5a == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_90 <= _pht_T_3;
        end else begin
          pht_90 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_91 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h5b == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_91 <= _pht_T_3;
        end else begin
          pht_91 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_92 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h5c == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_92 <= _pht_T_3;
        end else begin
          pht_92 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_93 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h5d == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_93 <= _pht_T_3;
        end else begin
          pht_93 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_94 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h5e == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_94 <= _pht_T_3;
        end else begin
          pht_94 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_95 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h5f == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_95 <= _pht_T_3;
        end else begin
          pht_95 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_96 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h60 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_96 <= _pht_T_3;
        end else begin
          pht_96 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_97 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h61 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_97 <= _pht_T_3;
        end else begin
          pht_97 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_98 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h62 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_98 <= _pht_T_3;
        end else begin
          pht_98 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_99 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h63 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_99 <= _pht_T_3;
        end else begin
          pht_99 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_100 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h64 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_100 <= _pht_T_3;
        end else begin
          pht_100 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_101 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h65 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_101 <= _pht_T_3;
        end else begin
          pht_101 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_102 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h66 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_102 <= _pht_T_3;
        end else begin
          pht_102 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_103 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h67 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_103 <= _pht_T_3;
        end else begin
          pht_103 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_104 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h68 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_104 <= _pht_T_3;
        end else begin
          pht_104 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_105 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h69 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_105 <= _pht_T_3;
        end else begin
          pht_105 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_106 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h6a == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_106 <= _pht_T_3;
        end else begin
          pht_106 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_107 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h6b == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_107 <= _pht_T_3;
        end else begin
          pht_107 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_108 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h6c == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_108 <= _pht_T_3;
        end else begin
          pht_108 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_109 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h6d == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_109 <= _pht_T_3;
        end else begin
          pht_109 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_110 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h6e == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_110 <= _pht_T_3;
        end else begin
          pht_110 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_111 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h6f == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_111 <= _pht_T_3;
        end else begin
          pht_111 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_112 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h70 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_112 <= _pht_T_3;
        end else begin
          pht_112 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_113 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h71 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_113 <= _pht_T_3;
        end else begin
          pht_113 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_114 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h72 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_114 <= _pht_T_3;
        end else begin
          pht_114 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_115 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h73 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_115 <= _pht_T_3;
        end else begin
          pht_115 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_116 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h74 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_116 <= _pht_T_3;
        end else begin
          pht_116 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_117 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h75 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_117 <= _pht_T_3;
        end else begin
          pht_117 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_118 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h76 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_118 <= _pht_T_3;
        end else begin
          pht_118 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_119 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h77 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_119 <= _pht_T_3;
        end else begin
          pht_119 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_120 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h78 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_120 <= _pht_T_3;
        end else begin
          pht_120 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_121 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h79 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_121 <= _pht_T_3;
        end else begin
          pht_121 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_122 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h7a == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_122 <= _pht_T_3;
        end else begin
          pht_122 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_123 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h7b == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_123 <= _pht_T_3;
        end else begin
          pht_123 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_124 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h7c == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_124 <= _pht_T_3;
        end else begin
          pht_124 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_125 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h7d == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_125 <= _pht_T_3;
        end else begin
          pht_125 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_126 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h7e == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_126 <= _pht_T_3;
        end else begin
          pht_126 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_127 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h7f == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_127 <= _pht_T_3;
        end else begin
          pht_127 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_128 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h80 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_128 <= _pht_T_3;
        end else begin
          pht_128 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_129 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h81 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_129 <= _pht_T_3;
        end else begin
          pht_129 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_130 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h82 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_130 <= _pht_T_3;
        end else begin
          pht_130 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_131 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h83 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_131 <= _pht_T_3;
        end else begin
          pht_131 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_132 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h84 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_132 <= _pht_T_3;
        end else begin
          pht_132 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_133 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h85 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_133 <= _pht_T_3;
        end else begin
          pht_133 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_134 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h86 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_134 <= _pht_T_3;
        end else begin
          pht_134 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_135 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h87 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_135 <= _pht_T_3;
        end else begin
          pht_135 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_136 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h88 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_136 <= _pht_T_3;
        end else begin
          pht_136 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_137 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h89 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_137 <= _pht_T_3;
        end else begin
          pht_137 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_138 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h8a == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_138 <= _pht_T_3;
        end else begin
          pht_138 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_139 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h8b == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_139 <= _pht_T_3;
        end else begin
          pht_139 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_140 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h8c == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_140 <= _pht_T_3;
        end else begin
          pht_140 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_141 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h8d == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_141 <= _pht_T_3;
        end else begin
          pht_141 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_142 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h8e == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_142 <= _pht_T_3;
        end else begin
          pht_142 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_143 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h8f == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_143 <= _pht_T_3;
        end else begin
          pht_143 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_144 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h90 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_144 <= _pht_T_3;
        end else begin
          pht_144 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_145 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h91 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_145 <= _pht_T_3;
        end else begin
          pht_145 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_146 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h92 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_146 <= _pht_T_3;
        end else begin
          pht_146 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_147 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h93 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_147 <= _pht_T_3;
        end else begin
          pht_147 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_148 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h94 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_148 <= _pht_T_3;
        end else begin
          pht_148 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_149 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h95 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_149 <= _pht_T_3;
        end else begin
          pht_149 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_150 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h96 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_150 <= _pht_T_3;
        end else begin
          pht_150 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_151 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h97 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_151 <= _pht_T_3;
        end else begin
          pht_151 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_152 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h98 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_152 <= _pht_T_3;
        end else begin
          pht_152 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_153 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h99 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_153 <= _pht_T_3;
        end else begin
          pht_153 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_154 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h9a == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_154 <= _pht_T_3;
        end else begin
          pht_154 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_155 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h9b == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_155 <= _pht_T_3;
        end else begin
          pht_155 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_156 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h9c == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_156 <= _pht_T_3;
        end else begin
          pht_156 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_157 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h9d == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_157 <= _pht_T_3;
        end else begin
          pht_157 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_158 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h9e == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_158 <= _pht_T_3;
        end else begin
          pht_158 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_159 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h9f == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_159 <= _pht_T_3;
        end else begin
          pht_159 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_160 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'ha0 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_160 <= _pht_T_3;
        end else begin
          pht_160 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_161 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'ha1 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_161 <= _pht_T_3;
        end else begin
          pht_161 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_162 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'ha2 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_162 <= _pht_T_3;
        end else begin
          pht_162 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_163 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'ha3 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_163 <= _pht_T_3;
        end else begin
          pht_163 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_164 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'ha4 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_164 <= _pht_T_3;
        end else begin
          pht_164 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_165 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'ha5 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_165 <= _pht_T_3;
        end else begin
          pht_165 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_166 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'ha6 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_166 <= _pht_T_3;
        end else begin
          pht_166 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_167 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'ha7 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_167 <= _pht_T_3;
        end else begin
          pht_167 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_168 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'ha8 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_168 <= _pht_T_3;
        end else begin
          pht_168 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_169 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'ha9 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_169 <= _pht_T_3;
        end else begin
          pht_169 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_170 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'haa == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_170 <= _pht_T_3;
        end else begin
          pht_170 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_171 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hab == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_171 <= _pht_T_3;
        end else begin
          pht_171 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_172 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hac == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_172 <= _pht_T_3;
        end else begin
          pht_172 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_173 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'had == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_173 <= _pht_T_3;
        end else begin
          pht_173 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_174 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hae == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_174 <= _pht_T_3;
        end else begin
          pht_174 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_175 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'haf == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_175 <= _pht_T_3;
        end else begin
          pht_175 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_176 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hb0 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_176 <= _pht_T_3;
        end else begin
          pht_176 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_177 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hb1 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_177 <= _pht_T_3;
        end else begin
          pht_177 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_178 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hb2 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_178 <= _pht_T_3;
        end else begin
          pht_178 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_179 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hb3 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_179 <= _pht_T_3;
        end else begin
          pht_179 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_180 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hb4 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_180 <= _pht_T_3;
        end else begin
          pht_180 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_181 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hb5 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_181 <= _pht_T_3;
        end else begin
          pht_181 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_182 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hb6 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_182 <= _pht_T_3;
        end else begin
          pht_182 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_183 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hb7 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_183 <= _pht_T_3;
        end else begin
          pht_183 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_184 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hb8 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_184 <= _pht_T_3;
        end else begin
          pht_184 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_185 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hb9 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_185 <= _pht_T_3;
        end else begin
          pht_185 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_186 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hba == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_186 <= _pht_T_3;
        end else begin
          pht_186 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_187 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hbb == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_187 <= _pht_T_3;
        end else begin
          pht_187 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_188 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hbc == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_188 <= _pht_T_3;
        end else begin
          pht_188 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_189 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hbd == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_189 <= _pht_T_3;
        end else begin
          pht_189 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_190 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hbe == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_190 <= _pht_T_3;
        end else begin
          pht_190 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_191 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hbf == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_191 <= _pht_T_3;
        end else begin
          pht_191 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_192 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hc0 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_192 <= _pht_T_3;
        end else begin
          pht_192 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_193 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hc1 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_193 <= _pht_T_3;
        end else begin
          pht_193 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_194 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hc2 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_194 <= _pht_T_3;
        end else begin
          pht_194 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_195 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hc3 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_195 <= _pht_T_3;
        end else begin
          pht_195 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_196 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hc4 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_196 <= _pht_T_3;
        end else begin
          pht_196 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_197 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hc5 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_197 <= _pht_T_3;
        end else begin
          pht_197 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_198 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hc6 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_198 <= _pht_T_3;
        end else begin
          pht_198 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_199 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hc7 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_199 <= _pht_T_3;
        end else begin
          pht_199 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_200 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hc8 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_200 <= _pht_T_3;
        end else begin
          pht_200 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_201 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hc9 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_201 <= _pht_T_3;
        end else begin
          pht_201 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_202 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hca == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_202 <= _pht_T_3;
        end else begin
          pht_202 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_203 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hcb == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_203 <= _pht_T_3;
        end else begin
          pht_203 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_204 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hcc == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_204 <= _pht_T_3;
        end else begin
          pht_204 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_205 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hcd == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_205 <= _pht_T_3;
        end else begin
          pht_205 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_206 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hce == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_206 <= _pht_T_3;
        end else begin
          pht_206 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_207 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hcf == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_207 <= _pht_T_3;
        end else begin
          pht_207 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_208 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hd0 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_208 <= _pht_T_3;
        end else begin
          pht_208 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_209 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hd1 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_209 <= _pht_T_3;
        end else begin
          pht_209 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_210 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hd2 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_210 <= _pht_T_3;
        end else begin
          pht_210 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_211 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hd3 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_211 <= _pht_T_3;
        end else begin
          pht_211 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_212 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hd4 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_212 <= _pht_T_3;
        end else begin
          pht_212 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_213 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hd5 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_213 <= _pht_T_3;
        end else begin
          pht_213 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_214 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hd6 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_214 <= _pht_T_3;
        end else begin
          pht_214 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_215 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hd7 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_215 <= _pht_T_3;
        end else begin
          pht_215 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_216 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hd8 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_216 <= _pht_T_3;
        end else begin
          pht_216 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_217 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hd9 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_217 <= _pht_T_3;
        end else begin
          pht_217 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_218 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hda == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_218 <= _pht_T_3;
        end else begin
          pht_218 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_219 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hdb == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_219 <= _pht_T_3;
        end else begin
          pht_219 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_220 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hdc == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_220 <= _pht_T_3;
        end else begin
          pht_220 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_221 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hdd == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_221 <= _pht_T_3;
        end else begin
          pht_221 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_222 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hde == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_222 <= _pht_T_3;
        end else begin
          pht_222 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_223 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hdf == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_223 <= _pht_T_3;
        end else begin
          pht_223 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_224 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'he0 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_224 <= _pht_T_3;
        end else begin
          pht_224 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_225 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'he1 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_225 <= _pht_T_3;
        end else begin
          pht_225 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_226 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'he2 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_226 <= _pht_T_3;
        end else begin
          pht_226 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_227 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'he3 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_227 <= _pht_T_3;
        end else begin
          pht_227 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_228 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'he4 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_228 <= _pht_T_3;
        end else begin
          pht_228 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_229 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'he5 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_229 <= _pht_T_3;
        end else begin
          pht_229 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_230 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'he6 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_230 <= _pht_T_3;
        end else begin
          pht_230 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_231 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'he7 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_231 <= _pht_T_3;
        end else begin
          pht_231 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_232 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'he8 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_232 <= _pht_T_3;
        end else begin
          pht_232 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_233 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'he9 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_233 <= _pht_T_3;
        end else begin
          pht_233 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_234 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hea == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_234 <= _pht_T_3;
        end else begin
          pht_234 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_235 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'heb == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_235 <= _pht_T_3;
        end else begin
          pht_235 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_236 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hec == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_236 <= _pht_T_3;
        end else begin
          pht_236 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_237 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hed == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_237 <= _pht_T_3;
        end else begin
          pht_237 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_238 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hee == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_238 <= _pht_T_3;
        end else begin
          pht_238 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_239 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hef == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_239 <= _pht_T_3;
        end else begin
          pht_239 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_240 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hf0 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_240 <= _pht_T_3;
        end else begin
          pht_240 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_241 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hf1 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_241 <= _pht_T_3;
        end else begin
          pht_241 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_242 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hf2 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_242 <= _pht_T_3;
        end else begin
          pht_242 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_243 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hf3 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_243 <= _pht_T_3;
        end else begin
          pht_243 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_244 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hf4 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_244 <= _pht_T_3;
        end else begin
          pht_244 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_245 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hf5 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_245 <= _pht_T_3;
        end else begin
          pht_245 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_246 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hf6 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_246 <= _pht_T_3;
        end else begin
          pht_246 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_247 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hf7 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_247 <= _pht_T_3;
        end else begin
          pht_247 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_248 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hf8 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_248 <= _pht_T_3;
        end else begin
          pht_248 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_249 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hf9 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_249 <= _pht_T_3;
        end else begin
          pht_249 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_250 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hfa == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_250 <= _pht_T_3;
        end else begin
          pht_250 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_251 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hfb == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_251 <= _pht_T_3;
        end else begin
          pht_251 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_252 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hfc == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_252 <= _pht_T_3;
        end else begin
          pht_252 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_253 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hfd == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_253 <= _pht_T_3;
        end else begin
          pht_253 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_254 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hfe == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_254 <= _pht_T_3;
        end else begin
          pht_254 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_255 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'hff == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_255 <= _pht_T_3;
        end else begin
          pht_255 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_256 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h100 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_256 <= _pht_T_3;
        end else begin
          pht_256 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_257 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h101 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_257 <= _pht_T_3;
        end else begin
          pht_257 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_258 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h102 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_258 <= _pht_T_3;
        end else begin
          pht_258 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_259 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h103 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_259 <= _pht_T_3;
        end else begin
          pht_259 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_260 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h104 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_260 <= _pht_T_3;
        end else begin
          pht_260 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_261 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h105 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_261 <= _pht_T_3;
        end else begin
          pht_261 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_262 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h106 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_262 <= _pht_T_3;
        end else begin
          pht_262 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_263 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h107 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_263 <= _pht_T_3;
        end else begin
          pht_263 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_264 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h108 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_264 <= _pht_T_3;
        end else begin
          pht_264 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_265 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h109 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_265 <= _pht_T_3;
        end else begin
          pht_265 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_266 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h10a == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_266 <= _pht_T_3;
        end else begin
          pht_266 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_267 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h10b == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_267 <= _pht_T_3;
        end else begin
          pht_267 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_268 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h10c == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_268 <= _pht_T_3;
        end else begin
          pht_268 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_269 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h10d == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_269 <= _pht_T_3;
        end else begin
          pht_269 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_270 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h10e == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_270 <= _pht_T_3;
        end else begin
          pht_270 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_271 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h10f == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_271 <= _pht_T_3;
        end else begin
          pht_271 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_272 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h110 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_272 <= _pht_T_3;
        end else begin
          pht_272 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_273 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h111 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_273 <= _pht_T_3;
        end else begin
          pht_273 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_274 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h112 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_274 <= _pht_T_3;
        end else begin
          pht_274 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_275 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h113 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_275 <= _pht_T_3;
        end else begin
          pht_275 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_276 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h114 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_276 <= _pht_T_3;
        end else begin
          pht_276 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_277 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h115 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_277 <= _pht_T_3;
        end else begin
          pht_277 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_278 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h116 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_278 <= _pht_T_3;
        end else begin
          pht_278 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_279 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h117 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_279 <= _pht_T_3;
        end else begin
          pht_279 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_280 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h118 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_280 <= _pht_T_3;
        end else begin
          pht_280 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_281 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h119 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_281 <= _pht_T_3;
        end else begin
          pht_281 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_282 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h11a == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_282 <= _pht_T_3;
        end else begin
          pht_282 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_283 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h11b == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_283 <= _pht_T_3;
        end else begin
          pht_283 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_284 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h11c == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_284 <= _pht_T_3;
        end else begin
          pht_284 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_285 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h11d == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_285 <= _pht_T_3;
        end else begin
          pht_285 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_286 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h11e == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_286 <= _pht_T_3;
        end else begin
          pht_286 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_287 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h11f == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_287 <= _pht_T_3;
        end else begin
          pht_287 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_288 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h120 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_288 <= _pht_T_3;
        end else begin
          pht_288 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_289 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h121 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_289 <= _pht_T_3;
        end else begin
          pht_289 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_290 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h122 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_290 <= _pht_T_3;
        end else begin
          pht_290 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_291 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h123 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_291 <= _pht_T_3;
        end else begin
          pht_291 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_292 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h124 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_292 <= _pht_T_3;
        end else begin
          pht_292 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_293 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h125 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_293 <= _pht_T_3;
        end else begin
          pht_293 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_294 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h126 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_294 <= _pht_T_3;
        end else begin
          pht_294 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_295 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h127 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_295 <= _pht_T_3;
        end else begin
          pht_295 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_296 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h128 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_296 <= _pht_T_3;
        end else begin
          pht_296 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_297 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h129 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_297 <= _pht_T_3;
        end else begin
          pht_297 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_298 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h12a == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_298 <= _pht_T_3;
        end else begin
          pht_298 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_299 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h12b == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_299 <= _pht_T_3;
        end else begin
          pht_299 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_300 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h12c == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_300 <= _pht_T_3;
        end else begin
          pht_300 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_301 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h12d == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_301 <= _pht_T_3;
        end else begin
          pht_301 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_302 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h12e == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_302 <= _pht_T_3;
        end else begin
          pht_302 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_303 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h12f == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_303 <= _pht_T_3;
        end else begin
          pht_303 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_304 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h130 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_304 <= _pht_T_3;
        end else begin
          pht_304 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_305 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h131 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_305 <= _pht_T_3;
        end else begin
          pht_305 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_306 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h132 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_306 <= _pht_T_3;
        end else begin
          pht_306 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_307 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h133 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_307 <= _pht_T_3;
        end else begin
          pht_307 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_308 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h134 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_308 <= _pht_T_3;
        end else begin
          pht_308 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_309 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h135 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_309 <= _pht_T_3;
        end else begin
          pht_309 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_310 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h136 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_310 <= _pht_T_3;
        end else begin
          pht_310 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_311 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h137 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_311 <= _pht_T_3;
        end else begin
          pht_311 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_312 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h138 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_312 <= _pht_T_3;
        end else begin
          pht_312 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_313 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h139 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_313 <= _pht_T_3;
        end else begin
          pht_313 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_314 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h13a == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_314 <= _pht_T_3;
        end else begin
          pht_314 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_315 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h13b == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_315 <= _pht_T_3;
        end else begin
          pht_315 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_316 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h13c == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_316 <= _pht_T_3;
        end else begin
          pht_316 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_317 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h13d == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_317 <= _pht_T_3;
        end else begin
          pht_317 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_318 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h13e == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_318 <= _pht_T_3;
        end else begin
          pht_318 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_319 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h13f == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_319 <= _pht_T_3;
        end else begin
          pht_319 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_320 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h140 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_320 <= _pht_T_3;
        end else begin
          pht_320 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_321 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h141 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_321 <= _pht_T_3;
        end else begin
          pht_321 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_322 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h142 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_322 <= _pht_T_3;
        end else begin
          pht_322 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_323 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h143 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_323 <= _pht_T_3;
        end else begin
          pht_323 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_324 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h144 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_324 <= _pht_T_3;
        end else begin
          pht_324 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_325 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h145 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_325 <= _pht_T_3;
        end else begin
          pht_325 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_326 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h146 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_326 <= _pht_T_3;
        end else begin
          pht_326 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_327 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h147 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_327 <= _pht_T_3;
        end else begin
          pht_327 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_328 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h148 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_328 <= _pht_T_3;
        end else begin
          pht_328 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_329 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h149 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_329 <= _pht_T_3;
        end else begin
          pht_329 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_330 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h14a == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_330 <= _pht_T_3;
        end else begin
          pht_330 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_331 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h14b == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_331 <= _pht_T_3;
        end else begin
          pht_331 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_332 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h14c == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_332 <= _pht_T_3;
        end else begin
          pht_332 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_333 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h14d == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_333 <= _pht_T_3;
        end else begin
          pht_333 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_334 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h14e == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_334 <= _pht_T_3;
        end else begin
          pht_334 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_335 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h14f == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_335 <= _pht_T_3;
        end else begin
          pht_335 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_336 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h150 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_336 <= _pht_T_3;
        end else begin
          pht_336 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_337 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h151 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_337 <= _pht_T_3;
        end else begin
          pht_337 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_338 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h152 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_338 <= _pht_T_3;
        end else begin
          pht_338 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_339 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h153 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_339 <= _pht_T_3;
        end else begin
          pht_339 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_340 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h154 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_340 <= _pht_T_3;
        end else begin
          pht_340 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_341 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h155 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_341 <= _pht_T_3;
        end else begin
          pht_341 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_342 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h156 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_342 <= _pht_T_3;
        end else begin
          pht_342 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_343 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h157 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_343 <= _pht_T_3;
        end else begin
          pht_343 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_344 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h158 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_344 <= _pht_T_3;
        end else begin
          pht_344 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_345 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h159 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_345 <= _pht_T_3;
        end else begin
          pht_345 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_346 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h15a == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_346 <= _pht_T_3;
        end else begin
          pht_346 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_347 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h15b == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_347 <= _pht_T_3;
        end else begin
          pht_347 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_348 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h15c == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_348 <= _pht_T_3;
        end else begin
          pht_348 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_349 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h15d == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_349 <= _pht_T_3;
        end else begin
          pht_349 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_350 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h15e == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_350 <= _pht_T_3;
        end else begin
          pht_350 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_351 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h15f == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_351 <= _pht_T_3;
        end else begin
          pht_351 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_352 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h160 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_352 <= _pht_T_3;
        end else begin
          pht_352 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_353 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h161 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_353 <= _pht_T_3;
        end else begin
          pht_353 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_354 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h162 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_354 <= _pht_T_3;
        end else begin
          pht_354 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_355 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h163 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_355 <= _pht_T_3;
        end else begin
          pht_355 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_356 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h164 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_356 <= _pht_T_3;
        end else begin
          pht_356 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_357 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h165 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_357 <= _pht_T_3;
        end else begin
          pht_357 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_358 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h166 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_358 <= _pht_T_3;
        end else begin
          pht_358 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_359 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h167 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_359 <= _pht_T_3;
        end else begin
          pht_359 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_360 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h168 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_360 <= _pht_T_3;
        end else begin
          pht_360 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_361 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h169 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_361 <= _pht_T_3;
        end else begin
          pht_361 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_362 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h16a == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_362 <= _pht_T_3;
        end else begin
          pht_362 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_363 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h16b == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_363 <= _pht_T_3;
        end else begin
          pht_363 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_364 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h16c == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_364 <= _pht_T_3;
        end else begin
          pht_364 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_365 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h16d == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_365 <= _pht_T_3;
        end else begin
          pht_365 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_366 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h16e == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_366 <= _pht_T_3;
        end else begin
          pht_366 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_367 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h16f == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_367 <= _pht_T_3;
        end else begin
          pht_367 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_368 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h170 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_368 <= _pht_T_3;
        end else begin
          pht_368 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_369 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h171 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_369 <= _pht_T_3;
        end else begin
          pht_369 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_370 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h172 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_370 <= _pht_T_3;
        end else begin
          pht_370 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_371 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h173 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_371 <= _pht_T_3;
        end else begin
          pht_371 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_372 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h174 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_372 <= _pht_T_3;
        end else begin
          pht_372 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_373 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h175 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_373 <= _pht_T_3;
        end else begin
          pht_373 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_374 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h176 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_374 <= _pht_T_3;
        end else begin
          pht_374 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_375 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h177 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_375 <= _pht_T_3;
        end else begin
          pht_375 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_376 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h178 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_376 <= _pht_T_3;
        end else begin
          pht_376 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_377 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h179 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_377 <= _pht_T_3;
        end else begin
          pht_377 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_378 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h17a == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_378 <= _pht_T_3;
        end else begin
          pht_378 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_379 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h17b == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_379 <= _pht_T_3;
        end else begin
          pht_379 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_380 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h17c == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_380 <= _pht_T_3;
        end else begin
          pht_380 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_381 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h17d == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_381 <= _pht_T_3;
        end else begin
          pht_381 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_382 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h17e == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_382 <= _pht_T_3;
        end else begin
          pht_382 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_383 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h17f == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_383 <= _pht_T_3;
        end else begin
          pht_383 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_384 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h180 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_384 <= _pht_T_3;
        end else begin
          pht_384 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_385 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h181 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_385 <= _pht_T_3;
        end else begin
          pht_385 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_386 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h182 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_386 <= _pht_T_3;
        end else begin
          pht_386 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_387 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h183 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_387 <= _pht_T_3;
        end else begin
          pht_387 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_388 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h184 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_388 <= _pht_T_3;
        end else begin
          pht_388 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_389 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h185 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_389 <= _pht_T_3;
        end else begin
          pht_389 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_390 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h186 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_390 <= _pht_T_3;
        end else begin
          pht_390 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_391 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h187 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_391 <= _pht_T_3;
        end else begin
          pht_391 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_392 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h188 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_392 <= _pht_T_3;
        end else begin
          pht_392 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_393 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h189 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_393 <= _pht_T_3;
        end else begin
          pht_393 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_394 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h18a == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_394 <= _pht_T_3;
        end else begin
          pht_394 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_395 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h18b == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_395 <= _pht_T_3;
        end else begin
          pht_395 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_396 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h18c == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_396 <= _pht_T_3;
        end else begin
          pht_396 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_397 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h18d == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_397 <= _pht_T_3;
        end else begin
          pht_397 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_398 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h18e == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_398 <= _pht_T_3;
        end else begin
          pht_398 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_399 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h18f == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_399 <= _pht_T_3;
        end else begin
          pht_399 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_400 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h190 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_400 <= _pht_T_3;
        end else begin
          pht_400 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_401 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h191 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_401 <= _pht_T_3;
        end else begin
          pht_401 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_402 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h192 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_402 <= _pht_T_3;
        end else begin
          pht_402 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_403 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h193 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_403 <= _pht_T_3;
        end else begin
          pht_403 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_404 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h194 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_404 <= _pht_T_3;
        end else begin
          pht_404 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_405 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h195 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_405 <= _pht_T_3;
        end else begin
          pht_405 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_406 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h196 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_406 <= _pht_T_3;
        end else begin
          pht_406 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_407 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h197 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_407 <= _pht_T_3;
        end else begin
          pht_407 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_408 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h198 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_408 <= _pht_T_3;
        end else begin
          pht_408 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_409 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h199 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_409 <= _pht_T_3;
        end else begin
          pht_409 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_410 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h19a == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_410 <= _pht_T_3;
        end else begin
          pht_410 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_411 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h19b == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_411 <= _pht_T_3;
        end else begin
          pht_411 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_412 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h19c == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_412 <= _pht_T_3;
        end else begin
          pht_412 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_413 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h19d == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_413 <= _pht_T_3;
        end else begin
          pht_413 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_414 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h19e == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_414 <= _pht_T_3;
        end else begin
          pht_414 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_415 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h19f == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_415 <= _pht_T_3;
        end else begin
          pht_415 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_416 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1a0 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_416 <= _pht_T_3;
        end else begin
          pht_416 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_417 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1a1 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_417 <= _pht_T_3;
        end else begin
          pht_417 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_418 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1a2 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_418 <= _pht_T_3;
        end else begin
          pht_418 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_419 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1a3 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_419 <= _pht_T_3;
        end else begin
          pht_419 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_420 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1a4 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_420 <= _pht_T_3;
        end else begin
          pht_420 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_421 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1a5 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_421 <= _pht_T_3;
        end else begin
          pht_421 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_422 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1a6 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_422 <= _pht_T_3;
        end else begin
          pht_422 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_423 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1a7 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_423 <= _pht_T_3;
        end else begin
          pht_423 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_424 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1a8 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_424 <= _pht_T_3;
        end else begin
          pht_424 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_425 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1a9 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_425 <= _pht_T_3;
        end else begin
          pht_425 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_426 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1aa == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_426 <= _pht_T_3;
        end else begin
          pht_426 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_427 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1ab == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_427 <= _pht_T_3;
        end else begin
          pht_427 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_428 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1ac == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_428 <= _pht_T_3;
        end else begin
          pht_428 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_429 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1ad == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_429 <= _pht_T_3;
        end else begin
          pht_429 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_430 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1ae == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_430 <= _pht_T_3;
        end else begin
          pht_430 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_431 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1af == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_431 <= _pht_T_3;
        end else begin
          pht_431 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_432 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1b0 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_432 <= _pht_T_3;
        end else begin
          pht_432 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_433 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1b1 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_433 <= _pht_T_3;
        end else begin
          pht_433 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_434 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1b2 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_434 <= _pht_T_3;
        end else begin
          pht_434 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_435 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1b3 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_435 <= _pht_T_3;
        end else begin
          pht_435 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_436 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1b4 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_436 <= _pht_T_3;
        end else begin
          pht_436 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_437 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1b5 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_437 <= _pht_T_3;
        end else begin
          pht_437 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_438 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1b6 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_438 <= _pht_T_3;
        end else begin
          pht_438 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_439 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1b7 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_439 <= _pht_T_3;
        end else begin
          pht_439 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_440 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1b8 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_440 <= _pht_T_3;
        end else begin
          pht_440 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_441 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1b9 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_441 <= _pht_T_3;
        end else begin
          pht_441 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_442 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1ba == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_442 <= _pht_T_3;
        end else begin
          pht_442 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_443 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1bb == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_443 <= _pht_T_3;
        end else begin
          pht_443 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_444 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1bc == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_444 <= _pht_T_3;
        end else begin
          pht_444 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_445 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1bd == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_445 <= _pht_T_3;
        end else begin
          pht_445 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_446 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1be == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_446 <= _pht_T_3;
        end else begin
          pht_446 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_447 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1bf == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_447 <= _pht_T_3;
        end else begin
          pht_447 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_448 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1c0 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_448 <= _pht_T_3;
        end else begin
          pht_448 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_449 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1c1 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_449 <= _pht_T_3;
        end else begin
          pht_449 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_450 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1c2 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_450 <= _pht_T_3;
        end else begin
          pht_450 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_451 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1c3 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_451 <= _pht_T_3;
        end else begin
          pht_451 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_452 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1c4 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_452 <= _pht_T_3;
        end else begin
          pht_452 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_453 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1c5 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_453 <= _pht_T_3;
        end else begin
          pht_453 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_454 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1c6 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_454 <= _pht_T_3;
        end else begin
          pht_454 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_455 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1c7 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_455 <= _pht_T_3;
        end else begin
          pht_455 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_456 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1c8 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_456 <= _pht_T_3;
        end else begin
          pht_456 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_457 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1c9 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_457 <= _pht_T_3;
        end else begin
          pht_457 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_458 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1ca == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_458 <= _pht_T_3;
        end else begin
          pht_458 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_459 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1cb == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_459 <= _pht_T_3;
        end else begin
          pht_459 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_460 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1cc == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_460 <= _pht_T_3;
        end else begin
          pht_460 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_461 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1cd == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_461 <= _pht_T_3;
        end else begin
          pht_461 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_462 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1ce == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_462 <= _pht_T_3;
        end else begin
          pht_462 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_463 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1cf == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_463 <= _pht_T_3;
        end else begin
          pht_463 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_464 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1d0 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_464 <= _pht_T_3;
        end else begin
          pht_464 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_465 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1d1 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_465 <= _pht_T_3;
        end else begin
          pht_465 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_466 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1d2 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_466 <= _pht_T_3;
        end else begin
          pht_466 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_467 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1d3 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_467 <= _pht_T_3;
        end else begin
          pht_467 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_468 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1d4 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_468 <= _pht_T_3;
        end else begin
          pht_468 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_469 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1d5 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_469 <= _pht_T_3;
        end else begin
          pht_469 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_470 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1d6 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_470 <= _pht_T_3;
        end else begin
          pht_470 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_471 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1d7 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_471 <= _pht_T_3;
        end else begin
          pht_471 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_472 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1d8 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_472 <= _pht_T_3;
        end else begin
          pht_472 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_473 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1d9 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_473 <= _pht_T_3;
        end else begin
          pht_473 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_474 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1da == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_474 <= _pht_T_3;
        end else begin
          pht_474 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_475 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1db == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_475 <= _pht_T_3;
        end else begin
          pht_475 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_476 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1dc == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_476 <= _pht_T_3;
        end else begin
          pht_476 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_477 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1dd == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_477 <= _pht_T_3;
        end else begin
          pht_477 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_478 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1de == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_478 <= _pht_T_3;
        end else begin
          pht_478 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_479 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1df == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_479 <= _pht_T_3;
        end else begin
          pht_479 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_480 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1e0 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_480 <= _pht_T_3;
        end else begin
          pht_480 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_481 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1e1 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_481 <= _pht_T_3;
        end else begin
          pht_481 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_482 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1e2 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_482 <= _pht_T_3;
        end else begin
          pht_482 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_483 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1e3 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_483 <= _pht_T_3;
        end else begin
          pht_483 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_484 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1e4 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_484 <= _pht_T_3;
        end else begin
          pht_484 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_485 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1e5 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_485 <= _pht_T_3;
        end else begin
          pht_485 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_486 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1e6 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_486 <= _pht_T_3;
        end else begin
          pht_486 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_487 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1e7 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_487 <= _pht_T_3;
        end else begin
          pht_487 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_488 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1e8 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_488 <= _pht_T_3;
        end else begin
          pht_488 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_489 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1e9 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_489 <= _pht_T_3;
        end else begin
          pht_489 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_490 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1ea == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_490 <= _pht_T_3;
        end else begin
          pht_490 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_491 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1eb == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_491 <= _pht_T_3;
        end else begin
          pht_491 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_492 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1ec == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_492 <= _pht_T_3;
        end else begin
          pht_492 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_493 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1ed == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_493 <= _pht_T_3;
        end else begin
          pht_493 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_494 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1ee == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_494 <= _pht_T_3;
        end else begin
          pht_494 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_495 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1ef == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_495 <= _pht_T_3;
        end else begin
          pht_495 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_496 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1f0 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_496 <= _pht_T_3;
        end else begin
          pht_496 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_497 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1f1 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_497 <= _pht_T_3;
        end else begin
          pht_497 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_498 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1f2 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_498 <= _pht_T_3;
        end else begin
          pht_498 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_499 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1f3 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_499 <= _pht_T_3;
        end else begin
          pht_499 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_500 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1f4 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_500 <= _pht_T_3;
        end else begin
          pht_500 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_501 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1f5 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_501 <= _pht_T_3;
        end else begin
          pht_501 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_502 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1f6 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_502 <= _pht_T_3;
        end else begin
          pht_502 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_503 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1f7 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_503 <= _pht_T_3;
        end else begin
          pht_503 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_504 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1f8 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_504 <= _pht_T_3;
        end else begin
          pht_504 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_505 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1f9 == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_505 <= _pht_T_3;
        end else begin
          pht_505 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_506 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1fa == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_506 <= _pht_T_3;
        end else begin
          pht_506 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_507 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1fb == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_507 <= _pht_T_3;
        end else begin
          pht_507 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_508 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1fc == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_508 <= _pht_T_3;
        end else begin
          pht_508 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_509 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1fd == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_509 <= _pht_T_3;
        end else begin
          pht_509 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_510 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1fe == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_510 <= _pht_T_3;
        end else begin
          pht_510 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 27:20]
      pht_511 <= 2'h1; // @[BPU.scala 27:20]
    end else if (io_jmp_packet_bp_update) begin // @[BPU.scala 53:33]
      if (9'h1ff == pht_widx) begin // @[BPU.scala 55:19]
        if (2'h3 == _GEN_1056) begin // @[Mux.scala 81:58]
          pht_511 <= _pht_T_3;
        end else begin
          pht_511 <= _pht_T_7;
        end
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_0_tag <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'h0 == btb_replace_idx) begin // @[BPU.scala 80:33]
        btb_0_tag <= io_jmp_packet_bp_pc[38:2]; // @[BPU.scala 80:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_0_target <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'h0 == btb_replace_idx) begin // @[BPU.scala 81:33]
        btb_0_target <= io_jmp_packet_target[38:2]; // @[BPU.scala 81:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_0_valid <= 1'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      btb_0_valid <= _GEN_2114;
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_1_tag <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'h1 == btb_replace_idx) begin // @[BPU.scala 80:33]
        btb_1_tag <= io_jmp_packet_bp_pc[38:2]; // @[BPU.scala 80:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_1_target <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'h1 == btb_replace_idx) begin // @[BPU.scala 81:33]
        btb_1_target <= io_jmp_packet_target[38:2]; // @[BPU.scala 81:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_1_valid <= 1'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      btb_1_valid <= _GEN_2115;
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_2_tag <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'h2 == btb_replace_idx) begin // @[BPU.scala 80:33]
        btb_2_tag <= io_jmp_packet_bp_pc[38:2]; // @[BPU.scala 80:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_2_target <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'h2 == btb_replace_idx) begin // @[BPU.scala 81:33]
        btb_2_target <= io_jmp_packet_target[38:2]; // @[BPU.scala 81:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_2_valid <= 1'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      btb_2_valid <= _GEN_2116;
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_3_tag <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'h3 == btb_replace_idx) begin // @[BPU.scala 80:33]
        btb_3_tag <= io_jmp_packet_bp_pc[38:2]; // @[BPU.scala 80:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_3_target <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'h3 == btb_replace_idx) begin // @[BPU.scala 81:33]
        btb_3_target <= io_jmp_packet_target[38:2]; // @[BPU.scala 81:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_3_valid <= 1'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      btb_3_valid <= _GEN_2117;
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_4_tag <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'h4 == btb_replace_idx) begin // @[BPU.scala 80:33]
        btb_4_tag <= io_jmp_packet_bp_pc[38:2]; // @[BPU.scala 80:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_4_target <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'h4 == btb_replace_idx) begin // @[BPU.scala 81:33]
        btb_4_target <= io_jmp_packet_target[38:2]; // @[BPU.scala 81:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_4_valid <= 1'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      btb_4_valid <= _GEN_2118;
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_5_tag <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'h5 == btb_replace_idx) begin // @[BPU.scala 80:33]
        btb_5_tag <= io_jmp_packet_bp_pc[38:2]; // @[BPU.scala 80:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_5_target <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'h5 == btb_replace_idx) begin // @[BPU.scala 81:33]
        btb_5_target <= io_jmp_packet_target[38:2]; // @[BPU.scala 81:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_5_valid <= 1'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      btb_5_valid <= _GEN_2119;
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_6_tag <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'h6 == btb_replace_idx) begin // @[BPU.scala 80:33]
        btb_6_tag <= io_jmp_packet_bp_pc[38:2]; // @[BPU.scala 80:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_6_target <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'h6 == btb_replace_idx) begin // @[BPU.scala 81:33]
        btb_6_target <= io_jmp_packet_target[38:2]; // @[BPU.scala 81:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_6_valid <= 1'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      btb_6_valid <= _GEN_2120;
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_7_tag <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'h7 == btb_replace_idx) begin // @[BPU.scala 80:33]
        btb_7_tag <= io_jmp_packet_bp_pc[38:2]; // @[BPU.scala 80:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_7_target <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'h7 == btb_replace_idx) begin // @[BPU.scala 81:33]
        btb_7_target <= io_jmp_packet_target[38:2]; // @[BPU.scala 81:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_7_valid <= 1'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      btb_7_valid <= _GEN_2121;
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_8_tag <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'h8 == btb_replace_idx) begin // @[BPU.scala 80:33]
        btb_8_tag <= io_jmp_packet_bp_pc[38:2]; // @[BPU.scala 80:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_8_target <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'h8 == btb_replace_idx) begin // @[BPU.scala 81:33]
        btb_8_target <= io_jmp_packet_target[38:2]; // @[BPU.scala 81:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_8_valid <= 1'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      btb_8_valid <= _GEN_2122;
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_9_tag <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'h9 == btb_replace_idx) begin // @[BPU.scala 80:33]
        btb_9_tag <= io_jmp_packet_bp_pc[38:2]; // @[BPU.scala 80:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_9_target <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'h9 == btb_replace_idx) begin // @[BPU.scala 81:33]
        btb_9_target <= io_jmp_packet_target[38:2]; // @[BPU.scala 81:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_9_valid <= 1'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      btb_9_valid <= _GEN_2123;
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_10_tag <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'ha == btb_replace_idx) begin // @[BPU.scala 80:33]
        btb_10_tag <= io_jmp_packet_bp_pc[38:2]; // @[BPU.scala 80:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_10_target <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'ha == btb_replace_idx) begin // @[BPU.scala 81:33]
        btb_10_target <= io_jmp_packet_target[38:2]; // @[BPU.scala 81:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_10_valid <= 1'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      btb_10_valid <= _GEN_2124;
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_11_tag <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'hb == btb_replace_idx) begin // @[BPU.scala 80:33]
        btb_11_tag <= io_jmp_packet_bp_pc[38:2]; // @[BPU.scala 80:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_11_target <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'hb == btb_replace_idx) begin // @[BPU.scala 81:33]
        btb_11_target <= io_jmp_packet_target[38:2]; // @[BPU.scala 81:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_11_valid <= 1'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      btb_11_valid <= _GEN_2125;
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_12_tag <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'hc == btb_replace_idx) begin // @[BPU.scala 80:33]
        btb_12_tag <= io_jmp_packet_bp_pc[38:2]; // @[BPU.scala 80:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_12_target <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'hc == btb_replace_idx) begin // @[BPU.scala 81:33]
        btb_12_target <= io_jmp_packet_target[38:2]; // @[BPU.scala 81:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_12_valid <= 1'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      btb_12_valid <= _GEN_2126;
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_13_tag <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'hd == btb_replace_idx) begin // @[BPU.scala 80:33]
        btb_13_tag <= io_jmp_packet_bp_pc[38:2]; // @[BPU.scala 80:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_13_target <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'hd == btb_replace_idx) begin // @[BPU.scala 81:33]
        btb_13_target <= io_jmp_packet_target[38:2]; // @[BPU.scala 81:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_13_valid <= 1'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      btb_13_valid <= _GEN_2127;
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_14_tag <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'he == btb_replace_idx) begin // @[BPU.scala 80:33]
        btb_14_tag <= io_jmp_packet_bp_pc[38:2]; // @[BPU.scala 80:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_14_target <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'he == btb_replace_idx) begin // @[BPU.scala 81:33]
        btb_14_target <= io_jmp_packet_target[38:2]; // @[BPU.scala 81:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_14_valid <= 1'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      btb_14_valid <= _GEN_2128;
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_15_tag <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'hf == btb_replace_idx) begin // @[BPU.scala 80:33]
        btb_15_tag <= io_jmp_packet_bp_pc[38:2]; // @[BPU.scala 80:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_15_target <= 37'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      if (4'hf == btb_replace_idx) begin // @[BPU.scala 81:33]
        btb_15_target <= io_jmp_packet_target[38:2]; // @[BPU.scala 81:33]
      end
    end
    if (reset) begin // @[BPU.scala 28:20]
      btb_15_valid <= 1'h0; // @[BPU.scala 28:20]
    end else if (io_jmp_packet_bp_update & io_jmp_packet_bp_taken) begin // @[BPU.scala 78:59]
      btb_15_valid <= _GEN_2129;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ghr = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  pht_0 = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  pht_1 = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  pht_2 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  pht_3 = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  pht_4 = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  pht_5 = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  pht_6 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  pht_7 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  pht_8 = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  pht_9 = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  pht_10 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  pht_11 = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  pht_12 = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  pht_13 = _RAND_14[1:0];
  _RAND_15 = {1{`RANDOM}};
  pht_14 = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  pht_15 = _RAND_16[1:0];
  _RAND_17 = {1{`RANDOM}};
  pht_16 = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  pht_17 = _RAND_18[1:0];
  _RAND_19 = {1{`RANDOM}};
  pht_18 = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  pht_19 = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  pht_20 = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  pht_21 = _RAND_22[1:0];
  _RAND_23 = {1{`RANDOM}};
  pht_22 = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  pht_23 = _RAND_24[1:0];
  _RAND_25 = {1{`RANDOM}};
  pht_24 = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  pht_25 = _RAND_26[1:0];
  _RAND_27 = {1{`RANDOM}};
  pht_26 = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  pht_27 = _RAND_28[1:0];
  _RAND_29 = {1{`RANDOM}};
  pht_28 = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  pht_29 = _RAND_30[1:0];
  _RAND_31 = {1{`RANDOM}};
  pht_30 = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  pht_31 = _RAND_32[1:0];
  _RAND_33 = {1{`RANDOM}};
  pht_32 = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  pht_33 = _RAND_34[1:0];
  _RAND_35 = {1{`RANDOM}};
  pht_34 = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  pht_35 = _RAND_36[1:0];
  _RAND_37 = {1{`RANDOM}};
  pht_36 = _RAND_37[1:0];
  _RAND_38 = {1{`RANDOM}};
  pht_37 = _RAND_38[1:0];
  _RAND_39 = {1{`RANDOM}};
  pht_38 = _RAND_39[1:0];
  _RAND_40 = {1{`RANDOM}};
  pht_39 = _RAND_40[1:0];
  _RAND_41 = {1{`RANDOM}};
  pht_40 = _RAND_41[1:0];
  _RAND_42 = {1{`RANDOM}};
  pht_41 = _RAND_42[1:0];
  _RAND_43 = {1{`RANDOM}};
  pht_42 = _RAND_43[1:0];
  _RAND_44 = {1{`RANDOM}};
  pht_43 = _RAND_44[1:0];
  _RAND_45 = {1{`RANDOM}};
  pht_44 = _RAND_45[1:0];
  _RAND_46 = {1{`RANDOM}};
  pht_45 = _RAND_46[1:0];
  _RAND_47 = {1{`RANDOM}};
  pht_46 = _RAND_47[1:0];
  _RAND_48 = {1{`RANDOM}};
  pht_47 = _RAND_48[1:0];
  _RAND_49 = {1{`RANDOM}};
  pht_48 = _RAND_49[1:0];
  _RAND_50 = {1{`RANDOM}};
  pht_49 = _RAND_50[1:0];
  _RAND_51 = {1{`RANDOM}};
  pht_50 = _RAND_51[1:0];
  _RAND_52 = {1{`RANDOM}};
  pht_51 = _RAND_52[1:0];
  _RAND_53 = {1{`RANDOM}};
  pht_52 = _RAND_53[1:0];
  _RAND_54 = {1{`RANDOM}};
  pht_53 = _RAND_54[1:0];
  _RAND_55 = {1{`RANDOM}};
  pht_54 = _RAND_55[1:0];
  _RAND_56 = {1{`RANDOM}};
  pht_55 = _RAND_56[1:0];
  _RAND_57 = {1{`RANDOM}};
  pht_56 = _RAND_57[1:0];
  _RAND_58 = {1{`RANDOM}};
  pht_57 = _RAND_58[1:0];
  _RAND_59 = {1{`RANDOM}};
  pht_58 = _RAND_59[1:0];
  _RAND_60 = {1{`RANDOM}};
  pht_59 = _RAND_60[1:0];
  _RAND_61 = {1{`RANDOM}};
  pht_60 = _RAND_61[1:0];
  _RAND_62 = {1{`RANDOM}};
  pht_61 = _RAND_62[1:0];
  _RAND_63 = {1{`RANDOM}};
  pht_62 = _RAND_63[1:0];
  _RAND_64 = {1{`RANDOM}};
  pht_63 = _RAND_64[1:0];
  _RAND_65 = {1{`RANDOM}};
  pht_64 = _RAND_65[1:0];
  _RAND_66 = {1{`RANDOM}};
  pht_65 = _RAND_66[1:0];
  _RAND_67 = {1{`RANDOM}};
  pht_66 = _RAND_67[1:0];
  _RAND_68 = {1{`RANDOM}};
  pht_67 = _RAND_68[1:0];
  _RAND_69 = {1{`RANDOM}};
  pht_68 = _RAND_69[1:0];
  _RAND_70 = {1{`RANDOM}};
  pht_69 = _RAND_70[1:0];
  _RAND_71 = {1{`RANDOM}};
  pht_70 = _RAND_71[1:0];
  _RAND_72 = {1{`RANDOM}};
  pht_71 = _RAND_72[1:0];
  _RAND_73 = {1{`RANDOM}};
  pht_72 = _RAND_73[1:0];
  _RAND_74 = {1{`RANDOM}};
  pht_73 = _RAND_74[1:0];
  _RAND_75 = {1{`RANDOM}};
  pht_74 = _RAND_75[1:0];
  _RAND_76 = {1{`RANDOM}};
  pht_75 = _RAND_76[1:0];
  _RAND_77 = {1{`RANDOM}};
  pht_76 = _RAND_77[1:0];
  _RAND_78 = {1{`RANDOM}};
  pht_77 = _RAND_78[1:0];
  _RAND_79 = {1{`RANDOM}};
  pht_78 = _RAND_79[1:0];
  _RAND_80 = {1{`RANDOM}};
  pht_79 = _RAND_80[1:0];
  _RAND_81 = {1{`RANDOM}};
  pht_80 = _RAND_81[1:0];
  _RAND_82 = {1{`RANDOM}};
  pht_81 = _RAND_82[1:0];
  _RAND_83 = {1{`RANDOM}};
  pht_82 = _RAND_83[1:0];
  _RAND_84 = {1{`RANDOM}};
  pht_83 = _RAND_84[1:0];
  _RAND_85 = {1{`RANDOM}};
  pht_84 = _RAND_85[1:0];
  _RAND_86 = {1{`RANDOM}};
  pht_85 = _RAND_86[1:0];
  _RAND_87 = {1{`RANDOM}};
  pht_86 = _RAND_87[1:0];
  _RAND_88 = {1{`RANDOM}};
  pht_87 = _RAND_88[1:0];
  _RAND_89 = {1{`RANDOM}};
  pht_88 = _RAND_89[1:0];
  _RAND_90 = {1{`RANDOM}};
  pht_89 = _RAND_90[1:0];
  _RAND_91 = {1{`RANDOM}};
  pht_90 = _RAND_91[1:0];
  _RAND_92 = {1{`RANDOM}};
  pht_91 = _RAND_92[1:0];
  _RAND_93 = {1{`RANDOM}};
  pht_92 = _RAND_93[1:0];
  _RAND_94 = {1{`RANDOM}};
  pht_93 = _RAND_94[1:0];
  _RAND_95 = {1{`RANDOM}};
  pht_94 = _RAND_95[1:0];
  _RAND_96 = {1{`RANDOM}};
  pht_95 = _RAND_96[1:0];
  _RAND_97 = {1{`RANDOM}};
  pht_96 = _RAND_97[1:0];
  _RAND_98 = {1{`RANDOM}};
  pht_97 = _RAND_98[1:0];
  _RAND_99 = {1{`RANDOM}};
  pht_98 = _RAND_99[1:0];
  _RAND_100 = {1{`RANDOM}};
  pht_99 = _RAND_100[1:0];
  _RAND_101 = {1{`RANDOM}};
  pht_100 = _RAND_101[1:0];
  _RAND_102 = {1{`RANDOM}};
  pht_101 = _RAND_102[1:0];
  _RAND_103 = {1{`RANDOM}};
  pht_102 = _RAND_103[1:0];
  _RAND_104 = {1{`RANDOM}};
  pht_103 = _RAND_104[1:0];
  _RAND_105 = {1{`RANDOM}};
  pht_104 = _RAND_105[1:0];
  _RAND_106 = {1{`RANDOM}};
  pht_105 = _RAND_106[1:0];
  _RAND_107 = {1{`RANDOM}};
  pht_106 = _RAND_107[1:0];
  _RAND_108 = {1{`RANDOM}};
  pht_107 = _RAND_108[1:0];
  _RAND_109 = {1{`RANDOM}};
  pht_108 = _RAND_109[1:0];
  _RAND_110 = {1{`RANDOM}};
  pht_109 = _RAND_110[1:0];
  _RAND_111 = {1{`RANDOM}};
  pht_110 = _RAND_111[1:0];
  _RAND_112 = {1{`RANDOM}};
  pht_111 = _RAND_112[1:0];
  _RAND_113 = {1{`RANDOM}};
  pht_112 = _RAND_113[1:0];
  _RAND_114 = {1{`RANDOM}};
  pht_113 = _RAND_114[1:0];
  _RAND_115 = {1{`RANDOM}};
  pht_114 = _RAND_115[1:0];
  _RAND_116 = {1{`RANDOM}};
  pht_115 = _RAND_116[1:0];
  _RAND_117 = {1{`RANDOM}};
  pht_116 = _RAND_117[1:0];
  _RAND_118 = {1{`RANDOM}};
  pht_117 = _RAND_118[1:0];
  _RAND_119 = {1{`RANDOM}};
  pht_118 = _RAND_119[1:0];
  _RAND_120 = {1{`RANDOM}};
  pht_119 = _RAND_120[1:0];
  _RAND_121 = {1{`RANDOM}};
  pht_120 = _RAND_121[1:0];
  _RAND_122 = {1{`RANDOM}};
  pht_121 = _RAND_122[1:0];
  _RAND_123 = {1{`RANDOM}};
  pht_122 = _RAND_123[1:0];
  _RAND_124 = {1{`RANDOM}};
  pht_123 = _RAND_124[1:0];
  _RAND_125 = {1{`RANDOM}};
  pht_124 = _RAND_125[1:0];
  _RAND_126 = {1{`RANDOM}};
  pht_125 = _RAND_126[1:0];
  _RAND_127 = {1{`RANDOM}};
  pht_126 = _RAND_127[1:0];
  _RAND_128 = {1{`RANDOM}};
  pht_127 = _RAND_128[1:0];
  _RAND_129 = {1{`RANDOM}};
  pht_128 = _RAND_129[1:0];
  _RAND_130 = {1{`RANDOM}};
  pht_129 = _RAND_130[1:0];
  _RAND_131 = {1{`RANDOM}};
  pht_130 = _RAND_131[1:0];
  _RAND_132 = {1{`RANDOM}};
  pht_131 = _RAND_132[1:0];
  _RAND_133 = {1{`RANDOM}};
  pht_132 = _RAND_133[1:0];
  _RAND_134 = {1{`RANDOM}};
  pht_133 = _RAND_134[1:0];
  _RAND_135 = {1{`RANDOM}};
  pht_134 = _RAND_135[1:0];
  _RAND_136 = {1{`RANDOM}};
  pht_135 = _RAND_136[1:0];
  _RAND_137 = {1{`RANDOM}};
  pht_136 = _RAND_137[1:0];
  _RAND_138 = {1{`RANDOM}};
  pht_137 = _RAND_138[1:0];
  _RAND_139 = {1{`RANDOM}};
  pht_138 = _RAND_139[1:0];
  _RAND_140 = {1{`RANDOM}};
  pht_139 = _RAND_140[1:0];
  _RAND_141 = {1{`RANDOM}};
  pht_140 = _RAND_141[1:0];
  _RAND_142 = {1{`RANDOM}};
  pht_141 = _RAND_142[1:0];
  _RAND_143 = {1{`RANDOM}};
  pht_142 = _RAND_143[1:0];
  _RAND_144 = {1{`RANDOM}};
  pht_143 = _RAND_144[1:0];
  _RAND_145 = {1{`RANDOM}};
  pht_144 = _RAND_145[1:0];
  _RAND_146 = {1{`RANDOM}};
  pht_145 = _RAND_146[1:0];
  _RAND_147 = {1{`RANDOM}};
  pht_146 = _RAND_147[1:0];
  _RAND_148 = {1{`RANDOM}};
  pht_147 = _RAND_148[1:0];
  _RAND_149 = {1{`RANDOM}};
  pht_148 = _RAND_149[1:0];
  _RAND_150 = {1{`RANDOM}};
  pht_149 = _RAND_150[1:0];
  _RAND_151 = {1{`RANDOM}};
  pht_150 = _RAND_151[1:0];
  _RAND_152 = {1{`RANDOM}};
  pht_151 = _RAND_152[1:0];
  _RAND_153 = {1{`RANDOM}};
  pht_152 = _RAND_153[1:0];
  _RAND_154 = {1{`RANDOM}};
  pht_153 = _RAND_154[1:0];
  _RAND_155 = {1{`RANDOM}};
  pht_154 = _RAND_155[1:0];
  _RAND_156 = {1{`RANDOM}};
  pht_155 = _RAND_156[1:0];
  _RAND_157 = {1{`RANDOM}};
  pht_156 = _RAND_157[1:0];
  _RAND_158 = {1{`RANDOM}};
  pht_157 = _RAND_158[1:0];
  _RAND_159 = {1{`RANDOM}};
  pht_158 = _RAND_159[1:0];
  _RAND_160 = {1{`RANDOM}};
  pht_159 = _RAND_160[1:0];
  _RAND_161 = {1{`RANDOM}};
  pht_160 = _RAND_161[1:0];
  _RAND_162 = {1{`RANDOM}};
  pht_161 = _RAND_162[1:0];
  _RAND_163 = {1{`RANDOM}};
  pht_162 = _RAND_163[1:0];
  _RAND_164 = {1{`RANDOM}};
  pht_163 = _RAND_164[1:0];
  _RAND_165 = {1{`RANDOM}};
  pht_164 = _RAND_165[1:0];
  _RAND_166 = {1{`RANDOM}};
  pht_165 = _RAND_166[1:0];
  _RAND_167 = {1{`RANDOM}};
  pht_166 = _RAND_167[1:0];
  _RAND_168 = {1{`RANDOM}};
  pht_167 = _RAND_168[1:0];
  _RAND_169 = {1{`RANDOM}};
  pht_168 = _RAND_169[1:0];
  _RAND_170 = {1{`RANDOM}};
  pht_169 = _RAND_170[1:0];
  _RAND_171 = {1{`RANDOM}};
  pht_170 = _RAND_171[1:0];
  _RAND_172 = {1{`RANDOM}};
  pht_171 = _RAND_172[1:0];
  _RAND_173 = {1{`RANDOM}};
  pht_172 = _RAND_173[1:0];
  _RAND_174 = {1{`RANDOM}};
  pht_173 = _RAND_174[1:0];
  _RAND_175 = {1{`RANDOM}};
  pht_174 = _RAND_175[1:0];
  _RAND_176 = {1{`RANDOM}};
  pht_175 = _RAND_176[1:0];
  _RAND_177 = {1{`RANDOM}};
  pht_176 = _RAND_177[1:0];
  _RAND_178 = {1{`RANDOM}};
  pht_177 = _RAND_178[1:0];
  _RAND_179 = {1{`RANDOM}};
  pht_178 = _RAND_179[1:0];
  _RAND_180 = {1{`RANDOM}};
  pht_179 = _RAND_180[1:0];
  _RAND_181 = {1{`RANDOM}};
  pht_180 = _RAND_181[1:0];
  _RAND_182 = {1{`RANDOM}};
  pht_181 = _RAND_182[1:0];
  _RAND_183 = {1{`RANDOM}};
  pht_182 = _RAND_183[1:0];
  _RAND_184 = {1{`RANDOM}};
  pht_183 = _RAND_184[1:0];
  _RAND_185 = {1{`RANDOM}};
  pht_184 = _RAND_185[1:0];
  _RAND_186 = {1{`RANDOM}};
  pht_185 = _RAND_186[1:0];
  _RAND_187 = {1{`RANDOM}};
  pht_186 = _RAND_187[1:0];
  _RAND_188 = {1{`RANDOM}};
  pht_187 = _RAND_188[1:0];
  _RAND_189 = {1{`RANDOM}};
  pht_188 = _RAND_189[1:0];
  _RAND_190 = {1{`RANDOM}};
  pht_189 = _RAND_190[1:0];
  _RAND_191 = {1{`RANDOM}};
  pht_190 = _RAND_191[1:0];
  _RAND_192 = {1{`RANDOM}};
  pht_191 = _RAND_192[1:0];
  _RAND_193 = {1{`RANDOM}};
  pht_192 = _RAND_193[1:0];
  _RAND_194 = {1{`RANDOM}};
  pht_193 = _RAND_194[1:0];
  _RAND_195 = {1{`RANDOM}};
  pht_194 = _RAND_195[1:0];
  _RAND_196 = {1{`RANDOM}};
  pht_195 = _RAND_196[1:0];
  _RAND_197 = {1{`RANDOM}};
  pht_196 = _RAND_197[1:0];
  _RAND_198 = {1{`RANDOM}};
  pht_197 = _RAND_198[1:0];
  _RAND_199 = {1{`RANDOM}};
  pht_198 = _RAND_199[1:0];
  _RAND_200 = {1{`RANDOM}};
  pht_199 = _RAND_200[1:0];
  _RAND_201 = {1{`RANDOM}};
  pht_200 = _RAND_201[1:0];
  _RAND_202 = {1{`RANDOM}};
  pht_201 = _RAND_202[1:0];
  _RAND_203 = {1{`RANDOM}};
  pht_202 = _RAND_203[1:0];
  _RAND_204 = {1{`RANDOM}};
  pht_203 = _RAND_204[1:0];
  _RAND_205 = {1{`RANDOM}};
  pht_204 = _RAND_205[1:0];
  _RAND_206 = {1{`RANDOM}};
  pht_205 = _RAND_206[1:0];
  _RAND_207 = {1{`RANDOM}};
  pht_206 = _RAND_207[1:0];
  _RAND_208 = {1{`RANDOM}};
  pht_207 = _RAND_208[1:0];
  _RAND_209 = {1{`RANDOM}};
  pht_208 = _RAND_209[1:0];
  _RAND_210 = {1{`RANDOM}};
  pht_209 = _RAND_210[1:0];
  _RAND_211 = {1{`RANDOM}};
  pht_210 = _RAND_211[1:0];
  _RAND_212 = {1{`RANDOM}};
  pht_211 = _RAND_212[1:0];
  _RAND_213 = {1{`RANDOM}};
  pht_212 = _RAND_213[1:0];
  _RAND_214 = {1{`RANDOM}};
  pht_213 = _RAND_214[1:0];
  _RAND_215 = {1{`RANDOM}};
  pht_214 = _RAND_215[1:0];
  _RAND_216 = {1{`RANDOM}};
  pht_215 = _RAND_216[1:0];
  _RAND_217 = {1{`RANDOM}};
  pht_216 = _RAND_217[1:0];
  _RAND_218 = {1{`RANDOM}};
  pht_217 = _RAND_218[1:0];
  _RAND_219 = {1{`RANDOM}};
  pht_218 = _RAND_219[1:0];
  _RAND_220 = {1{`RANDOM}};
  pht_219 = _RAND_220[1:0];
  _RAND_221 = {1{`RANDOM}};
  pht_220 = _RAND_221[1:0];
  _RAND_222 = {1{`RANDOM}};
  pht_221 = _RAND_222[1:0];
  _RAND_223 = {1{`RANDOM}};
  pht_222 = _RAND_223[1:0];
  _RAND_224 = {1{`RANDOM}};
  pht_223 = _RAND_224[1:0];
  _RAND_225 = {1{`RANDOM}};
  pht_224 = _RAND_225[1:0];
  _RAND_226 = {1{`RANDOM}};
  pht_225 = _RAND_226[1:0];
  _RAND_227 = {1{`RANDOM}};
  pht_226 = _RAND_227[1:0];
  _RAND_228 = {1{`RANDOM}};
  pht_227 = _RAND_228[1:0];
  _RAND_229 = {1{`RANDOM}};
  pht_228 = _RAND_229[1:0];
  _RAND_230 = {1{`RANDOM}};
  pht_229 = _RAND_230[1:0];
  _RAND_231 = {1{`RANDOM}};
  pht_230 = _RAND_231[1:0];
  _RAND_232 = {1{`RANDOM}};
  pht_231 = _RAND_232[1:0];
  _RAND_233 = {1{`RANDOM}};
  pht_232 = _RAND_233[1:0];
  _RAND_234 = {1{`RANDOM}};
  pht_233 = _RAND_234[1:0];
  _RAND_235 = {1{`RANDOM}};
  pht_234 = _RAND_235[1:0];
  _RAND_236 = {1{`RANDOM}};
  pht_235 = _RAND_236[1:0];
  _RAND_237 = {1{`RANDOM}};
  pht_236 = _RAND_237[1:0];
  _RAND_238 = {1{`RANDOM}};
  pht_237 = _RAND_238[1:0];
  _RAND_239 = {1{`RANDOM}};
  pht_238 = _RAND_239[1:0];
  _RAND_240 = {1{`RANDOM}};
  pht_239 = _RAND_240[1:0];
  _RAND_241 = {1{`RANDOM}};
  pht_240 = _RAND_241[1:0];
  _RAND_242 = {1{`RANDOM}};
  pht_241 = _RAND_242[1:0];
  _RAND_243 = {1{`RANDOM}};
  pht_242 = _RAND_243[1:0];
  _RAND_244 = {1{`RANDOM}};
  pht_243 = _RAND_244[1:0];
  _RAND_245 = {1{`RANDOM}};
  pht_244 = _RAND_245[1:0];
  _RAND_246 = {1{`RANDOM}};
  pht_245 = _RAND_246[1:0];
  _RAND_247 = {1{`RANDOM}};
  pht_246 = _RAND_247[1:0];
  _RAND_248 = {1{`RANDOM}};
  pht_247 = _RAND_248[1:0];
  _RAND_249 = {1{`RANDOM}};
  pht_248 = _RAND_249[1:0];
  _RAND_250 = {1{`RANDOM}};
  pht_249 = _RAND_250[1:0];
  _RAND_251 = {1{`RANDOM}};
  pht_250 = _RAND_251[1:0];
  _RAND_252 = {1{`RANDOM}};
  pht_251 = _RAND_252[1:0];
  _RAND_253 = {1{`RANDOM}};
  pht_252 = _RAND_253[1:0];
  _RAND_254 = {1{`RANDOM}};
  pht_253 = _RAND_254[1:0];
  _RAND_255 = {1{`RANDOM}};
  pht_254 = _RAND_255[1:0];
  _RAND_256 = {1{`RANDOM}};
  pht_255 = _RAND_256[1:0];
  _RAND_257 = {1{`RANDOM}};
  pht_256 = _RAND_257[1:0];
  _RAND_258 = {1{`RANDOM}};
  pht_257 = _RAND_258[1:0];
  _RAND_259 = {1{`RANDOM}};
  pht_258 = _RAND_259[1:0];
  _RAND_260 = {1{`RANDOM}};
  pht_259 = _RAND_260[1:0];
  _RAND_261 = {1{`RANDOM}};
  pht_260 = _RAND_261[1:0];
  _RAND_262 = {1{`RANDOM}};
  pht_261 = _RAND_262[1:0];
  _RAND_263 = {1{`RANDOM}};
  pht_262 = _RAND_263[1:0];
  _RAND_264 = {1{`RANDOM}};
  pht_263 = _RAND_264[1:0];
  _RAND_265 = {1{`RANDOM}};
  pht_264 = _RAND_265[1:0];
  _RAND_266 = {1{`RANDOM}};
  pht_265 = _RAND_266[1:0];
  _RAND_267 = {1{`RANDOM}};
  pht_266 = _RAND_267[1:0];
  _RAND_268 = {1{`RANDOM}};
  pht_267 = _RAND_268[1:0];
  _RAND_269 = {1{`RANDOM}};
  pht_268 = _RAND_269[1:0];
  _RAND_270 = {1{`RANDOM}};
  pht_269 = _RAND_270[1:0];
  _RAND_271 = {1{`RANDOM}};
  pht_270 = _RAND_271[1:0];
  _RAND_272 = {1{`RANDOM}};
  pht_271 = _RAND_272[1:0];
  _RAND_273 = {1{`RANDOM}};
  pht_272 = _RAND_273[1:0];
  _RAND_274 = {1{`RANDOM}};
  pht_273 = _RAND_274[1:0];
  _RAND_275 = {1{`RANDOM}};
  pht_274 = _RAND_275[1:0];
  _RAND_276 = {1{`RANDOM}};
  pht_275 = _RAND_276[1:0];
  _RAND_277 = {1{`RANDOM}};
  pht_276 = _RAND_277[1:0];
  _RAND_278 = {1{`RANDOM}};
  pht_277 = _RAND_278[1:0];
  _RAND_279 = {1{`RANDOM}};
  pht_278 = _RAND_279[1:0];
  _RAND_280 = {1{`RANDOM}};
  pht_279 = _RAND_280[1:0];
  _RAND_281 = {1{`RANDOM}};
  pht_280 = _RAND_281[1:0];
  _RAND_282 = {1{`RANDOM}};
  pht_281 = _RAND_282[1:0];
  _RAND_283 = {1{`RANDOM}};
  pht_282 = _RAND_283[1:0];
  _RAND_284 = {1{`RANDOM}};
  pht_283 = _RAND_284[1:0];
  _RAND_285 = {1{`RANDOM}};
  pht_284 = _RAND_285[1:0];
  _RAND_286 = {1{`RANDOM}};
  pht_285 = _RAND_286[1:0];
  _RAND_287 = {1{`RANDOM}};
  pht_286 = _RAND_287[1:0];
  _RAND_288 = {1{`RANDOM}};
  pht_287 = _RAND_288[1:0];
  _RAND_289 = {1{`RANDOM}};
  pht_288 = _RAND_289[1:0];
  _RAND_290 = {1{`RANDOM}};
  pht_289 = _RAND_290[1:0];
  _RAND_291 = {1{`RANDOM}};
  pht_290 = _RAND_291[1:0];
  _RAND_292 = {1{`RANDOM}};
  pht_291 = _RAND_292[1:0];
  _RAND_293 = {1{`RANDOM}};
  pht_292 = _RAND_293[1:0];
  _RAND_294 = {1{`RANDOM}};
  pht_293 = _RAND_294[1:0];
  _RAND_295 = {1{`RANDOM}};
  pht_294 = _RAND_295[1:0];
  _RAND_296 = {1{`RANDOM}};
  pht_295 = _RAND_296[1:0];
  _RAND_297 = {1{`RANDOM}};
  pht_296 = _RAND_297[1:0];
  _RAND_298 = {1{`RANDOM}};
  pht_297 = _RAND_298[1:0];
  _RAND_299 = {1{`RANDOM}};
  pht_298 = _RAND_299[1:0];
  _RAND_300 = {1{`RANDOM}};
  pht_299 = _RAND_300[1:0];
  _RAND_301 = {1{`RANDOM}};
  pht_300 = _RAND_301[1:0];
  _RAND_302 = {1{`RANDOM}};
  pht_301 = _RAND_302[1:0];
  _RAND_303 = {1{`RANDOM}};
  pht_302 = _RAND_303[1:0];
  _RAND_304 = {1{`RANDOM}};
  pht_303 = _RAND_304[1:0];
  _RAND_305 = {1{`RANDOM}};
  pht_304 = _RAND_305[1:0];
  _RAND_306 = {1{`RANDOM}};
  pht_305 = _RAND_306[1:0];
  _RAND_307 = {1{`RANDOM}};
  pht_306 = _RAND_307[1:0];
  _RAND_308 = {1{`RANDOM}};
  pht_307 = _RAND_308[1:0];
  _RAND_309 = {1{`RANDOM}};
  pht_308 = _RAND_309[1:0];
  _RAND_310 = {1{`RANDOM}};
  pht_309 = _RAND_310[1:0];
  _RAND_311 = {1{`RANDOM}};
  pht_310 = _RAND_311[1:0];
  _RAND_312 = {1{`RANDOM}};
  pht_311 = _RAND_312[1:0];
  _RAND_313 = {1{`RANDOM}};
  pht_312 = _RAND_313[1:0];
  _RAND_314 = {1{`RANDOM}};
  pht_313 = _RAND_314[1:0];
  _RAND_315 = {1{`RANDOM}};
  pht_314 = _RAND_315[1:0];
  _RAND_316 = {1{`RANDOM}};
  pht_315 = _RAND_316[1:0];
  _RAND_317 = {1{`RANDOM}};
  pht_316 = _RAND_317[1:0];
  _RAND_318 = {1{`RANDOM}};
  pht_317 = _RAND_318[1:0];
  _RAND_319 = {1{`RANDOM}};
  pht_318 = _RAND_319[1:0];
  _RAND_320 = {1{`RANDOM}};
  pht_319 = _RAND_320[1:0];
  _RAND_321 = {1{`RANDOM}};
  pht_320 = _RAND_321[1:0];
  _RAND_322 = {1{`RANDOM}};
  pht_321 = _RAND_322[1:0];
  _RAND_323 = {1{`RANDOM}};
  pht_322 = _RAND_323[1:0];
  _RAND_324 = {1{`RANDOM}};
  pht_323 = _RAND_324[1:0];
  _RAND_325 = {1{`RANDOM}};
  pht_324 = _RAND_325[1:0];
  _RAND_326 = {1{`RANDOM}};
  pht_325 = _RAND_326[1:0];
  _RAND_327 = {1{`RANDOM}};
  pht_326 = _RAND_327[1:0];
  _RAND_328 = {1{`RANDOM}};
  pht_327 = _RAND_328[1:0];
  _RAND_329 = {1{`RANDOM}};
  pht_328 = _RAND_329[1:0];
  _RAND_330 = {1{`RANDOM}};
  pht_329 = _RAND_330[1:0];
  _RAND_331 = {1{`RANDOM}};
  pht_330 = _RAND_331[1:0];
  _RAND_332 = {1{`RANDOM}};
  pht_331 = _RAND_332[1:0];
  _RAND_333 = {1{`RANDOM}};
  pht_332 = _RAND_333[1:0];
  _RAND_334 = {1{`RANDOM}};
  pht_333 = _RAND_334[1:0];
  _RAND_335 = {1{`RANDOM}};
  pht_334 = _RAND_335[1:0];
  _RAND_336 = {1{`RANDOM}};
  pht_335 = _RAND_336[1:0];
  _RAND_337 = {1{`RANDOM}};
  pht_336 = _RAND_337[1:0];
  _RAND_338 = {1{`RANDOM}};
  pht_337 = _RAND_338[1:0];
  _RAND_339 = {1{`RANDOM}};
  pht_338 = _RAND_339[1:0];
  _RAND_340 = {1{`RANDOM}};
  pht_339 = _RAND_340[1:0];
  _RAND_341 = {1{`RANDOM}};
  pht_340 = _RAND_341[1:0];
  _RAND_342 = {1{`RANDOM}};
  pht_341 = _RAND_342[1:0];
  _RAND_343 = {1{`RANDOM}};
  pht_342 = _RAND_343[1:0];
  _RAND_344 = {1{`RANDOM}};
  pht_343 = _RAND_344[1:0];
  _RAND_345 = {1{`RANDOM}};
  pht_344 = _RAND_345[1:0];
  _RAND_346 = {1{`RANDOM}};
  pht_345 = _RAND_346[1:0];
  _RAND_347 = {1{`RANDOM}};
  pht_346 = _RAND_347[1:0];
  _RAND_348 = {1{`RANDOM}};
  pht_347 = _RAND_348[1:0];
  _RAND_349 = {1{`RANDOM}};
  pht_348 = _RAND_349[1:0];
  _RAND_350 = {1{`RANDOM}};
  pht_349 = _RAND_350[1:0];
  _RAND_351 = {1{`RANDOM}};
  pht_350 = _RAND_351[1:0];
  _RAND_352 = {1{`RANDOM}};
  pht_351 = _RAND_352[1:0];
  _RAND_353 = {1{`RANDOM}};
  pht_352 = _RAND_353[1:0];
  _RAND_354 = {1{`RANDOM}};
  pht_353 = _RAND_354[1:0];
  _RAND_355 = {1{`RANDOM}};
  pht_354 = _RAND_355[1:0];
  _RAND_356 = {1{`RANDOM}};
  pht_355 = _RAND_356[1:0];
  _RAND_357 = {1{`RANDOM}};
  pht_356 = _RAND_357[1:0];
  _RAND_358 = {1{`RANDOM}};
  pht_357 = _RAND_358[1:0];
  _RAND_359 = {1{`RANDOM}};
  pht_358 = _RAND_359[1:0];
  _RAND_360 = {1{`RANDOM}};
  pht_359 = _RAND_360[1:0];
  _RAND_361 = {1{`RANDOM}};
  pht_360 = _RAND_361[1:0];
  _RAND_362 = {1{`RANDOM}};
  pht_361 = _RAND_362[1:0];
  _RAND_363 = {1{`RANDOM}};
  pht_362 = _RAND_363[1:0];
  _RAND_364 = {1{`RANDOM}};
  pht_363 = _RAND_364[1:0];
  _RAND_365 = {1{`RANDOM}};
  pht_364 = _RAND_365[1:0];
  _RAND_366 = {1{`RANDOM}};
  pht_365 = _RAND_366[1:0];
  _RAND_367 = {1{`RANDOM}};
  pht_366 = _RAND_367[1:0];
  _RAND_368 = {1{`RANDOM}};
  pht_367 = _RAND_368[1:0];
  _RAND_369 = {1{`RANDOM}};
  pht_368 = _RAND_369[1:0];
  _RAND_370 = {1{`RANDOM}};
  pht_369 = _RAND_370[1:0];
  _RAND_371 = {1{`RANDOM}};
  pht_370 = _RAND_371[1:0];
  _RAND_372 = {1{`RANDOM}};
  pht_371 = _RAND_372[1:0];
  _RAND_373 = {1{`RANDOM}};
  pht_372 = _RAND_373[1:0];
  _RAND_374 = {1{`RANDOM}};
  pht_373 = _RAND_374[1:0];
  _RAND_375 = {1{`RANDOM}};
  pht_374 = _RAND_375[1:0];
  _RAND_376 = {1{`RANDOM}};
  pht_375 = _RAND_376[1:0];
  _RAND_377 = {1{`RANDOM}};
  pht_376 = _RAND_377[1:0];
  _RAND_378 = {1{`RANDOM}};
  pht_377 = _RAND_378[1:0];
  _RAND_379 = {1{`RANDOM}};
  pht_378 = _RAND_379[1:0];
  _RAND_380 = {1{`RANDOM}};
  pht_379 = _RAND_380[1:0];
  _RAND_381 = {1{`RANDOM}};
  pht_380 = _RAND_381[1:0];
  _RAND_382 = {1{`RANDOM}};
  pht_381 = _RAND_382[1:0];
  _RAND_383 = {1{`RANDOM}};
  pht_382 = _RAND_383[1:0];
  _RAND_384 = {1{`RANDOM}};
  pht_383 = _RAND_384[1:0];
  _RAND_385 = {1{`RANDOM}};
  pht_384 = _RAND_385[1:0];
  _RAND_386 = {1{`RANDOM}};
  pht_385 = _RAND_386[1:0];
  _RAND_387 = {1{`RANDOM}};
  pht_386 = _RAND_387[1:0];
  _RAND_388 = {1{`RANDOM}};
  pht_387 = _RAND_388[1:0];
  _RAND_389 = {1{`RANDOM}};
  pht_388 = _RAND_389[1:0];
  _RAND_390 = {1{`RANDOM}};
  pht_389 = _RAND_390[1:0];
  _RAND_391 = {1{`RANDOM}};
  pht_390 = _RAND_391[1:0];
  _RAND_392 = {1{`RANDOM}};
  pht_391 = _RAND_392[1:0];
  _RAND_393 = {1{`RANDOM}};
  pht_392 = _RAND_393[1:0];
  _RAND_394 = {1{`RANDOM}};
  pht_393 = _RAND_394[1:0];
  _RAND_395 = {1{`RANDOM}};
  pht_394 = _RAND_395[1:0];
  _RAND_396 = {1{`RANDOM}};
  pht_395 = _RAND_396[1:0];
  _RAND_397 = {1{`RANDOM}};
  pht_396 = _RAND_397[1:0];
  _RAND_398 = {1{`RANDOM}};
  pht_397 = _RAND_398[1:0];
  _RAND_399 = {1{`RANDOM}};
  pht_398 = _RAND_399[1:0];
  _RAND_400 = {1{`RANDOM}};
  pht_399 = _RAND_400[1:0];
  _RAND_401 = {1{`RANDOM}};
  pht_400 = _RAND_401[1:0];
  _RAND_402 = {1{`RANDOM}};
  pht_401 = _RAND_402[1:0];
  _RAND_403 = {1{`RANDOM}};
  pht_402 = _RAND_403[1:0];
  _RAND_404 = {1{`RANDOM}};
  pht_403 = _RAND_404[1:0];
  _RAND_405 = {1{`RANDOM}};
  pht_404 = _RAND_405[1:0];
  _RAND_406 = {1{`RANDOM}};
  pht_405 = _RAND_406[1:0];
  _RAND_407 = {1{`RANDOM}};
  pht_406 = _RAND_407[1:0];
  _RAND_408 = {1{`RANDOM}};
  pht_407 = _RAND_408[1:0];
  _RAND_409 = {1{`RANDOM}};
  pht_408 = _RAND_409[1:0];
  _RAND_410 = {1{`RANDOM}};
  pht_409 = _RAND_410[1:0];
  _RAND_411 = {1{`RANDOM}};
  pht_410 = _RAND_411[1:0];
  _RAND_412 = {1{`RANDOM}};
  pht_411 = _RAND_412[1:0];
  _RAND_413 = {1{`RANDOM}};
  pht_412 = _RAND_413[1:0];
  _RAND_414 = {1{`RANDOM}};
  pht_413 = _RAND_414[1:0];
  _RAND_415 = {1{`RANDOM}};
  pht_414 = _RAND_415[1:0];
  _RAND_416 = {1{`RANDOM}};
  pht_415 = _RAND_416[1:0];
  _RAND_417 = {1{`RANDOM}};
  pht_416 = _RAND_417[1:0];
  _RAND_418 = {1{`RANDOM}};
  pht_417 = _RAND_418[1:0];
  _RAND_419 = {1{`RANDOM}};
  pht_418 = _RAND_419[1:0];
  _RAND_420 = {1{`RANDOM}};
  pht_419 = _RAND_420[1:0];
  _RAND_421 = {1{`RANDOM}};
  pht_420 = _RAND_421[1:0];
  _RAND_422 = {1{`RANDOM}};
  pht_421 = _RAND_422[1:0];
  _RAND_423 = {1{`RANDOM}};
  pht_422 = _RAND_423[1:0];
  _RAND_424 = {1{`RANDOM}};
  pht_423 = _RAND_424[1:0];
  _RAND_425 = {1{`RANDOM}};
  pht_424 = _RAND_425[1:0];
  _RAND_426 = {1{`RANDOM}};
  pht_425 = _RAND_426[1:0];
  _RAND_427 = {1{`RANDOM}};
  pht_426 = _RAND_427[1:0];
  _RAND_428 = {1{`RANDOM}};
  pht_427 = _RAND_428[1:0];
  _RAND_429 = {1{`RANDOM}};
  pht_428 = _RAND_429[1:0];
  _RAND_430 = {1{`RANDOM}};
  pht_429 = _RAND_430[1:0];
  _RAND_431 = {1{`RANDOM}};
  pht_430 = _RAND_431[1:0];
  _RAND_432 = {1{`RANDOM}};
  pht_431 = _RAND_432[1:0];
  _RAND_433 = {1{`RANDOM}};
  pht_432 = _RAND_433[1:0];
  _RAND_434 = {1{`RANDOM}};
  pht_433 = _RAND_434[1:0];
  _RAND_435 = {1{`RANDOM}};
  pht_434 = _RAND_435[1:0];
  _RAND_436 = {1{`RANDOM}};
  pht_435 = _RAND_436[1:0];
  _RAND_437 = {1{`RANDOM}};
  pht_436 = _RAND_437[1:0];
  _RAND_438 = {1{`RANDOM}};
  pht_437 = _RAND_438[1:0];
  _RAND_439 = {1{`RANDOM}};
  pht_438 = _RAND_439[1:0];
  _RAND_440 = {1{`RANDOM}};
  pht_439 = _RAND_440[1:0];
  _RAND_441 = {1{`RANDOM}};
  pht_440 = _RAND_441[1:0];
  _RAND_442 = {1{`RANDOM}};
  pht_441 = _RAND_442[1:0];
  _RAND_443 = {1{`RANDOM}};
  pht_442 = _RAND_443[1:0];
  _RAND_444 = {1{`RANDOM}};
  pht_443 = _RAND_444[1:0];
  _RAND_445 = {1{`RANDOM}};
  pht_444 = _RAND_445[1:0];
  _RAND_446 = {1{`RANDOM}};
  pht_445 = _RAND_446[1:0];
  _RAND_447 = {1{`RANDOM}};
  pht_446 = _RAND_447[1:0];
  _RAND_448 = {1{`RANDOM}};
  pht_447 = _RAND_448[1:0];
  _RAND_449 = {1{`RANDOM}};
  pht_448 = _RAND_449[1:0];
  _RAND_450 = {1{`RANDOM}};
  pht_449 = _RAND_450[1:0];
  _RAND_451 = {1{`RANDOM}};
  pht_450 = _RAND_451[1:0];
  _RAND_452 = {1{`RANDOM}};
  pht_451 = _RAND_452[1:0];
  _RAND_453 = {1{`RANDOM}};
  pht_452 = _RAND_453[1:0];
  _RAND_454 = {1{`RANDOM}};
  pht_453 = _RAND_454[1:0];
  _RAND_455 = {1{`RANDOM}};
  pht_454 = _RAND_455[1:0];
  _RAND_456 = {1{`RANDOM}};
  pht_455 = _RAND_456[1:0];
  _RAND_457 = {1{`RANDOM}};
  pht_456 = _RAND_457[1:0];
  _RAND_458 = {1{`RANDOM}};
  pht_457 = _RAND_458[1:0];
  _RAND_459 = {1{`RANDOM}};
  pht_458 = _RAND_459[1:0];
  _RAND_460 = {1{`RANDOM}};
  pht_459 = _RAND_460[1:0];
  _RAND_461 = {1{`RANDOM}};
  pht_460 = _RAND_461[1:0];
  _RAND_462 = {1{`RANDOM}};
  pht_461 = _RAND_462[1:0];
  _RAND_463 = {1{`RANDOM}};
  pht_462 = _RAND_463[1:0];
  _RAND_464 = {1{`RANDOM}};
  pht_463 = _RAND_464[1:0];
  _RAND_465 = {1{`RANDOM}};
  pht_464 = _RAND_465[1:0];
  _RAND_466 = {1{`RANDOM}};
  pht_465 = _RAND_466[1:0];
  _RAND_467 = {1{`RANDOM}};
  pht_466 = _RAND_467[1:0];
  _RAND_468 = {1{`RANDOM}};
  pht_467 = _RAND_468[1:0];
  _RAND_469 = {1{`RANDOM}};
  pht_468 = _RAND_469[1:0];
  _RAND_470 = {1{`RANDOM}};
  pht_469 = _RAND_470[1:0];
  _RAND_471 = {1{`RANDOM}};
  pht_470 = _RAND_471[1:0];
  _RAND_472 = {1{`RANDOM}};
  pht_471 = _RAND_472[1:0];
  _RAND_473 = {1{`RANDOM}};
  pht_472 = _RAND_473[1:0];
  _RAND_474 = {1{`RANDOM}};
  pht_473 = _RAND_474[1:0];
  _RAND_475 = {1{`RANDOM}};
  pht_474 = _RAND_475[1:0];
  _RAND_476 = {1{`RANDOM}};
  pht_475 = _RAND_476[1:0];
  _RAND_477 = {1{`RANDOM}};
  pht_476 = _RAND_477[1:0];
  _RAND_478 = {1{`RANDOM}};
  pht_477 = _RAND_478[1:0];
  _RAND_479 = {1{`RANDOM}};
  pht_478 = _RAND_479[1:0];
  _RAND_480 = {1{`RANDOM}};
  pht_479 = _RAND_480[1:0];
  _RAND_481 = {1{`RANDOM}};
  pht_480 = _RAND_481[1:0];
  _RAND_482 = {1{`RANDOM}};
  pht_481 = _RAND_482[1:0];
  _RAND_483 = {1{`RANDOM}};
  pht_482 = _RAND_483[1:0];
  _RAND_484 = {1{`RANDOM}};
  pht_483 = _RAND_484[1:0];
  _RAND_485 = {1{`RANDOM}};
  pht_484 = _RAND_485[1:0];
  _RAND_486 = {1{`RANDOM}};
  pht_485 = _RAND_486[1:0];
  _RAND_487 = {1{`RANDOM}};
  pht_486 = _RAND_487[1:0];
  _RAND_488 = {1{`RANDOM}};
  pht_487 = _RAND_488[1:0];
  _RAND_489 = {1{`RANDOM}};
  pht_488 = _RAND_489[1:0];
  _RAND_490 = {1{`RANDOM}};
  pht_489 = _RAND_490[1:0];
  _RAND_491 = {1{`RANDOM}};
  pht_490 = _RAND_491[1:0];
  _RAND_492 = {1{`RANDOM}};
  pht_491 = _RAND_492[1:0];
  _RAND_493 = {1{`RANDOM}};
  pht_492 = _RAND_493[1:0];
  _RAND_494 = {1{`RANDOM}};
  pht_493 = _RAND_494[1:0];
  _RAND_495 = {1{`RANDOM}};
  pht_494 = _RAND_495[1:0];
  _RAND_496 = {1{`RANDOM}};
  pht_495 = _RAND_496[1:0];
  _RAND_497 = {1{`RANDOM}};
  pht_496 = _RAND_497[1:0];
  _RAND_498 = {1{`RANDOM}};
  pht_497 = _RAND_498[1:0];
  _RAND_499 = {1{`RANDOM}};
  pht_498 = _RAND_499[1:0];
  _RAND_500 = {1{`RANDOM}};
  pht_499 = _RAND_500[1:0];
  _RAND_501 = {1{`RANDOM}};
  pht_500 = _RAND_501[1:0];
  _RAND_502 = {1{`RANDOM}};
  pht_501 = _RAND_502[1:0];
  _RAND_503 = {1{`RANDOM}};
  pht_502 = _RAND_503[1:0];
  _RAND_504 = {1{`RANDOM}};
  pht_503 = _RAND_504[1:0];
  _RAND_505 = {1{`RANDOM}};
  pht_504 = _RAND_505[1:0];
  _RAND_506 = {1{`RANDOM}};
  pht_505 = _RAND_506[1:0];
  _RAND_507 = {1{`RANDOM}};
  pht_506 = _RAND_507[1:0];
  _RAND_508 = {1{`RANDOM}};
  pht_507 = _RAND_508[1:0];
  _RAND_509 = {1{`RANDOM}};
  pht_508 = _RAND_509[1:0];
  _RAND_510 = {1{`RANDOM}};
  pht_509 = _RAND_510[1:0];
  _RAND_511 = {1{`RANDOM}};
  pht_510 = _RAND_511[1:0];
  _RAND_512 = {1{`RANDOM}};
  pht_511 = _RAND_512[1:0];
  _RAND_513 = {2{`RANDOM}};
  btb_0_tag = _RAND_513[36:0];
  _RAND_514 = {2{`RANDOM}};
  btb_0_target = _RAND_514[36:0];
  _RAND_515 = {1{`RANDOM}};
  btb_0_valid = _RAND_515[0:0];
  _RAND_516 = {2{`RANDOM}};
  btb_1_tag = _RAND_516[36:0];
  _RAND_517 = {2{`RANDOM}};
  btb_1_target = _RAND_517[36:0];
  _RAND_518 = {1{`RANDOM}};
  btb_1_valid = _RAND_518[0:0];
  _RAND_519 = {2{`RANDOM}};
  btb_2_tag = _RAND_519[36:0];
  _RAND_520 = {2{`RANDOM}};
  btb_2_target = _RAND_520[36:0];
  _RAND_521 = {1{`RANDOM}};
  btb_2_valid = _RAND_521[0:0];
  _RAND_522 = {2{`RANDOM}};
  btb_3_tag = _RAND_522[36:0];
  _RAND_523 = {2{`RANDOM}};
  btb_3_target = _RAND_523[36:0];
  _RAND_524 = {1{`RANDOM}};
  btb_3_valid = _RAND_524[0:0];
  _RAND_525 = {2{`RANDOM}};
  btb_4_tag = _RAND_525[36:0];
  _RAND_526 = {2{`RANDOM}};
  btb_4_target = _RAND_526[36:0];
  _RAND_527 = {1{`RANDOM}};
  btb_4_valid = _RAND_527[0:0];
  _RAND_528 = {2{`RANDOM}};
  btb_5_tag = _RAND_528[36:0];
  _RAND_529 = {2{`RANDOM}};
  btb_5_target = _RAND_529[36:0];
  _RAND_530 = {1{`RANDOM}};
  btb_5_valid = _RAND_530[0:0];
  _RAND_531 = {2{`RANDOM}};
  btb_6_tag = _RAND_531[36:0];
  _RAND_532 = {2{`RANDOM}};
  btb_6_target = _RAND_532[36:0];
  _RAND_533 = {1{`RANDOM}};
  btb_6_valid = _RAND_533[0:0];
  _RAND_534 = {2{`RANDOM}};
  btb_7_tag = _RAND_534[36:0];
  _RAND_535 = {2{`RANDOM}};
  btb_7_target = _RAND_535[36:0];
  _RAND_536 = {1{`RANDOM}};
  btb_7_valid = _RAND_536[0:0];
  _RAND_537 = {2{`RANDOM}};
  btb_8_tag = _RAND_537[36:0];
  _RAND_538 = {2{`RANDOM}};
  btb_8_target = _RAND_538[36:0];
  _RAND_539 = {1{`RANDOM}};
  btb_8_valid = _RAND_539[0:0];
  _RAND_540 = {2{`RANDOM}};
  btb_9_tag = _RAND_540[36:0];
  _RAND_541 = {2{`RANDOM}};
  btb_9_target = _RAND_541[36:0];
  _RAND_542 = {1{`RANDOM}};
  btb_9_valid = _RAND_542[0:0];
  _RAND_543 = {2{`RANDOM}};
  btb_10_tag = _RAND_543[36:0];
  _RAND_544 = {2{`RANDOM}};
  btb_10_target = _RAND_544[36:0];
  _RAND_545 = {1{`RANDOM}};
  btb_10_valid = _RAND_545[0:0];
  _RAND_546 = {2{`RANDOM}};
  btb_11_tag = _RAND_546[36:0];
  _RAND_547 = {2{`RANDOM}};
  btb_11_target = _RAND_547[36:0];
  _RAND_548 = {1{`RANDOM}};
  btb_11_valid = _RAND_548[0:0];
  _RAND_549 = {2{`RANDOM}};
  btb_12_tag = _RAND_549[36:0];
  _RAND_550 = {2{`RANDOM}};
  btb_12_target = _RAND_550[36:0];
  _RAND_551 = {1{`RANDOM}};
  btb_12_valid = _RAND_551[0:0];
  _RAND_552 = {2{`RANDOM}};
  btb_13_tag = _RAND_552[36:0];
  _RAND_553 = {2{`RANDOM}};
  btb_13_target = _RAND_553[36:0];
  _RAND_554 = {1{`RANDOM}};
  btb_13_valid = _RAND_554[0:0];
  _RAND_555 = {2{`RANDOM}};
  btb_14_tag = _RAND_555[36:0];
  _RAND_556 = {2{`RANDOM}};
  btb_14_target = _RAND_556[36:0];
  _RAND_557 = {1{`RANDOM}};
  btb_14_valid = _RAND_557[0:0];
  _RAND_558 = {2{`RANDOM}};
  btb_15_tag = _RAND_558[36:0];
  _RAND_559 = {2{`RANDOM}};
  btb_15_target = _RAND_559[36:0];
  _RAND_560 = {1{`RANDOM}};
  btb_15_valid = _RAND_560[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IF0(
  input         clock,
  input         reset,
  input         io_jmp_packet_valid,
  input  [63:0] io_jmp_packet_target,
  input         io_jmp_packet_bp_update,
  input         io_jmp_packet_bp_taken,
  input  [63:0] io_jmp_packet_bp_pc,
  input         io_req_ready,
  output        io_req_valid,
  output [38:0] io_req_bits_addr,
  output [38:0] io_req_addr,
  output [63:0] io_bp_npc,
  input         io_stall_b
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  bpu_clock; // @[IFU.scala 21:21]
  wire  bpu_reset; // @[IFU.scala 21:21]
  wire [63:0] bpu_io_pc; // @[IFU.scala 21:21]
  wire [63:0] bpu_io_jmp_packet_target; // @[IFU.scala 21:21]
  wire  bpu_io_jmp_packet_bp_update; // @[IFU.scala 21:21]
  wire  bpu_io_jmp_packet_bp_taken; // @[IFU.scala 21:21]
  wire [63:0] bpu_io_jmp_packet_bp_pc; // @[IFU.scala 21:21]
  wire [63:0] bpu_io_out; // @[IFU.scala 21:21]
  wire  _pc_update_T = io_req_ready & io_req_valid; // @[Decoupled.scala 51:35]
  wire  pc_update = io_jmp_packet_valid | _pc_update_T; // @[IFU.scala 15:41]
  reg [63:0] pc; // @[Reg.scala 35:20]
  wire [63:0] jmp_target = {io_jmp_packet_target[63:2],2'h0}; // @[Cat.scala 33:92]
  wire [63:0] pc_next_raw = bpu_io_out; // @[IFU.scala 19:25 24:23]
  wire [63:0] _io_req_addr_T = io_jmp_packet_valid ? jmp_target : pc; // @[IFU.scala 33:26]
  BPU bpu ( // @[IFU.scala 21:21]
    .clock(bpu_clock),
    .reset(bpu_reset),
    .io_pc(bpu_io_pc),
    .io_jmp_packet_target(bpu_io_jmp_packet_target),
    .io_jmp_packet_bp_update(bpu_io_jmp_packet_bp_update),
    .io_jmp_packet_bp_taken(bpu_io_jmp_packet_bp_taken),
    .io_jmp_packet_bp_pc(bpu_io_jmp_packet_bp_pc),
    .io_out(bpu_io_out)
  );
  assign io_req_valid = io_stall_b; // @[IFU.scala 36:20]
  assign io_req_bits_addr = {io_req_addr[38:3],3'h0}; // @[Cat.scala 33:92]
  assign io_req_addr = _io_req_addr_T[38:0]; // @[IFU.scala 33:20]
  assign io_bp_npc = bpu_io_out; // @[IFU.scala 19:25 24:23]
  assign bpu_clock = clock;
  assign bpu_reset = reset;
  assign bpu_io_pc = io_jmp_packet_valid & _pc_update_T ? jmp_target : pc; // @[IFU.scala 22:29]
  assign bpu_io_jmp_packet_target = io_jmp_packet_target; // @[IFU.scala 23:23]
  assign bpu_io_jmp_packet_bp_update = io_jmp_packet_bp_update; // @[IFU.scala 23:23]
  assign bpu_io_jmp_packet_bp_taken = io_jmp_packet_bp_taken; // @[IFU.scala 23:23]
  assign bpu_io_jmp_packet_bp_pc = io_jmp_packet_bp_pc; // @[IFU.scala 23:23]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 35:20]
      pc <= 64'h10000; // @[Reg.scala 35:20]
    end else if (pc_update) begin // @[Reg.scala 36:18]
      if (io_jmp_packet_valid & ~_pc_update_T) begin // @[IFU.scala 31:20]
        pc <= jmp_target;
      end else begin
        pc <= pc_next_raw;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  pc = _RAND_0[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IF1(
  input   clock,
  input   reset,
  input   io_jmp_packet_valid,
  output  io_resp_ready,
  input   io_resp_valid,
  input   io_stall_b,
  output  io_out_valid,
  input   io_req_fire,
  input   io_pc_queue_empty
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[IFU.scala 51:50]
  wire  _jmp_r_T = io_resp_ready & io_resp_valid; // @[Decoupled.scala 51:35]
  wire  _jmp_r_T_6 = io_jmp_packet_valid & ~_jmp_r_T & state != 2'h2 & ~io_pc_queue_empty; // @[IFU.scala 54:64]
  reg  jmp_r; // @[Utils.scala 36:20]
  wire  _GEN_0 = _jmp_r_T_6 | jmp_r; // @[Utils.scala 41:19 36:20 41:23]
  wire  _state_to_wait_T_1 = ~jmp_r; // @[IFU.scala 58:81]
  wire  _state_to_wait_T_3 = ~io_jmp_packet_valid; // @[IFU.scala 58:91]
  wire [1:0] _state_T = io_jmp_packet_valid ? 2'h0 : 2'h1; // @[IFU.scala 68:21]
  wire [1:0] _GEN_4 = io_jmp_packet_valid ? 2'h0 : state; // @[IFU.scala 72:33 73:15 51:50]
  assign io_resp_ready = (io_stall_b | io_jmp_packet_valid) & state == 2'h1 | state == 2'h0; // @[IFU.scala 78:80]
  assign io_out_valid = _jmp_r_T & _state_to_wait_T_3 & _state_to_wait_T_1; // @[IFU.scala 81:56]
  always @(posedge clock) begin
    if (reset) begin // @[IFU.scala 51:50]
      state <= 2'h0; // @[IFU.scala 51:50]
    end else if (2'h0 == state) begin // @[IFU.scala 60:17]
      if (io_req_fire) begin // @[IFU.scala 62:25]
        state <= 2'h1; // @[IFU.scala 63:15]
      end
    end else if (2'h1 == state) begin // @[IFU.scala 60:17]
      if (_jmp_r_T) begin // @[IFU.scala 67:26]
        state <= _state_T; // @[IFU.scala 68:15]
      end
    end else if (2'h2 == state) begin // @[IFU.scala 60:17]
      state <= _GEN_4;
    end
    if (reset) begin // @[Utils.scala 36:20]
      jmp_r <= 1'h0; // @[Utils.scala 36:20]
    end else if (_jmp_r_T) begin // @[Utils.scala 42:18]
      jmp_r <= 1'h0; // @[Utils.scala 42:22]
    end else begin
      jmp_r <= _GEN_0;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  jmp_r = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [38:0] io_enq_bits,
  input         io_deq_ready,
  output        io_deq_valid,
  output [38:0] io_deq_bits,
  output        io_count
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [38:0] ram [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [38:0] ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [38:0] ram_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_MPORT_en; // @[Decoupled.scala 273:95]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 278:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  assign ram_io_deq_bits_MPORT_en = 1'h1;
  assign ram_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_MPORT_data = io_enq_bits;
  assign ram_MPORT_addr = 1'h0;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = io_deq_ready | empty; // @[Decoupled.scala 303:16 323:{24,39}]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits = ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_count = maybe_full; // @[Decoupled.scala 329:62]
  always @(posedge clock) begin
    if (ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram[initvar] = _RAND_0[38:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  maybe_full = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_1(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [63:0] io_enq_bits,
  input         io_deq_ready,
  output        io_deq_valid,
  output [63:0] io_deq_bits
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] ram [0:0]; // @[Decoupled.scala 273:95]
  wire  ram_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire  ram_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [63:0] ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [63:0] ram_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_MPORT_en; // @[Decoupled.scala 273:95]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 278:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  assign ram_io_deq_bits_MPORT_en = 1'h1;
  assign ram_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_MPORT_data = io_enq_bits;
  assign ram_MPORT_addr = 1'h0;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = io_deq_ready | empty; // @[Decoupled.scala 303:16 323:{24,39}]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits = ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  always @(posedge clock) begin
    if (ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram[initvar] = _RAND_0[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  maybe_full = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IFU(
  input         clock,
  input         reset,
  input         io_jmp_packet_valid,
  input  [63:0] io_jmp_packet_target,
  input         io_jmp_packet_bp_update,
  input         io_jmp_packet_bp_taken,
  input  [63:0] io_jmp_packet_bp_pc,
  input         io_imem_req_ready,
  output        io_imem_req_valid,
  output [38:0] io_imem_req_bits_addr,
  output        io_imem_resp_ready,
  input         io_imem_resp_valid,
  input  [63:0] io_imem_resp_bits_rdata,
  input         io_imem_resp_bits_page_fault,
  input         io_imem_resp_bits_access_fault,
  output [63:0] io_out_pc,
  output [31:0] io_out_instr,
  output        io_out_valid,
  output        io_out_page_fault,
  output        io_out_access_fault,
  output [63:0] io_out_bp_npc,
  input         io_stall_b
);
  wire  if0_clock; // @[IFU.scala 96:19]
  wire  if0_reset; // @[IFU.scala 96:19]
  wire  if0_io_jmp_packet_valid; // @[IFU.scala 96:19]
  wire [63:0] if0_io_jmp_packet_target; // @[IFU.scala 96:19]
  wire  if0_io_jmp_packet_bp_update; // @[IFU.scala 96:19]
  wire  if0_io_jmp_packet_bp_taken; // @[IFU.scala 96:19]
  wire [63:0] if0_io_jmp_packet_bp_pc; // @[IFU.scala 96:19]
  wire  if0_io_req_ready; // @[IFU.scala 96:19]
  wire  if0_io_req_valid; // @[IFU.scala 96:19]
  wire [38:0] if0_io_req_bits_addr; // @[IFU.scala 96:19]
  wire [38:0] if0_io_req_addr; // @[IFU.scala 96:19]
  wire [63:0] if0_io_bp_npc; // @[IFU.scala 96:19]
  wire  if0_io_stall_b; // @[IFU.scala 96:19]
  wire  if1_clock; // @[IFU.scala 97:19]
  wire  if1_reset; // @[IFU.scala 97:19]
  wire  if1_io_jmp_packet_valid; // @[IFU.scala 97:19]
  wire  if1_io_resp_ready; // @[IFU.scala 97:19]
  wire  if1_io_resp_valid; // @[IFU.scala 97:19]
  wire  if1_io_stall_b; // @[IFU.scala 97:19]
  wire  if1_io_out_valid; // @[IFU.scala 97:19]
  wire  if1_io_req_fire; // @[IFU.scala 97:19]
  wire  if1_io_pc_queue_empty; // @[IFU.scala 97:19]
  wire  pc_queue_clock; // @[IFU.scala 99:28]
  wire  pc_queue_reset; // @[IFU.scala 99:28]
  wire  pc_queue_io_enq_ready; // @[IFU.scala 99:28]
  wire  pc_queue_io_enq_valid; // @[IFU.scala 99:28]
  wire [38:0] pc_queue_io_enq_bits; // @[IFU.scala 99:28]
  wire  pc_queue_io_deq_ready; // @[IFU.scala 99:28]
  wire  pc_queue_io_deq_valid; // @[IFU.scala 99:28]
  wire [38:0] pc_queue_io_deq_bits; // @[IFU.scala 99:28]
  wire  pc_queue_io_count; // @[IFU.scala 99:28]
  wire  bp_npc_queue_clock; // @[IFU.scala 100:28]
  wire  bp_npc_queue_reset; // @[IFU.scala 100:28]
  wire  bp_npc_queue_io_enq_ready; // @[IFU.scala 100:28]
  wire  bp_npc_queue_io_enq_valid; // @[IFU.scala 100:28]
  wire [63:0] bp_npc_queue_io_enq_bits; // @[IFU.scala 100:28]
  wire  bp_npc_queue_io_deq_ready; // @[IFU.scala 100:28]
  wire  bp_npc_queue_io_deq_valid; // @[IFU.scala 100:28]
  wire [63:0] bp_npc_queue_io_deq_bits; // @[IFU.scala 100:28]
  wire [24:0] _io_out_pc_T_2 = pc_queue_io_deq_bits[38] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 77:12]
  IF0 if0 ( // @[IFU.scala 96:19]
    .clock(if0_clock),
    .reset(if0_reset),
    .io_jmp_packet_valid(if0_io_jmp_packet_valid),
    .io_jmp_packet_target(if0_io_jmp_packet_target),
    .io_jmp_packet_bp_update(if0_io_jmp_packet_bp_update),
    .io_jmp_packet_bp_taken(if0_io_jmp_packet_bp_taken),
    .io_jmp_packet_bp_pc(if0_io_jmp_packet_bp_pc),
    .io_req_ready(if0_io_req_ready),
    .io_req_valid(if0_io_req_valid),
    .io_req_bits_addr(if0_io_req_bits_addr),
    .io_req_addr(if0_io_req_addr),
    .io_bp_npc(if0_io_bp_npc),
    .io_stall_b(if0_io_stall_b)
  );
  IF1 if1 ( // @[IFU.scala 97:19]
    .clock(if1_clock),
    .reset(if1_reset),
    .io_jmp_packet_valid(if1_io_jmp_packet_valid),
    .io_resp_ready(if1_io_resp_ready),
    .io_resp_valid(if1_io_resp_valid),
    .io_stall_b(if1_io_stall_b),
    .io_out_valid(if1_io_out_valid),
    .io_req_fire(if1_io_req_fire),
    .io_pc_queue_empty(if1_io_pc_queue_empty)
  );
  Queue pc_queue ( // @[IFU.scala 99:28]
    .clock(pc_queue_clock),
    .reset(pc_queue_reset),
    .io_enq_ready(pc_queue_io_enq_ready),
    .io_enq_valid(pc_queue_io_enq_valid),
    .io_enq_bits(pc_queue_io_enq_bits),
    .io_deq_ready(pc_queue_io_deq_ready),
    .io_deq_valid(pc_queue_io_deq_valid),
    .io_deq_bits(pc_queue_io_deq_bits),
    .io_count(pc_queue_io_count)
  );
  Queue_1 bp_npc_queue ( // @[IFU.scala 100:28]
    .clock(bp_npc_queue_clock),
    .reset(bp_npc_queue_reset),
    .io_enq_ready(bp_npc_queue_io_enq_ready),
    .io_enq_valid(bp_npc_queue_io_enq_valid),
    .io_enq_bits(bp_npc_queue_io_enq_bits),
    .io_deq_ready(bp_npc_queue_io_deq_ready),
    .io_deq_valid(bp_npc_queue_io_deq_valid),
    .io_deq_bits(bp_npc_queue_io_deq_bits)
  );
  assign io_imem_req_valid = if0_io_req_valid; // @[IFU.scala 103:21]
  assign io_imem_req_bits_addr = if0_io_req_bits_addr; // @[IFU.scala 103:21]
  assign io_imem_resp_ready = if1_io_resp_ready; // @[IFU.scala 107:25]
  assign io_out_pc = {_io_out_pc_T_2,pc_queue_io_deq_bits}; // @[Cat.scala 33:92]
  assign io_out_instr = io_out_pc[2] ? io_imem_resp_bits_rdata[63:32] : io_imem_resp_bits_rdata[31:0]; // @[IFU.scala 122:29]
  assign io_out_valid = if1_io_out_valid; // @[IFU.scala 120:23]
  assign io_out_page_fault = io_imem_resp_bits_page_fault; // @[IFU.scala 123:23]
  assign io_out_access_fault = io_imem_resp_bits_access_fault; // @[IFU.scala 124:23]
  assign io_out_bp_npc = bp_npc_queue_io_deq_bits; // @[IFU.scala 125:23]
  assign if0_clock = clock;
  assign if0_reset = reset;
  assign if0_io_jmp_packet_valid = io_jmp_packet_valid; // @[IFU.scala 102:21]
  assign if0_io_jmp_packet_target = io_jmp_packet_target; // @[IFU.scala 102:21]
  assign if0_io_jmp_packet_bp_update = io_jmp_packet_bp_update; // @[IFU.scala 102:21]
  assign if0_io_jmp_packet_bp_taken = io_jmp_packet_bp_taken; // @[IFU.scala 102:21]
  assign if0_io_jmp_packet_bp_pc = io_jmp_packet_bp_pc; // @[IFU.scala 102:21]
  assign if0_io_req_ready = io_imem_req_ready; // @[IFU.scala 103:21]
  assign if0_io_stall_b = pc_queue_io_enq_ready & io_stall_b; // @[IFU.scala 104:46]
  assign if1_clock = clock;
  assign if1_reset = reset;
  assign if1_io_jmp_packet_valid = io_jmp_packet_valid; // @[IFU.scala 106:25]
  assign if1_io_resp_valid = io_imem_resp_valid; // @[IFU.scala 107:25]
  assign if1_io_stall_b = io_stall_b; // @[IFU.scala 108:25]
  assign if1_io_req_fire = io_imem_req_ready & io_imem_req_valid; // @[Decoupled.scala 51:35]
  assign if1_io_pc_queue_empty = ~pc_queue_io_count; // @[IFU.scala 110:47]
  assign pc_queue_clock = clock;
  assign pc_queue_reset = reset;
  assign pc_queue_io_enq_valid = io_imem_req_ready & io_imem_req_valid; // @[Decoupled.scala 51:35]
  assign pc_queue_io_enq_bits = if0_io_req_addr; // @[IFU.scala 112:25]
  assign pc_queue_io_deq_ready = io_imem_resp_ready & io_imem_resp_valid; // @[Decoupled.scala 51:35]
  assign bp_npc_queue_clock = clock;
  assign bp_npc_queue_reset = reset;
  assign bp_npc_queue_io_enq_valid = io_imem_req_ready & io_imem_req_valid; // @[Decoupled.scala 51:35]
  assign bp_npc_queue_io_enq_bits = if0_io_bp_npc; // @[IFU.scala 116:29]
  assign bp_npc_queue_io_deq_ready = io_imem_resp_ready & io_imem_resp_valid; // @[Decoupled.scala 51:35]
endmodule
module MaxPeriodFibonacciLFSR_1(
  input   clock,
  input   reset,
  output  io_out_0,
  output  io_out_1,
  output  io_out_2,
  output  io_out_3,
  output  io_out_4
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg  state_0; // @[PRNG.scala 55:49]
  reg  state_1; // @[PRNG.scala 55:49]
  reg  state_2; // @[PRNG.scala 55:49]
  reg  state_3; // @[PRNG.scala 55:49]
  reg  state_4; // @[PRNG.scala 55:49]
  wire  _T = state_4 ^ state_2; // @[LFSR.scala 15:41]
  assign io_out_0 = state_0; // @[PRNG.scala 78:10]
  assign io_out_1 = state_1; // @[PRNG.scala 78:10]
  assign io_out_2 = state_2; // @[PRNG.scala 78:10]
  assign io_out_3 = state_3; // @[PRNG.scala 78:10]
  assign io_out_4 = state_4; // @[PRNG.scala 78:10]
  always @(posedge clock) begin
    state_0 <= reset | _T; // @[PRNG.scala 55:{49,49}]
    if (reset) begin // @[PRNG.scala 55:49]
      state_1 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_1 <= state_0;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_2 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_2 <= state_1;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_3 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_3 <= state_2;
    end
    if (reset) begin // @[PRNG.scala 55:49]
      state_4 <= 1'h0; // @[PRNG.scala 55:49]
    end else begin
      state_4 <= state_3;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  state_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  state_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  state_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  state_4 = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLB(
  input         clock,
  input         reset,
  input         io_sfence_vma,
  input  [8:0]  io_vaddr_vpn2,
  input  [8:0]  io_vaddr_vpn1,
  input  [8:0]  io_vaddr_vpn0,
  output [1:0]  io_rpte_ppn2,
  output [8:0]  io_rpte_ppn1,
  output [8:0]  io_rpte_ppn0,
  output        io_rpte_flag_d,
  output        io_rpte_flag_a,
  output        io_rpte_flag_u,
  output        io_rpte_flag_x,
  output        io_rpte_flag_w,
  output        io_rpte_flag_r,
  output        io_rpte_flag_v,
  output [1:0]  io_rlevel,
  output        io_hit,
  input         io_wen,
  input  [8:0]  io_wvaddr_vpn2,
  input  [8:0]  io_wvaddr_vpn1,
  input  [8:0]  io_wvaddr_vpn0,
  input  [1:0]  io_wpte_ppn2,
  input  [8:0]  io_wpte_ppn1,
  input  [8:0]  io_wpte_ppn0,
  input         io_wpte_flag_d,
  input         io_wpte_flag_a,
  input         io_wpte_flag_g,
  input         io_wpte_flag_u,
  input         io_wpte_flag_x,
  input         io_wpte_flag_w,
  input         io_wpte_flag_r,
  input         io_wpte_flag_v,
  input  [1:0]  io_wlevel,
  input  [15:0] io_satp_asid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
`endif // RANDOMIZE_REG_INIT
  wire  replace_idx_prng_clock; // @[PRNG.scala 91:22]
  wire  replace_idx_prng_reset; // @[PRNG.scala 91:22]
  wire  replace_idx_prng_io_out_0; // @[PRNG.scala 91:22]
  wire  replace_idx_prng_io_out_1; // @[PRNG.scala 91:22]
  wire  replace_idx_prng_io_out_2; // @[PRNG.scala 91:22]
  wire  replace_idx_prng_io_out_3; // @[PRNG.scala 91:22]
  wire  replace_idx_prng_io_out_4; // @[PRNG.scala 91:22]
  wire  _T_2 = ~reset; // @[TLB.scala 48:9]
  wire [4:0] replace_idx = {replace_idx_prng_io_out_4,replace_idx_prng_io_out_3,replace_idx_prng_io_out_2,
    replace_idx_prng_io_out_1,replace_idx_prng_io_out_0}; // @[PRNG.scala 95:17]
  reg  array4kb_0_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_0_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_0_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_0_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_0_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_0_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_0_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_0_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_0_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_0_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_0_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_0_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_0_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_0_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_0_asid; // @[TLB.scala 64:31]
  reg  array4kb_1_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_1_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_1_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_1_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_1_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_1_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_1_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_1_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_1_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_1_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_1_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_1_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_1_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_1_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_1_asid; // @[TLB.scala 64:31]
  reg  array4kb_2_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_2_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_2_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_2_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_2_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_2_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_2_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_2_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_2_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_2_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_2_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_2_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_2_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_2_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_2_asid; // @[TLB.scala 64:31]
  reg  array4kb_3_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_3_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_3_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_3_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_3_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_3_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_3_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_3_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_3_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_3_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_3_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_3_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_3_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_3_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_3_asid; // @[TLB.scala 64:31]
  reg  array4kb_4_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_4_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_4_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_4_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_4_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_4_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_4_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_4_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_4_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_4_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_4_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_4_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_4_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_4_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_4_asid; // @[TLB.scala 64:31]
  reg  array4kb_5_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_5_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_5_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_5_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_5_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_5_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_5_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_5_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_5_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_5_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_5_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_5_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_5_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_5_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_5_asid; // @[TLB.scala 64:31]
  reg  array4kb_6_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_6_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_6_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_6_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_6_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_6_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_6_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_6_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_6_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_6_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_6_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_6_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_6_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_6_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_6_asid; // @[TLB.scala 64:31]
  reg  array4kb_7_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_7_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_7_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_7_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_7_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_7_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_7_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_7_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_7_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_7_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_7_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_7_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_7_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_7_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_7_asid; // @[TLB.scala 64:31]
  reg  array4kb_8_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_8_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_8_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_8_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_8_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_8_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_8_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_8_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_8_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_8_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_8_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_8_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_8_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_8_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_8_asid; // @[TLB.scala 64:31]
  reg  array4kb_9_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_9_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_9_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_9_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_9_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_9_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_9_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_9_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_9_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_9_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_9_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_9_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_9_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_9_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_9_asid; // @[TLB.scala 64:31]
  reg  array4kb_10_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_10_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_10_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_10_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_10_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_10_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_10_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_10_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_10_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_10_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_10_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_10_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_10_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_10_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_10_asid; // @[TLB.scala 64:31]
  reg  array4kb_11_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_11_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_11_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_11_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_11_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_11_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_11_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_11_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_11_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_11_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_11_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_11_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_11_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_11_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_11_asid; // @[TLB.scala 64:31]
  reg  array4kb_12_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_12_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_12_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_12_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_12_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_12_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_12_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_12_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_12_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_12_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_12_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_12_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_12_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_12_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_12_asid; // @[TLB.scala 64:31]
  reg  array4kb_13_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_13_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_13_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_13_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_13_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_13_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_13_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_13_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_13_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_13_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_13_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_13_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_13_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_13_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_13_asid; // @[TLB.scala 64:31]
  reg  array4kb_14_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_14_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_14_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_14_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_14_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_14_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_14_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_14_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_14_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_14_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_14_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_14_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_14_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_14_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_14_asid; // @[TLB.scala 64:31]
  reg  array4kb_15_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_15_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_15_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_15_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_15_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_15_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_15_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_15_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_15_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_15_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_15_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_15_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_15_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_15_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_15_asid; // @[TLB.scala 64:31]
  reg  array4kb_16_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_16_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_16_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_16_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_16_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_16_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_16_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_16_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_16_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_16_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_16_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_16_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_16_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_16_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_16_asid; // @[TLB.scala 64:31]
  reg  array4kb_17_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_17_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_17_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_17_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_17_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_17_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_17_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_17_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_17_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_17_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_17_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_17_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_17_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_17_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_17_asid; // @[TLB.scala 64:31]
  reg  array4kb_18_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_18_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_18_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_18_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_18_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_18_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_18_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_18_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_18_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_18_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_18_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_18_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_18_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_18_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_18_asid; // @[TLB.scala 64:31]
  reg  array4kb_19_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_19_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_19_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_19_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_19_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_19_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_19_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_19_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_19_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_19_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_19_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_19_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_19_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_19_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_19_asid; // @[TLB.scala 64:31]
  reg  array4kb_20_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_20_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_20_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_20_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_20_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_20_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_20_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_20_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_20_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_20_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_20_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_20_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_20_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_20_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_20_asid; // @[TLB.scala 64:31]
  reg  array4kb_21_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_21_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_21_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_21_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_21_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_21_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_21_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_21_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_21_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_21_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_21_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_21_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_21_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_21_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_21_asid; // @[TLB.scala 64:31]
  reg  array4kb_22_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_22_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_22_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_22_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_22_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_22_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_22_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_22_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_22_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_22_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_22_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_22_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_22_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_22_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_22_asid; // @[TLB.scala 64:31]
  reg  array4kb_23_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_23_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_23_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_23_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_23_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_23_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_23_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_23_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_23_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_23_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_23_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_23_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_23_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_23_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_23_asid; // @[TLB.scala 64:31]
  reg  array4kb_24_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_24_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_24_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_24_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_24_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_24_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_24_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_24_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_24_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_24_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_24_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_24_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_24_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_24_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_24_asid; // @[TLB.scala 64:31]
  reg  array4kb_25_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_25_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_25_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_25_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_25_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_25_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_25_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_25_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_25_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_25_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_25_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_25_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_25_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_25_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_25_asid; // @[TLB.scala 64:31]
  reg  array4kb_26_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_26_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_26_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_26_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_26_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_26_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_26_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_26_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_26_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_26_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_26_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_26_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_26_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_26_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_26_asid; // @[TLB.scala 64:31]
  reg  array4kb_27_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_27_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_27_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_27_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_27_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_27_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_27_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_27_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_27_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_27_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_27_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_27_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_27_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_27_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_27_asid; // @[TLB.scala 64:31]
  reg  array4kb_28_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_28_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_28_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_28_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_28_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_28_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_28_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_28_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_28_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_28_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_28_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_28_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_28_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_28_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_28_asid; // @[TLB.scala 64:31]
  reg  array4kb_29_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_29_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_29_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_29_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_29_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_29_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_29_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_29_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_29_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_29_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_29_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_29_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_29_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_29_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_29_asid; // @[TLB.scala 64:31]
  reg  array4kb_30_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_30_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_30_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_30_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_30_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_30_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_30_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_30_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_30_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_30_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_30_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_30_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_30_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_30_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_30_asid; // @[TLB.scala 64:31]
  reg  array4kb_31_flag_d; // @[TLB.scala 64:31]
  reg  array4kb_31_flag_a; // @[TLB.scala 64:31]
  reg  array4kb_31_flag_g; // @[TLB.scala 64:31]
  reg  array4kb_31_flag_u; // @[TLB.scala 64:31]
  reg  array4kb_31_flag_x; // @[TLB.scala 64:31]
  reg  array4kb_31_flag_w; // @[TLB.scala 64:31]
  reg  array4kb_31_flag_r; // @[TLB.scala 64:31]
  reg  array4kb_31_flag_v; // @[TLB.scala 64:31]
  reg [8:0] array4kb_31_vpn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_31_vpn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_31_vpn0; // @[TLB.scala 64:31]
  reg [1:0] array4kb_31_ppn2; // @[TLB.scala 64:31]
  reg [8:0] array4kb_31_ppn1; // @[TLB.scala 64:31]
  reg [8:0] array4kb_31_ppn0; // @[TLB.scala 64:31]
  reg [15:0] array4kb_31_asid; // @[TLB.scala 64:31]
  reg  array4kb_valid_0; // @[TLB.scala 65:31]
  reg  array4kb_valid_1; // @[TLB.scala 65:31]
  reg  array4kb_valid_2; // @[TLB.scala 65:31]
  reg  array4kb_valid_3; // @[TLB.scala 65:31]
  reg  array4kb_valid_4; // @[TLB.scala 65:31]
  reg  array4kb_valid_5; // @[TLB.scala 65:31]
  reg  array4kb_valid_6; // @[TLB.scala 65:31]
  reg  array4kb_valid_7; // @[TLB.scala 65:31]
  reg  array4kb_valid_8; // @[TLB.scala 65:31]
  reg  array4kb_valid_9; // @[TLB.scala 65:31]
  reg  array4kb_valid_10; // @[TLB.scala 65:31]
  reg  array4kb_valid_11; // @[TLB.scala 65:31]
  reg  array4kb_valid_12; // @[TLB.scala 65:31]
  reg  array4kb_valid_13; // @[TLB.scala 65:31]
  reg  array4kb_valid_14; // @[TLB.scala 65:31]
  reg  array4kb_valid_15; // @[TLB.scala 65:31]
  reg  array4kb_valid_16; // @[TLB.scala 65:31]
  reg  array4kb_valid_17; // @[TLB.scala 65:31]
  reg  array4kb_valid_18; // @[TLB.scala 65:31]
  reg  array4kb_valid_19; // @[TLB.scala 65:31]
  reg  array4kb_valid_20; // @[TLB.scala 65:31]
  reg  array4kb_valid_21; // @[TLB.scala 65:31]
  reg  array4kb_valid_22; // @[TLB.scala 65:31]
  reg  array4kb_valid_23; // @[TLB.scala 65:31]
  reg  array4kb_valid_24; // @[TLB.scala 65:31]
  reg  array4kb_valid_25; // @[TLB.scala 65:31]
  reg  array4kb_valid_26; // @[TLB.scala 65:31]
  reg  array4kb_valid_27; // @[TLB.scala 65:31]
  reg  array4kb_valid_28; // @[TLB.scala 65:31]
  reg  array4kb_valid_29; // @[TLB.scala 65:31]
  reg  array4kb_valid_30; // @[TLB.scala 65:31]
  reg  array4kb_valid_31; // @[TLB.scala 65:31]
  wire [26:0] _T_8 = {array4kb_0_vpn2,array4kb_0_vpn1,array4kb_0_vpn0}; // @[Cat.scala 33:92]
  wire [17:0] hi_1 = {io_vaddr_vpn2,io_vaddr_vpn1}; // @[Cat.scala 33:92]
  wire [26:0] _T_9 = {io_vaddr_vpn2,io_vaddr_vpn1,io_vaddr_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_0 = array4kb_valid_0 & _T_8 == _T_9 & (array4kb_0_asid == io_satp_asid | array4kb_0_flag_g); // @[TLB.scala 71:71 72:22 68:35]
  wire  _GEN_2 = array4kb_valid_0 & _T_8 == _T_9 & array4kb_0_flag_d; // @[TLB.scala 71:71 73:22 66:35]
  wire  _GEN_3 = array4kb_valid_0 & _T_8 == _T_9 & array4kb_0_flag_a; // @[TLB.scala 71:71 73:22 66:35]
  wire  _GEN_5 = array4kb_valid_0 & _T_8 == _T_9 & array4kb_0_flag_u; // @[TLB.scala 71:71 73:22 66:35]
  wire  _GEN_6 = array4kb_valid_0 & _T_8 == _T_9 & array4kb_0_flag_x; // @[TLB.scala 71:71 73:22 66:35]
  wire  _GEN_7 = array4kb_valid_0 & _T_8 == _T_9 & array4kb_0_flag_w; // @[TLB.scala 71:71 73:22 66:35]
  wire  _GEN_8 = array4kb_valid_0 & _T_8 == _T_9 & array4kb_0_flag_r; // @[TLB.scala 71:71 73:22 66:35]
  wire  _GEN_9 = array4kb_valid_0 & _T_8 == _T_9 & array4kb_0_flag_v; // @[TLB.scala 71:71 73:22 66:35]
  wire [1:0] _GEN_13 = array4kb_valid_0 & _T_8 == _T_9 ? array4kb_0_ppn2 : 2'h0; // @[TLB.scala 71:71 73:22 66:35]
  wire [8:0] _GEN_14 = array4kb_valid_0 & _T_8 == _T_9 ? array4kb_0_ppn1 : 9'h0; // @[TLB.scala 71:71 73:22 66:35]
  wire [8:0] _GEN_15 = array4kb_valid_0 & _T_8 == _T_9 ? array4kb_0_ppn0 : 9'h0; // @[TLB.scala 71:71 73:22 66:35]
  wire [26:0] _T_12 = {array4kb_1_vpn2,array4kb_1_vpn1,array4kb_1_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_17 = array4kb_valid_1 & _T_12 == _T_9 ? array4kb_1_asid == io_satp_asid | array4kb_1_flag_g : _GEN_0; // @[TLB.scala 71:71 72:22]
  wire  _GEN_19 = array4kb_valid_1 & _T_12 == _T_9 ? array4kb_1_flag_d : _GEN_2; // @[TLB.scala 71:71 73:22]
  wire  _GEN_20 = array4kb_valid_1 & _T_12 == _T_9 ? array4kb_1_flag_a : _GEN_3; // @[TLB.scala 71:71 73:22]
  wire  _GEN_22 = array4kb_valid_1 & _T_12 == _T_9 ? array4kb_1_flag_u : _GEN_5; // @[TLB.scala 71:71 73:22]
  wire  _GEN_23 = array4kb_valid_1 & _T_12 == _T_9 ? array4kb_1_flag_x : _GEN_6; // @[TLB.scala 71:71 73:22]
  wire  _GEN_24 = array4kb_valid_1 & _T_12 == _T_9 ? array4kb_1_flag_w : _GEN_7; // @[TLB.scala 71:71 73:22]
  wire  _GEN_25 = array4kb_valid_1 & _T_12 == _T_9 ? array4kb_1_flag_r : _GEN_8; // @[TLB.scala 71:71 73:22]
  wire  _GEN_26 = array4kb_valid_1 & _T_12 == _T_9 ? array4kb_1_flag_v : _GEN_9; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_30 = array4kb_valid_1 & _T_12 == _T_9 ? array4kb_1_ppn2 : _GEN_13; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_31 = array4kb_valid_1 & _T_12 == _T_9 ? array4kb_1_ppn1 : _GEN_14; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_32 = array4kb_valid_1 & _T_12 == _T_9 ? array4kb_1_ppn0 : _GEN_15; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_16 = {array4kb_2_vpn2,array4kb_2_vpn1,array4kb_2_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_34 = array4kb_valid_2 & _T_16 == _T_9 ? array4kb_2_asid == io_satp_asid | array4kb_2_flag_g : _GEN_17; // @[TLB.scala 71:71 72:22]
  wire  _GEN_36 = array4kb_valid_2 & _T_16 == _T_9 ? array4kb_2_flag_d : _GEN_19; // @[TLB.scala 71:71 73:22]
  wire  _GEN_37 = array4kb_valid_2 & _T_16 == _T_9 ? array4kb_2_flag_a : _GEN_20; // @[TLB.scala 71:71 73:22]
  wire  _GEN_39 = array4kb_valid_2 & _T_16 == _T_9 ? array4kb_2_flag_u : _GEN_22; // @[TLB.scala 71:71 73:22]
  wire  _GEN_40 = array4kb_valid_2 & _T_16 == _T_9 ? array4kb_2_flag_x : _GEN_23; // @[TLB.scala 71:71 73:22]
  wire  _GEN_41 = array4kb_valid_2 & _T_16 == _T_9 ? array4kb_2_flag_w : _GEN_24; // @[TLB.scala 71:71 73:22]
  wire  _GEN_42 = array4kb_valid_2 & _T_16 == _T_9 ? array4kb_2_flag_r : _GEN_25; // @[TLB.scala 71:71 73:22]
  wire  _GEN_43 = array4kb_valid_2 & _T_16 == _T_9 ? array4kb_2_flag_v : _GEN_26; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_47 = array4kb_valid_2 & _T_16 == _T_9 ? array4kb_2_ppn2 : _GEN_30; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_48 = array4kb_valid_2 & _T_16 == _T_9 ? array4kb_2_ppn1 : _GEN_31; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_49 = array4kb_valid_2 & _T_16 == _T_9 ? array4kb_2_ppn0 : _GEN_32; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_20 = {array4kb_3_vpn2,array4kb_3_vpn1,array4kb_3_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_51 = array4kb_valid_3 & _T_20 == _T_9 ? array4kb_3_asid == io_satp_asid | array4kb_3_flag_g : _GEN_34; // @[TLB.scala 71:71 72:22]
  wire  _GEN_53 = array4kb_valid_3 & _T_20 == _T_9 ? array4kb_3_flag_d : _GEN_36; // @[TLB.scala 71:71 73:22]
  wire  _GEN_54 = array4kb_valid_3 & _T_20 == _T_9 ? array4kb_3_flag_a : _GEN_37; // @[TLB.scala 71:71 73:22]
  wire  _GEN_56 = array4kb_valid_3 & _T_20 == _T_9 ? array4kb_3_flag_u : _GEN_39; // @[TLB.scala 71:71 73:22]
  wire  _GEN_57 = array4kb_valid_3 & _T_20 == _T_9 ? array4kb_3_flag_x : _GEN_40; // @[TLB.scala 71:71 73:22]
  wire  _GEN_58 = array4kb_valid_3 & _T_20 == _T_9 ? array4kb_3_flag_w : _GEN_41; // @[TLB.scala 71:71 73:22]
  wire  _GEN_59 = array4kb_valid_3 & _T_20 == _T_9 ? array4kb_3_flag_r : _GEN_42; // @[TLB.scala 71:71 73:22]
  wire  _GEN_60 = array4kb_valid_3 & _T_20 == _T_9 ? array4kb_3_flag_v : _GEN_43; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_64 = array4kb_valid_3 & _T_20 == _T_9 ? array4kb_3_ppn2 : _GEN_47; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_65 = array4kb_valid_3 & _T_20 == _T_9 ? array4kb_3_ppn1 : _GEN_48; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_66 = array4kb_valid_3 & _T_20 == _T_9 ? array4kb_3_ppn0 : _GEN_49; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_24 = {array4kb_4_vpn2,array4kb_4_vpn1,array4kb_4_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_68 = array4kb_valid_4 & _T_24 == _T_9 ? array4kb_4_asid == io_satp_asid | array4kb_4_flag_g : _GEN_51; // @[TLB.scala 71:71 72:22]
  wire  _GEN_70 = array4kb_valid_4 & _T_24 == _T_9 ? array4kb_4_flag_d : _GEN_53; // @[TLB.scala 71:71 73:22]
  wire  _GEN_71 = array4kb_valid_4 & _T_24 == _T_9 ? array4kb_4_flag_a : _GEN_54; // @[TLB.scala 71:71 73:22]
  wire  _GEN_73 = array4kb_valid_4 & _T_24 == _T_9 ? array4kb_4_flag_u : _GEN_56; // @[TLB.scala 71:71 73:22]
  wire  _GEN_74 = array4kb_valid_4 & _T_24 == _T_9 ? array4kb_4_flag_x : _GEN_57; // @[TLB.scala 71:71 73:22]
  wire  _GEN_75 = array4kb_valid_4 & _T_24 == _T_9 ? array4kb_4_flag_w : _GEN_58; // @[TLB.scala 71:71 73:22]
  wire  _GEN_76 = array4kb_valid_4 & _T_24 == _T_9 ? array4kb_4_flag_r : _GEN_59; // @[TLB.scala 71:71 73:22]
  wire  _GEN_77 = array4kb_valid_4 & _T_24 == _T_9 ? array4kb_4_flag_v : _GEN_60; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_81 = array4kb_valid_4 & _T_24 == _T_9 ? array4kb_4_ppn2 : _GEN_64; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_82 = array4kb_valid_4 & _T_24 == _T_9 ? array4kb_4_ppn1 : _GEN_65; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_83 = array4kb_valid_4 & _T_24 == _T_9 ? array4kb_4_ppn0 : _GEN_66; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_28 = {array4kb_5_vpn2,array4kb_5_vpn1,array4kb_5_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_85 = array4kb_valid_5 & _T_28 == _T_9 ? array4kb_5_asid == io_satp_asid | array4kb_5_flag_g : _GEN_68; // @[TLB.scala 71:71 72:22]
  wire  _GEN_87 = array4kb_valid_5 & _T_28 == _T_9 ? array4kb_5_flag_d : _GEN_70; // @[TLB.scala 71:71 73:22]
  wire  _GEN_88 = array4kb_valid_5 & _T_28 == _T_9 ? array4kb_5_flag_a : _GEN_71; // @[TLB.scala 71:71 73:22]
  wire  _GEN_90 = array4kb_valid_5 & _T_28 == _T_9 ? array4kb_5_flag_u : _GEN_73; // @[TLB.scala 71:71 73:22]
  wire  _GEN_91 = array4kb_valid_5 & _T_28 == _T_9 ? array4kb_5_flag_x : _GEN_74; // @[TLB.scala 71:71 73:22]
  wire  _GEN_92 = array4kb_valid_5 & _T_28 == _T_9 ? array4kb_5_flag_w : _GEN_75; // @[TLB.scala 71:71 73:22]
  wire  _GEN_93 = array4kb_valid_5 & _T_28 == _T_9 ? array4kb_5_flag_r : _GEN_76; // @[TLB.scala 71:71 73:22]
  wire  _GEN_94 = array4kb_valid_5 & _T_28 == _T_9 ? array4kb_5_flag_v : _GEN_77; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_98 = array4kb_valid_5 & _T_28 == _T_9 ? array4kb_5_ppn2 : _GEN_81; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_99 = array4kb_valid_5 & _T_28 == _T_9 ? array4kb_5_ppn1 : _GEN_82; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_100 = array4kb_valid_5 & _T_28 == _T_9 ? array4kb_5_ppn0 : _GEN_83; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_32 = {array4kb_6_vpn2,array4kb_6_vpn1,array4kb_6_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_102 = array4kb_valid_6 & _T_32 == _T_9 ? array4kb_6_asid == io_satp_asid | array4kb_6_flag_g : _GEN_85; // @[TLB.scala 71:71 72:22]
  wire  _GEN_104 = array4kb_valid_6 & _T_32 == _T_9 ? array4kb_6_flag_d : _GEN_87; // @[TLB.scala 71:71 73:22]
  wire  _GEN_105 = array4kb_valid_6 & _T_32 == _T_9 ? array4kb_6_flag_a : _GEN_88; // @[TLB.scala 71:71 73:22]
  wire  _GEN_107 = array4kb_valid_6 & _T_32 == _T_9 ? array4kb_6_flag_u : _GEN_90; // @[TLB.scala 71:71 73:22]
  wire  _GEN_108 = array4kb_valid_6 & _T_32 == _T_9 ? array4kb_6_flag_x : _GEN_91; // @[TLB.scala 71:71 73:22]
  wire  _GEN_109 = array4kb_valid_6 & _T_32 == _T_9 ? array4kb_6_flag_w : _GEN_92; // @[TLB.scala 71:71 73:22]
  wire  _GEN_110 = array4kb_valid_6 & _T_32 == _T_9 ? array4kb_6_flag_r : _GEN_93; // @[TLB.scala 71:71 73:22]
  wire  _GEN_111 = array4kb_valid_6 & _T_32 == _T_9 ? array4kb_6_flag_v : _GEN_94; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_115 = array4kb_valid_6 & _T_32 == _T_9 ? array4kb_6_ppn2 : _GEN_98; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_116 = array4kb_valid_6 & _T_32 == _T_9 ? array4kb_6_ppn1 : _GEN_99; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_117 = array4kb_valid_6 & _T_32 == _T_9 ? array4kb_6_ppn0 : _GEN_100; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_36 = {array4kb_7_vpn2,array4kb_7_vpn1,array4kb_7_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_119 = array4kb_valid_7 & _T_36 == _T_9 ? array4kb_7_asid == io_satp_asid | array4kb_7_flag_g : _GEN_102; // @[TLB.scala 71:71 72:22]
  wire  _GEN_121 = array4kb_valid_7 & _T_36 == _T_9 ? array4kb_7_flag_d : _GEN_104; // @[TLB.scala 71:71 73:22]
  wire  _GEN_122 = array4kb_valid_7 & _T_36 == _T_9 ? array4kb_7_flag_a : _GEN_105; // @[TLB.scala 71:71 73:22]
  wire  _GEN_124 = array4kb_valid_7 & _T_36 == _T_9 ? array4kb_7_flag_u : _GEN_107; // @[TLB.scala 71:71 73:22]
  wire  _GEN_125 = array4kb_valid_7 & _T_36 == _T_9 ? array4kb_7_flag_x : _GEN_108; // @[TLB.scala 71:71 73:22]
  wire  _GEN_126 = array4kb_valid_7 & _T_36 == _T_9 ? array4kb_7_flag_w : _GEN_109; // @[TLB.scala 71:71 73:22]
  wire  _GEN_127 = array4kb_valid_7 & _T_36 == _T_9 ? array4kb_7_flag_r : _GEN_110; // @[TLB.scala 71:71 73:22]
  wire  _GEN_128 = array4kb_valid_7 & _T_36 == _T_9 ? array4kb_7_flag_v : _GEN_111; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_132 = array4kb_valid_7 & _T_36 == _T_9 ? array4kb_7_ppn2 : _GEN_115; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_133 = array4kb_valid_7 & _T_36 == _T_9 ? array4kb_7_ppn1 : _GEN_116; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_134 = array4kb_valid_7 & _T_36 == _T_9 ? array4kb_7_ppn0 : _GEN_117; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_40 = {array4kb_8_vpn2,array4kb_8_vpn1,array4kb_8_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_136 = array4kb_valid_8 & _T_40 == _T_9 ? array4kb_8_asid == io_satp_asid | array4kb_8_flag_g : _GEN_119; // @[TLB.scala 71:71 72:22]
  wire  _GEN_138 = array4kb_valid_8 & _T_40 == _T_9 ? array4kb_8_flag_d : _GEN_121; // @[TLB.scala 71:71 73:22]
  wire  _GEN_139 = array4kb_valid_8 & _T_40 == _T_9 ? array4kb_8_flag_a : _GEN_122; // @[TLB.scala 71:71 73:22]
  wire  _GEN_141 = array4kb_valid_8 & _T_40 == _T_9 ? array4kb_8_flag_u : _GEN_124; // @[TLB.scala 71:71 73:22]
  wire  _GEN_142 = array4kb_valid_8 & _T_40 == _T_9 ? array4kb_8_flag_x : _GEN_125; // @[TLB.scala 71:71 73:22]
  wire  _GEN_143 = array4kb_valid_8 & _T_40 == _T_9 ? array4kb_8_flag_w : _GEN_126; // @[TLB.scala 71:71 73:22]
  wire  _GEN_144 = array4kb_valid_8 & _T_40 == _T_9 ? array4kb_8_flag_r : _GEN_127; // @[TLB.scala 71:71 73:22]
  wire  _GEN_145 = array4kb_valid_8 & _T_40 == _T_9 ? array4kb_8_flag_v : _GEN_128; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_149 = array4kb_valid_8 & _T_40 == _T_9 ? array4kb_8_ppn2 : _GEN_132; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_150 = array4kb_valid_8 & _T_40 == _T_9 ? array4kb_8_ppn1 : _GEN_133; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_151 = array4kb_valid_8 & _T_40 == _T_9 ? array4kb_8_ppn0 : _GEN_134; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_44 = {array4kb_9_vpn2,array4kb_9_vpn1,array4kb_9_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_153 = array4kb_valid_9 & _T_44 == _T_9 ? array4kb_9_asid == io_satp_asid | array4kb_9_flag_g : _GEN_136; // @[TLB.scala 71:71 72:22]
  wire  _GEN_155 = array4kb_valid_9 & _T_44 == _T_9 ? array4kb_9_flag_d : _GEN_138; // @[TLB.scala 71:71 73:22]
  wire  _GEN_156 = array4kb_valid_9 & _T_44 == _T_9 ? array4kb_9_flag_a : _GEN_139; // @[TLB.scala 71:71 73:22]
  wire  _GEN_158 = array4kb_valid_9 & _T_44 == _T_9 ? array4kb_9_flag_u : _GEN_141; // @[TLB.scala 71:71 73:22]
  wire  _GEN_159 = array4kb_valid_9 & _T_44 == _T_9 ? array4kb_9_flag_x : _GEN_142; // @[TLB.scala 71:71 73:22]
  wire  _GEN_160 = array4kb_valid_9 & _T_44 == _T_9 ? array4kb_9_flag_w : _GEN_143; // @[TLB.scala 71:71 73:22]
  wire  _GEN_161 = array4kb_valid_9 & _T_44 == _T_9 ? array4kb_9_flag_r : _GEN_144; // @[TLB.scala 71:71 73:22]
  wire  _GEN_162 = array4kb_valid_9 & _T_44 == _T_9 ? array4kb_9_flag_v : _GEN_145; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_166 = array4kb_valid_9 & _T_44 == _T_9 ? array4kb_9_ppn2 : _GEN_149; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_167 = array4kb_valid_9 & _T_44 == _T_9 ? array4kb_9_ppn1 : _GEN_150; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_168 = array4kb_valid_9 & _T_44 == _T_9 ? array4kb_9_ppn0 : _GEN_151; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_48 = {array4kb_10_vpn2,array4kb_10_vpn1,array4kb_10_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_170 = array4kb_valid_10 & _T_48 == _T_9 ? array4kb_10_asid == io_satp_asid | array4kb_10_flag_g : _GEN_153; // @[TLB.scala 71:71 72:22]
  wire  _GEN_172 = array4kb_valid_10 & _T_48 == _T_9 ? array4kb_10_flag_d : _GEN_155; // @[TLB.scala 71:71 73:22]
  wire  _GEN_173 = array4kb_valid_10 & _T_48 == _T_9 ? array4kb_10_flag_a : _GEN_156; // @[TLB.scala 71:71 73:22]
  wire  _GEN_175 = array4kb_valid_10 & _T_48 == _T_9 ? array4kb_10_flag_u : _GEN_158; // @[TLB.scala 71:71 73:22]
  wire  _GEN_176 = array4kb_valid_10 & _T_48 == _T_9 ? array4kb_10_flag_x : _GEN_159; // @[TLB.scala 71:71 73:22]
  wire  _GEN_177 = array4kb_valid_10 & _T_48 == _T_9 ? array4kb_10_flag_w : _GEN_160; // @[TLB.scala 71:71 73:22]
  wire  _GEN_178 = array4kb_valid_10 & _T_48 == _T_9 ? array4kb_10_flag_r : _GEN_161; // @[TLB.scala 71:71 73:22]
  wire  _GEN_179 = array4kb_valid_10 & _T_48 == _T_9 ? array4kb_10_flag_v : _GEN_162; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_183 = array4kb_valid_10 & _T_48 == _T_9 ? array4kb_10_ppn2 : _GEN_166; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_184 = array4kb_valid_10 & _T_48 == _T_9 ? array4kb_10_ppn1 : _GEN_167; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_185 = array4kb_valid_10 & _T_48 == _T_9 ? array4kb_10_ppn0 : _GEN_168; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_52 = {array4kb_11_vpn2,array4kb_11_vpn1,array4kb_11_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_187 = array4kb_valid_11 & _T_52 == _T_9 ? array4kb_11_asid == io_satp_asid | array4kb_11_flag_g : _GEN_170; // @[TLB.scala 71:71 72:22]
  wire  _GEN_189 = array4kb_valid_11 & _T_52 == _T_9 ? array4kb_11_flag_d : _GEN_172; // @[TLB.scala 71:71 73:22]
  wire  _GEN_190 = array4kb_valid_11 & _T_52 == _T_9 ? array4kb_11_flag_a : _GEN_173; // @[TLB.scala 71:71 73:22]
  wire  _GEN_192 = array4kb_valid_11 & _T_52 == _T_9 ? array4kb_11_flag_u : _GEN_175; // @[TLB.scala 71:71 73:22]
  wire  _GEN_193 = array4kb_valid_11 & _T_52 == _T_9 ? array4kb_11_flag_x : _GEN_176; // @[TLB.scala 71:71 73:22]
  wire  _GEN_194 = array4kb_valid_11 & _T_52 == _T_9 ? array4kb_11_flag_w : _GEN_177; // @[TLB.scala 71:71 73:22]
  wire  _GEN_195 = array4kb_valid_11 & _T_52 == _T_9 ? array4kb_11_flag_r : _GEN_178; // @[TLB.scala 71:71 73:22]
  wire  _GEN_196 = array4kb_valid_11 & _T_52 == _T_9 ? array4kb_11_flag_v : _GEN_179; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_200 = array4kb_valid_11 & _T_52 == _T_9 ? array4kb_11_ppn2 : _GEN_183; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_201 = array4kb_valid_11 & _T_52 == _T_9 ? array4kb_11_ppn1 : _GEN_184; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_202 = array4kb_valid_11 & _T_52 == _T_9 ? array4kb_11_ppn0 : _GEN_185; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_56 = {array4kb_12_vpn2,array4kb_12_vpn1,array4kb_12_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_204 = array4kb_valid_12 & _T_56 == _T_9 ? array4kb_12_asid == io_satp_asid | array4kb_12_flag_g : _GEN_187; // @[TLB.scala 71:71 72:22]
  wire  _GEN_206 = array4kb_valid_12 & _T_56 == _T_9 ? array4kb_12_flag_d : _GEN_189; // @[TLB.scala 71:71 73:22]
  wire  _GEN_207 = array4kb_valid_12 & _T_56 == _T_9 ? array4kb_12_flag_a : _GEN_190; // @[TLB.scala 71:71 73:22]
  wire  _GEN_209 = array4kb_valid_12 & _T_56 == _T_9 ? array4kb_12_flag_u : _GEN_192; // @[TLB.scala 71:71 73:22]
  wire  _GEN_210 = array4kb_valid_12 & _T_56 == _T_9 ? array4kb_12_flag_x : _GEN_193; // @[TLB.scala 71:71 73:22]
  wire  _GEN_211 = array4kb_valid_12 & _T_56 == _T_9 ? array4kb_12_flag_w : _GEN_194; // @[TLB.scala 71:71 73:22]
  wire  _GEN_212 = array4kb_valid_12 & _T_56 == _T_9 ? array4kb_12_flag_r : _GEN_195; // @[TLB.scala 71:71 73:22]
  wire  _GEN_213 = array4kb_valid_12 & _T_56 == _T_9 ? array4kb_12_flag_v : _GEN_196; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_217 = array4kb_valid_12 & _T_56 == _T_9 ? array4kb_12_ppn2 : _GEN_200; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_218 = array4kb_valid_12 & _T_56 == _T_9 ? array4kb_12_ppn1 : _GEN_201; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_219 = array4kb_valid_12 & _T_56 == _T_9 ? array4kb_12_ppn0 : _GEN_202; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_60 = {array4kb_13_vpn2,array4kb_13_vpn1,array4kb_13_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_221 = array4kb_valid_13 & _T_60 == _T_9 ? array4kb_13_asid == io_satp_asid | array4kb_13_flag_g : _GEN_204; // @[TLB.scala 71:71 72:22]
  wire  _GEN_223 = array4kb_valid_13 & _T_60 == _T_9 ? array4kb_13_flag_d : _GEN_206; // @[TLB.scala 71:71 73:22]
  wire  _GEN_224 = array4kb_valid_13 & _T_60 == _T_9 ? array4kb_13_flag_a : _GEN_207; // @[TLB.scala 71:71 73:22]
  wire  _GEN_226 = array4kb_valid_13 & _T_60 == _T_9 ? array4kb_13_flag_u : _GEN_209; // @[TLB.scala 71:71 73:22]
  wire  _GEN_227 = array4kb_valid_13 & _T_60 == _T_9 ? array4kb_13_flag_x : _GEN_210; // @[TLB.scala 71:71 73:22]
  wire  _GEN_228 = array4kb_valid_13 & _T_60 == _T_9 ? array4kb_13_flag_w : _GEN_211; // @[TLB.scala 71:71 73:22]
  wire  _GEN_229 = array4kb_valid_13 & _T_60 == _T_9 ? array4kb_13_flag_r : _GEN_212; // @[TLB.scala 71:71 73:22]
  wire  _GEN_230 = array4kb_valid_13 & _T_60 == _T_9 ? array4kb_13_flag_v : _GEN_213; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_234 = array4kb_valid_13 & _T_60 == _T_9 ? array4kb_13_ppn2 : _GEN_217; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_235 = array4kb_valid_13 & _T_60 == _T_9 ? array4kb_13_ppn1 : _GEN_218; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_236 = array4kb_valid_13 & _T_60 == _T_9 ? array4kb_13_ppn0 : _GEN_219; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_64 = {array4kb_14_vpn2,array4kb_14_vpn1,array4kb_14_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_238 = array4kb_valid_14 & _T_64 == _T_9 ? array4kb_14_asid == io_satp_asid | array4kb_14_flag_g : _GEN_221; // @[TLB.scala 71:71 72:22]
  wire  _GEN_240 = array4kb_valid_14 & _T_64 == _T_9 ? array4kb_14_flag_d : _GEN_223; // @[TLB.scala 71:71 73:22]
  wire  _GEN_241 = array4kb_valid_14 & _T_64 == _T_9 ? array4kb_14_flag_a : _GEN_224; // @[TLB.scala 71:71 73:22]
  wire  _GEN_243 = array4kb_valid_14 & _T_64 == _T_9 ? array4kb_14_flag_u : _GEN_226; // @[TLB.scala 71:71 73:22]
  wire  _GEN_244 = array4kb_valid_14 & _T_64 == _T_9 ? array4kb_14_flag_x : _GEN_227; // @[TLB.scala 71:71 73:22]
  wire  _GEN_245 = array4kb_valid_14 & _T_64 == _T_9 ? array4kb_14_flag_w : _GEN_228; // @[TLB.scala 71:71 73:22]
  wire  _GEN_246 = array4kb_valid_14 & _T_64 == _T_9 ? array4kb_14_flag_r : _GEN_229; // @[TLB.scala 71:71 73:22]
  wire  _GEN_247 = array4kb_valid_14 & _T_64 == _T_9 ? array4kb_14_flag_v : _GEN_230; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_251 = array4kb_valid_14 & _T_64 == _T_9 ? array4kb_14_ppn2 : _GEN_234; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_252 = array4kb_valid_14 & _T_64 == _T_9 ? array4kb_14_ppn1 : _GEN_235; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_253 = array4kb_valid_14 & _T_64 == _T_9 ? array4kb_14_ppn0 : _GEN_236; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_68 = {array4kb_15_vpn2,array4kb_15_vpn1,array4kb_15_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_255 = array4kb_valid_15 & _T_68 == _T_9 ? array4kb_15_asid == io_satp_asid | array4kb_15_flag_g : _GEN_238; // @[TLB.scala 71:71 72:22]
  wire  _GEN_257 = array4kb_valid_15 & _T_68 == _T_9 ? array4kb_15_flag_d : _GEN_240; // @[TLB.scala 71:71 73:22]
  wire  _GEN_258 = array4kb_valid_15 & _T_68 == _T_9 ? array4kb_15_flag_a : _GEN_241; // @[TLB.scala 71:71 73:22]
  wire  _GEN_260 = array4kb_valid_15 & _T_68 == _T_9 ? array4kb_15_flag_u : _GEN_243; // @[TLB.scala 71:71 73:22]
  wire  _GEN_261 = array4kb_valid_15 & _T_68 == _T_9 ? array4kb_15_flag_x : _GEN_244; // @[TLB.scala 71:71 73:22]
  wire  _GEN_262 = array4kb_valid_15 & _T_68 == _T_9 ? array4kb_15_flag_w : _GEN_245; // @[TLB.scala 71:71 73:22]
  wire  _GEN_263 = array4kb_valid_15 & _T_68 == _T_9 ? array4kb_15_flag_r : _GEN_246; // @[TLB.scala 71:71 73:22]
  wire  _GEN_264 = array4kb_valid_15 & _T_68 == _T_9 ? array4kb_15_flag_v : _GEN_247; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_268 = array4kb_valid_15 & _T_68 == _T_9 ? array4kb_15_ppn2 : _GEN_251; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_269 = array4kb_valid_15 & _T_68 == _T_9 ? array4kb_15_ppn1 : _GEN_252; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_270 = array4kb_valid_15 & _T_68 == _T_9 ? array4kb_15_ppn0 : _GEN_253; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_72 = {array4kb_16_vpn2,array4kb_16_vpn1,array4kb_16_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_272 = array4kb_valid_16 & _T_72 == _T_9 ? array4kb_16_asid == io_satp_asid | array4kb_16_flag_g : _GEN_255; // @[TLB.scala 71:71 72:22]
  wire  _GEN_274 = array4kb_valid_16 & _T_72 == _T_9 ? array4kb_16_flag_d : _GEN_257; // @[TLB.scala 71:71 73:22]
  wire  _GEN_275 = array4kb_valid_16 & _T_72 == _T_9 ? array4kb_16_flag_a : _GEN_258; // @[TLB.scala 71:71 73:22]
  wire  _GEN_277 = array4kb_valid_16 & _T_72 == _T_9 ? array4kb_16_flag_u : _GEN_260; // @[TLB.scala 71:71 73:22]
  wire  _GEN_278 = array4kb_valid_16 & _T_72 == _T_9 ? array4kb_16_flag_x : _GEN_261; // @[TLB.scala 71:71 73:22]
  wire  _GEN_279 = array4kb_valid_16 & _T_72 == _T_9 ? array4kb_16_flag_w : _GEN_262; // @[TLB.scala 71:71 73:22]
  wire  _GEN_280 = array4kb_valid_16 & _T_72 == _T_9 ? array4kb_16_flag_r : _GEN_263; // @[TLB.scala 71:71 73:22]
  wire  _GEN_281 = array4kb_valid_16 & _T_72 == _T_9 ? array4kb_16_flag_v : _GEN_264; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_285 = array4kb_valid_16 & _T_72 == _T_9 ? array4kb_16_ppn2 : _GEN_268; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_286 = array4kb_valid_16 & _T_72 == _T_9 ? array4kb_16_ppn1 : _GEN_269; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_287 = array4kb_valid_16 & _T_72 == _T_9 ? array4kb_16_ppn0 : _GEN_270; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_76 = {array4kb_17_vpn2,array4kb_17_vpn1,array4kb_17_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_289 = array4kb_valid_17 & _T_76 == _T_9 ? array4kb_17_asid == io_satp_asid | array4kb_17_flag_g : _GEN_272; // @[TLB.scala 71:71 72:22]
  wire  _GEN_291 = array4kb_valid_17 & _T_76 == _T_9 ? array4kb_17_flag_d : _GEN_274; // @[TLB.scala 71:71 73:22]
  wire  _GEN_292 = array4kb_valid_17 & _T_76 == _T_9 ? array4kb_17_flag_a : _GEN_275; // @[TLB.scala 71:71 73:22]
  wire  _GEN_294 = array4kb_valid_17 & _T_76 == _T_9 ? array4kb_17_flag_u : _GEN_277; // @[TLB.scala 71:71 73:22]
  wire  _GEN_295 = array4kb_valid_17 & _T_76 == _T_9 ? array4kb_17_flag_x : _GEN_278; // @[TLB.scala 71:71 73:22]
  wire  _GEN_296 = array4kb_valid_17 & _T_76 == _T_9 ? array4kb_17_flag_w : _GEN_279; // @[TLB.scala 71:71 73:22]
  wire  _GEN_297 = array4kb_valid_17 & _T_76 == _T_9 ? array4kb_17_flag_r : _GEN_280; // @[TLB.scala 71:71 73:22]
  wire  _GEN_298 = array4kb_valid_17 & _T_76 == _T_9 ? array4kb_17_flag_v : _GEN_281; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_302 = array4kb_valid_17 & _T_76 == _T_9 ? array4kb_17_ppn2 : _GEN_285; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_303 = array4kb_valid_17 & _T_76 == _T_9 ? array4kb_17_ppn1 : _GEN_286; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_304 = array4kb_valid_17 & _T_76 == _T_9 ? array4kb_17_ppn0 : _GEN_287; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_80 = {array4kb_18_vpn2,array4kb_18_vpn1,array4kb_18_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_306 = array4kb_valid_18 & _T_80 == _T_9 ? array4kb_18_asid == io_satp_asid | array4kb_18_flag_g : _GEN_289; // @[TLB.scala 71:71 72:22]
  wire  _GEN_308 = array4kb_valid_18 & _T_80 == _T_9 ? array4kb_18_flag_d : _GEN_291; // @[TLB.scala 71:71 73:22]
  wire  _GEN_309 = array4kb_valid_18 & _T_80 == _T_9 ? array4kb_18_flag_a : _GEN_292; // @[TLB.scala 71:71 73:22]
  wire  _GEN_311 = array4kb_valid_18 & _T_80 == _T_9 ? array4kb_18_flag_u : _GEN_294; // @[TLB.scala 71:71 73:22]
  wire  _GEN_312 = array4kb_valid_18 & _T_80 == _T_9 ? array4kb_18_flag_x : _GEN_295; // @[TLB.scala 71:71 73:22]
  wire  _GEN_313 = array4kb_valid_18 & _T_80 == _T_9 ? array4kb_18_flag_w : _GEN_296; // @[TLB.scala 71:71 73:22]
  wire  _GEN_314 = array4kb_valid_18 & _T_80 == _T_9 ? array4kb_18_flag_r : _GEN_297; // @[TLB.scala 71:71 73:22]
  wire  _GEN_315 = array4kb_valid_18 & _T_80 == _T_9 ? array4kb_18_flag_v : _GEN_298; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_319 = array4kb_valid_18 & _T_80 == _T_9 ? array4kb_18_ppn2 : _GEN_302; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_320 = array4kb_valid_18 & _T_80 == _T_9 ? array4kb_18_ppn1 : _GEN_303; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_321 = array4kb_valid_18 & _T_80 == _T_9 ? array4kb_18_ppn0 : _GEN_304; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_84 = {array4kb_19_vpn2,array4kb_19_vpn1,array4kb_19_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_323 = array4kb_valid_19 & _T_84 == _T_9 ? array4kb_19_asid == io_satp_asid | array4kb_19_flag_g : _GEN_306; // @[TLB.scala 71:71 72:22]
  wire  _GEN_325 = array4kb_valid_19 & _T_84 == _T_9 ? array4kb_19_flag_d : _GEN_308; // @[TLB.scala 71:71 73:22]
  wire  _GEN_326 = array4kb_valid_19 & _T_84 == _T_9 ? array4kb_19_flag_a : _GEN_309; // @[TLB.scala 71:71 73:22]
  wire  _GEN_328 = array4kb_valid_19 & _T_84 == _T_9 ? array4kb_19_flag_u : _GEN_311; // @[TLB.scala 71:71 73:22]
  wire  _GEN_329 = array4kb_valid_19 & _T_84 == _T_9 ? array4kb_19_flag_x : _GEN_312; // @[TLB.scala 71:71 73:22]
  wire  _GEN_330 = array4kb_valid_19 & _T_84 == _T_9 ? array4kb_19_flag_w : _GEN_313; // @[TLB.scala 71:71 73:22]
  wire  _GEN_331 = array4kb_valid_19 & _T_84 == _T_9 ? array4kb_19_flag_r : _GEN_314; // @[TLB.scala 71:71 73:22]
  wire  _GEN_332 = array4kb_valid_19 & _T_84 == _T_9 ? array4kb_19_flag_v : _GEN_315; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_336 = array4kb_valid_19 & _T_84 == _T_9 ? array4kb_19_ppn2 : _GEN_319; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_337 = array4kb_valid_19 & _T_84 == _T_9 ? array4kb_19_ppn1 : _GEN_320; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_338 = array4kb_valid_19 & _T_84 == _T_9 ? array4kb_19_ppn0 : _GEN_321; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_88 = {array4kb_20_vpn2,array4kb_20_vpn1,array4kb_20_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_340 = array4kb_valid_20 & _T_88 == _T_9 ? array4kb_20_asid == io_satp_asid | array4kb_20_flag_g : _GEN_323; // @[TLB.scala 71:71 72:22]
  wire  _GEN_342 = array4kb_valid_20 & _T_88 == _T_9 ? array4kb_20_flag_d : _GEN_325; // @[TLB.scala 71:71 73:22]
  wire  _GEN_343 = array4kb_valid_20 & _T_88 == _T_9 ? array4kb_20_flag_a : _GEN_326; // @[TLB.scala 71:71 73:22]
  wire  _GEN_345 = array4kb_valid_20 & _T_88 == _T_9 ? array4kb_20_flag_u : _GEN_328; // @[TLB.scala 71:71 73:22]
  wire  _GEN_346 = array4kb_valid_20 & _T_88 == _T_9 ? array4kb_20_flag_x : _GEN_329; // @[TLB.scala 71:71 73:22]
  wire  _GEN_347 = array4kb_valid_20 & _T_88 == _T_9 ? array4kb_20_flag_w : _GEN_330; // @[TLB.scala 71:71 73:22]
  wire  _GEN_348 = array4kb_valid_20 & _T_88 == _T_9 ? array4kb_20_flag_r : _GEN_331; // @[TLB.scala 71:71 73:22]
  wire  _GEN_349 = array4kb_valid_20 & _T_88 == _T_9 ? array4kb_20_flag_v : _GEN_332; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_353 = array4kb_valid_20 & _T_88 == _T_9 ? array4kb_20_ppn2 : _GEN_336; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_354 = array4kb_valid_20 & _T_88 == _T_9 ? array4kb_20_ppn1 : _GEN_337; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_355 = array4kb_valid_20 & _T_88 == _T_9 ? array4kb_20_ppn0 : _GEN_338; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_92 = {array4kb_21_vpn2,array4kb_21_vpn1,array4kb_21_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_357 = array4kb_valid_21 & _T_92 == _T_9 ? array4kb_21_asid == io_satp_asid | array4kb_21_flag_g : _GEN_340; // @[TLB.scala 71:71 72:22]
  wire  _GEN_359 = array4kb_valid_21 & _T_92 == _T_9 ? array4kb_21_flag_d : _GEN_342; // @[TLB.scala 71:71 73:22]
  wire  _GEN_360 = array4kb_valid_21 & _T_92 == _T_9 ? array4kb_21_flag_a : _GEN_343; // @[TLB.scala 71:71 73:22]
  wire  _GEN_362 = array4kb_valid_21 & _T_92 == _T_9 ? array4kb_21_flag_u : _GEN_345; // @[TLB.scala 71:71 73:22]
  wire  _GEN_363 = array4kb_valid_21 & _T_92 == _T_9 ? array4kb_21_flag_x : _GEN_346; // @[TLB.scala 71:71 73:22]
  wire  _GEN_364 = array4kb_valid_21 & _T_92 == _T_9 ? array4kb_21_flag_w : _GEN_347; // @[TLB.scala 71:71 73:22]
  wire  _GEN_365 = array4kb_valid_21 & _T_92 == _T_9 ? array4kb_21_flag_r : _GEN_348; // @[TLB.scala 71:71 73:22]
  wire  _GEN_366 = array4kb_valid_21 & _T_92 == _T_9 ? array4kb_21_flag_v : _GEN_349; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_370 = array4kb_valid_21 & _T_92 == _T_9 ? array4kb_21_ppn2 : _GEN_353; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_371 = array4kb_valid_21 & _T_92 == _T_9 ? array4kb_21_ppn1 : _GEN_354; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_372 = array4kb_valid_21 & _T_92 == _T_9 ? array4kb_21_ppn0 : _GEN_355; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_96 = {array4kb_22_vpn2,array4kb_22_vpn1,array4kb_22_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_374 = array4kb_valid_22 & _T_96 == _T_9 ? array4kb_22_asid == io_satp_asid | array4kb_22_flag_g : _GEN_357; // @[TLB.scala 71:71 72:22]
  wire  _GEN_376 = array4kb_valid_22 & _T_96 == _T_9 ? array4kb_22_flag_d : _GEN_359; // @[TLB.scala 71:71 73:22]
  wire  _GEN_377 = array4kb_valid_22 & _T_96 == _T_9 ? array4kb_22_flag_a : _GEN_360; // @[TLB.scala 71:71 73:22]
  wire  _GEN_379 = array4kb_valid_22 & _T_96 == _T_9 ? array4kb_22_flag_u : _GEN_362; // @[TLB.scala 71:71 73:22]
  wire  _GEN_380 = array4kb_valid_22 & _T_96 == _T_9 ? array4kb_22_flag_x : _GEN_363; // @[TLB.scala 71:71 73:22]
  wire  _GEN_381 = array4kb_valid_22 & _T_96 == _T_9 ? array4kb_22_flag_w : _GEN_364; // @[TLB.scala 71:71 73:22]
  wire  _GEN_382 = array4kb_valid_22 & _T_96 == _T_9 ? array4kb_22_flag_r : _GEN_365; // @[TLB.scala 71:71 73:22]
  wire  _GEN_383 = array4kb_valid_22 & _T_96 == _T_9 ? array4kb_22_flag_v : _GEN_366; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_387 = array4kb_valid_22 & _T_96 == _T_9 ? array4kb_22_ppn2 : _GEN_370; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_388 = array4kb_valid_22 & _T_96 == _T_9 ? array4kb_22_ppn1 : _GEN_371; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_389 = array4kb_valid_22 & _T_96 == _T_9 ? array4kb_22_ppn0 : _GEN_372; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_100 = {array4kb_23_vpn2,array4kb_23_vpn1,array4kb_23_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_391 = array4kb_valid_23 & _T_100 == _T_9 ? array4kb_23_asid == io_satp_asid | array4kb_23_flag_g : _GEN_374
    ; // @[TLB.scala 71:71 72:22]
  wire  _GEN_393 = array4kb_valid_23 & _T_100 == _T_9 ? array4kb_23_flag_d : _GEN_376; // @[TLB.scala 71:71 73:22]
  wire  _GEN_394 = array4kb_valid_23 & _T_100 == _T_9 ? array4kb_23_flag_a : _GEN_377; // @[TLB.scala 71:71 73:22]
  wire  _GEN_396 = array4kb_valid_23 & _T_100 == _T_9 ? array4kb_23_flag_u : _GEN_379; // @[TLB.scala 71:71 73:22]
  wire  _GEN_397 = array4kb_valid_23 & _T_100 == _T_9 ? array4kb_23_flag_x : _GEN_380; // @[TLB.scala 71:71 73:22]
  wire  _GEN_398 = array4kb_valid_23 & _T_100 == _T_9 ? array4kb_23_flag_w : _GEN_381; // @[TLB.scala 71:71 73:22]
  wire  _GEN_399 = array4kb_valid_23 & _T_100 == _T_9 ? array4kb_23_flag_r : _GEN_382; // @[TLB.scala 71:71 73:22]
  wire  _GEN_400 = array4kb_valid_23 & _T_100 == _T_9 ? array4kb_23_flag_v : _GEN_383; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_404 = array4kb_valid_23 & _T_100 == _T_9 ? array4kb_23_ppn2 : _GEN_387; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_405 = array4kb_valid_23 & _T_100 == _T_9 ? array4kb_23_ppn1 : _GEN_388; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_406 = array4kb_valid_23 & _T_100 == _T_9 ? array4kb_23_ppn0 : _GEN_389; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_104 = {array4kb_24_vpn2,array4kb_24_vpn1,array4kb_24_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_408 = array4kb_valid_24 & _T_104 == _T_9 ? array4kb_24_asid == io_satp_asid | array4kb_24_flag_g : _GEN_391
    ; // @[TLB.scala 71:71 72:22]
  wire  _GEN_410 = array4kb_valid_24 & _T_104 == _T_9 ? array4kb_24_flag_d : _GEN_393; // @[TLB.scala 71:71 73:22]
  wire  _GEN_411 = array4kb_valid_24 & _T_104 == _T_9 ? array4kb_24_flag_a : _GEN_394; // @[TLB.scala 71:71 73:22]
  wire  _GEN_413 = array4kb_valid_24 & _T_104 == _T_9 ? array4kb_24_flag_u : _GEN_396; // @[TLB.scala 71:71 73:22]
  wire  _GEN_414 = array4kb_valid_24 & _T_104 == _T_9 ? array4kb_24_flag_x : _GEN_397; // @[TLB.scala 71:71 73:22]
  wire  _GEN_415 = array4kb_valid_24 & _T_104 == _T_9 ? array4kb_24_flag_w : _GEN_398; // @[TLB.scala 71:71 73:22]
  wire  _GEN_416 = array4kb_valid_24 & _T_104 == _T_9 ? array4kb_24_flag_r : _GEN_399; // @[TLB.scala 71:71 73:22]
  wire  _GEN_417 = array4kb_valid_24 & _T_104 == _T_9 ? array4kb_24_flag_v : _GEN_400; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_421 = array4kb_valid_24 & _T_104 == _T_9 ? array4kb_24_ppn2 : _GEN_404; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_422 = array4kb_valid_24 & _T_104 == _T_9 ? array4kb_24_ppn1 : _GEN_405; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_423 = array4kb_valid_24 & _T_104 == _T_9 ? array4kb_24_ppn0 : _GEN_406; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_108 = {array4kb_25_vpn2,array4kb_25_vpn1,array4kb_25_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_425 = array4kb_valid_25 & _T_108 == _T_9 ? array4kb_25_asid == io_satp_asid | array4kb_25_flag_g : _GEN_408
    ; // @[TLB.scala 71:71 72:22]
  wire  _GEN_427 = array4kb_valid_25 & _T_108 == _T_9 ? array4kb_25_flag_d : _GEN_410; // @[TLB.scala 71:71 73:22]
  wire  _GEN_428 = array4kb_valid_25 & _T_108 == _T_9 ? array4kb_25_flag_a : _GEN_411; // @[TLB.scala 71:71 73:22]
  wire  _GEN_430 = array4kb_valid_25 & _T_108 == _T_9 ? array4kb_25_flag_u : _GEN_413; // @[TLB.scala 71:71 73:22]
  wire  _GEN_431 = array4kb_valid_25 & _T_108 == _T_9 ? array4kb_25_flag_x : _GEN_414; // @[TLB.scala 71:71 73:22]
  wire  _GEN_432 = array4kb_valid_25 & _T_108 == _T_9 ? array4kb_25_flag_w : _GEN_415; // @[TLB.scala 71:71 73:22]
  wire  _GEN_433 = array4kb_valid_25 & _T_108 == _T_9 ? array4kb_25_flag_r : _GEN_416; // @[TLB.scala 71:71 73:22]
  wire  _GEN_434 = array4kb_valid_25 & _T_108 == _T_9 ? array4kb_25_flag_v : _GEN_417; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_438 = array4kb_valid_25 & _T_108 == _T_9 ? array4kb_25_ppn2 : _GEN_421; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_439 = array4kb_valid_25 & _T_108 == _T_9 ? array4kb_25_ppn1 : _GEN_422; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_440 = array4kb_valid_25 & _T_108 == _T_9 ? array4kb_25_ppn0 : _GEN_423; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_112 = {array4kb_26_vpn2,array4kb_26_vpn1,array4kb_26_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_442 = array4kb_valid_26 & _T_112 == _T_9 ? array4kb_26_asid == io_satp_asid | array4kb_26_flag_g : _GEN_425
    ; // @[TLB.scala 71:71 72:22]
  wire  _GEN_444 = array4kb_valid_26 & _T_112 == _T_9 ? array4kb_26_flag_d : _GEN_427; // @[TLB.scala 71:71 73:22]
  wire  _GEN_445 = array4kb_valid_26 & _T_112 == _T_9 ? array4kb_26_flag_a : _GEN_428; // @[TLB.scala 71:71 73:22]
  wire  _GEN_447 = array4kb_valid_26 & _T_112 == _T_9 ? array4kb_26_flag_u : _GEN_430; // @[TLB.scala 71:71 73:22]
  wire  _GEN_448 = array4kb_valid_26 & _T_112 == _T_9 ? array4kb_26_flag_x : _GEN_431; // @[TLB.scala 71:71 73:22]
  wire  _GEN_449 = array4kb_valid_26 & _T_112 == _T_9 ? array4kb_26_flag_w : _GEN_432; // @[TLB.scala 71:71 73:22]
  wire  _GEN_450 = array4kb_valid_26 & _T_112 == _T_9 ? array4kb_26_flag_r : _GEN_433; // @[TLB.scala 71:71 73:22]
  wire  _GEN_451 = array4kb_valid_26 & _T_112 == _T_9 ? array4kb_26_flag_v : _GEN_434; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_455 = array4kb_valid_26 & _T_112 == _T_9 ? array4kb_26_ppn2 : _GEN_438; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_456 = array4kb_valid_26 & _T_112 == _T_9 ? array4kb_26_ppn1 : _GEN_439; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_457 = array4kb_valid_26 & _T_112 == _T_9 ? array4kb_26_ppn0 : _GEN_440; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_116 = {array4kb_27_vpn2,array4kb_27_vpn1,array4kb_27_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_459 = array4kb_valid_27 & _T_116 == _T_9 ? array4kb_27_asid == io_satp_asid | array4kb_27_flag_g : _GEN_442
    ; // @[TLB.scala 71:71 72:22]
  wire  _GEN_461 = array4kb_valid_27 & _T_116 == _T_9 ? array4kb_27_flag_d : _GEN_444; // @[TLB.scala 71:71 73:22]
  wire  _GEN_462 = array4kb_valid_27 & _T_116 == _T_9 ? array4kb_27_flag_a : _GEN_445; // @[TLB.scala 71:71 73:22]
  wire  _GEN_464 = array4kb_valid_27 & _T_116 == _T_9 ? array4kb_27_flag_u : _GEN_447; // @[TLB.scala 71:71 73:22]
  wire  _GEN_465 = array4kb_valid_27 & _T_116 == _T_9 ? array4kb_27_flag_x : _GEN_448; // @[TLB.scala 71:71 73:22]
  wire  _GEN_466 = array4kb_valid_27 & _T_116 == _T_9 ? array4kb_27_flag_w : _GEN_449; // @[TLB.scala 71:71 73:22]
  wire  _GEN_467 = array4kb_valid_27 & _T_116 == _T_9 ? array4kb_27_flag_r : _GEN_450; // @[TLB.scala 71:71 73:22]
  wire  _GEN_468 = array4kb_valid_27 & _T_116 == _T_9 ? array4kb_27_flag_v : _GEN_451; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_472 = array4kb_valid_27 & _T_116 == _T_9 ? array4kb_27_ppn2 : _GEN_455; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_473 = array4kb_valid_27 & _T_116 == _T_9 ? array4kb_27_ppn1 : _GEN_456; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_474 = array4kb_valid_27 & _T_116 == _T_9 ? array4kb_27_ppn0 : _GEN_457; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_120 = {array4kb_28_vpn2,array4kb_28_vpn1,array4kb_28_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_476 = array4kb_valid_28 & _T_120 == _T_9 ? array4kb_28_asid == io_satp_asid | array4kb_28_flag_g : _GEN_459
    ; // @[TLB.scala 71:71 72:22]
  wire  _GEN_478 = array4kb_valid_28 & _T_120 == _T_9 ? array4kb_28_flag_d : _GEN_461; // @[TLB.scala 71:71 73:22]
  wire  _GEN_479 = array4kb_valid_28 & _T_120 == _T_9 ? array4kb_28_flag_a : _GEN_462; // @[TLB.scala 71:71 73:22]
  wire  _GEN_481 = array4kb_valid_28 & _T_120 == _T_9 ? array4kb_28_flag_u : _GEN_464; // @[TLB.scala 71:71 73:22]
  wire  _GEN_482 = array4kb_valid_28 & _T_120 == _T_9 ? array4kb_28_flag_x : _GEN_465; // @[TLB.scala 71:71 73:22]
  wire  _GEN_483 = array4kb_valid_28 & _T_120 == _T_9 ? array4kb_28_flag_w : _GEN_466; // @[TLB.scala 71:71 73:22]
  wire  _GEN_484 = array4kb_valid_28 & _T_120 == _T_9 ? array4kb_28_flag_r : _GEN_467; // @[TLB.scala 71:71 73:22]
  wire  _GEN_485 = array4kb_valid_28 & _T_120 == _T_9 ? array4kb_28_flag_v : _GEN_468; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_489 = array4kb_valid_28 & _T_120 == _T_9 ? array4kb_28_ppn2 : _GEN_472; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_490 = array4kb_valid_28 & _T_120 == _T_9 ? array4kb_28_ppn1 : _GEN_473; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_491 = array4kb_valid_28 & _T_120 == _T_9 ? array4kb_28_ppn0 : _GEN_474; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_124 = {array4kb_29_vpn2,array4kb_29_vpn1,array4kb_29_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_493 = array4kb_valid_29 & _T_124 == _T_9 ? array4kb_29_asid == io_satp_asid | array4kb_29_flag_g : _GEN_476
    ; // @[TLB.scala 71:71 72:22]
  wire  _GEN_495 = array4kb_valid_29 & _T_124 == _T_9 ? array4kb_29_flag_d : _GEN_478; // @[TLB.scala 71:71 73:22]
  wire  _GEN_496 = array4kb_valid_29 & _T_124 == _T_9 ? array4kb_29_flag_a : _GEN_479; // @[TLB.scala 71:71 73:22]
  wire  _GEN_498 = array4kb_valid_29 & _T_124 == _T_9 ? array4kb_29_flag_u : _GEN_481; // @[TLB.scala 71:71 73:22]
  wire  _GEN_499 = array4kb_valid_29 & _T_124 == _T_9 ? array4kb_29_flag_x : _GEN_482; // @[TLB.scala 71:71 73:22]
  wire  _GEN_500 = array4kb_valid_29 & _T_124 == _T_9 ? array4kb_29_flag_w : _GEN_483; // @[TLB.scala 71:71 73:22]
  wire  _GEN_501 = array4kb_valid_29 & _T_124 == _T_9 ? array4kb_29_flag_r : _GEN_484; // @[TLB.scala 71:71 73:22]
  wire  _GEN_502 = array4kb_valid_29 & _T_124 == _T_9 ? array4kb_29_flag_v : _GEN_485; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_506 = array4kb_valid_29 & _T_124 == _T_9 ? array4kb_29_ppn2 : _GEN_489; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_507 = array4kb_valid_29 & _T_124 == _T_9 ? array4kb_29_ppn1 : _GEN_490; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_508 = array4kb_valid_29 & _T_124 == _T_9 ? array4kb_29_ppn0 : _GEN_491; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_128 = {array4kb_30_vpn2,array4kb_30_vpn1,array4kb_30_vpn0}; // @[Cat.scala 33:92]
  wire  _GEN_510 = array4kb_valid_30 & _T_128 == _T_9 ? array4kb_30_asid == io_satp_asid | array4kb_30_flag_g : _GEN_493
    ; // @[TLB.scala 71:71 72:22]
  wire  _GEN_512 = array4kb_valid_30 & _T_128 == _T_9 ? array4kb_30_flag_d : _GEN_495; // @[TLB.scala 71:71 73:22]
  wire  _GEN_513 = array4kb_valid_30 & _T_128 == _T_9 ? array4kb_30_flag_a : _GEN_496; // @[TLB.scala 71:71 73:22]
  wire  _GEN_515 = array4kb_valid_30 & _T_128 == _T_9 ? array4kb_30_flag_u : _GEN_498; // @[TLB.scala 71:71 73:22]
  wire  _GEN_516 = array4kb_valid_30 & _T_128 == _T_9 ? array4kb_30_flag_x : _GEN_499; // @[TLB.scala 71:71 73:22]
  wire  _GEN_517 = array4kb_valid_30 & _T_128 == _T_9 ? array4kb_30_flag_w : _GEN_500; // @[TLB.scala 71:71 73:22]
  wire  _GEN_518 = array4kb_valid_30 & _T_128 == _T_9 ? array4kb_30_flag_r : _GEN_501; // @[TLB.scala 71:71 73:22]
  wire  _GEN_519 = array4kb_valid_30 & _T_128 == _T_9 ? array4kb_30_flag_v : _GEN_502; // @[TLB.scala 71:71 73:22]
  wire [1:0] _GEN_523 = array4kb_valid_30 & _T_128 == _T_9 ? array4kb_30_ppn2 : _GEN_506; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_524 = array4kb_valid_30 & _T_128 == _T_9 ? array4kb_30_ppn1 : _GEN_507; // @[TLB.scala 71:71 73:22]
  wire [8:0] _GEN_525 = array4kb_valid_30 & _T_128 == _T_9 ? array4kb_30_ppn0 : _GEN_508; // @[TLB.scala 71:71 73:22]
  wire [26:0] _T_132 = {array4kb_31_vpn2,array4kb_31_vpn1,array4kb_31_vpn0}; // @[Cat.scala 33:92]
  wire  hit4kb = array4kb_valid_31 & _T_132 == _T_9 ? array4kb_31_asid == io_satp_asid | array4kb_31_flag_g : _GEN_510; // @[TLB.scala 71:71 72:22]
  wire  array4kb_rdata_flag_d = array4kb_valid_31 & _T_132 == _T_9 ? array4kb_31_flag_d : _GEN_512; // @[TLB.scala 71:71 73:22]
  wire  array4kb_rdata_flag_a = array4kb_valid_31 & _T_132 == _T_9 ? array4kb_31_flag_a : _GEN_513; // @[TLB.scala 71:71 73:22]
  wire  array4kb_rdata_flag_u = array4kb_valid_31 & _T_132 == _T_9 ? array4kb_31_flag_u : _GEN_515; // @[TLB.scala 71:71 73:22]
  wire  array4kb_rdata_flag_x = array4kb_valid_31 & _T_132 == _T_9 ? array4kb_31_flag_x : _GEN_516; // @[TLB.scala 71:71 73:22]
  wire  array4kb_rdata_flag_w = array4kb_valid_31 & _T_132 == _T_9 ? array4kb_31_flag_w : _GEN_517; // @[TLB.scala 71:71 73:22]
  wire  array4kb_rdata_flag_r = array4kb_valid_31 & _T_132 == _T_9 ? array4kb_31_flag_r : _GEN_518; // @[TLB.scala 71:71 73:22]
  wire  array4kb_rdata_flag_v = array4kb_valid_31 & _T_132 == _T_9 ? array4kb_31_flag_v : _GEN_519; // @[TLB.scala 71:71 73:22]
  wire [1:0] array4kb_rdata_ppn2 = array4kb_valid_31 & _T_132 == _T_9 ? array4kb_31_ppn2 : _GEN_523; // @[TLB.scala 71:71 73:22]
  wire [8:0] array4kb_rdata_ppn1 = array4kb_valid_31 & _T_132 == _T_9 ? array4kb_31_ppn1 : _GEN_524; // @[TLB.scala 71:71 73:22]
  wire [8:0] array4kb_rdata_ppn0 = array4kb_valid_31 & _T_132 == _T_9 ? array4kb_31_ppn0 : _GEN_525; // @[TLB.scala 71:71 73:22]
  wire  _GEN_1056 = 5'h0 == replace_idx | array4kb_valid_0; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1057 = 5'h1 == replace_idx | array4kb_valid_1; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1058 = 5'h2 == replace_idx | array4kb_valid_2; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1059 = 5'h3 == replace_idx | array4kb_valid_3; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1060 = 5'h4 == replace_idx | array4kb_valid_4; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1061 = 5'h5 == replace_idx | array4kb_valid_5; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1062 = 5'h6 == replace_idx | array4kb_valid_6; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1063 = 5'h7 == replace_idx | array4kb_valid_7; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1064 = 5'h8 == replace_idx | array4kb_valid_8; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1065 = 5'h9 == replace_idx | array4kb_valid_9; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1066 = 5'ha == replace_idx | array4kb_valid_10; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1067 = 5'hb == replace_idx | array4kb_valid_11; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1068 = 5'hc == replace_idx | array4kb_valid_12; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1069 = 5'hd == replace_idx | array4kb_valid_13; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1070 = 5'he == replace_idx | array4kb_valid_14; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1071 = 5'hf == replace_idx | array4kb_valid_15; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1072 = 5'h10 == replace_idx | array4kb_valid_16; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1073 = 5'h11 == replace_idx | array4kb_valid_17; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1074 = 5'h12 == replace_idx | array4kb_valid_18; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1075 = 5'h13 == replace_idx | array4kb_valid_19; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1076 = 5'h14 == replace_idx | array4kb_valid_20; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1077 = 5'h15 == replace_idx | array4kb_valid_21; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1078 = 5'h16 == replace_idx | array4kb_valid_22; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1079 = 5'h17 == replace_idx | array4kb_valid_23; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1080 = 5'h18 == replace_idx | array4kb_valid_24; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1081 = 5'h19 == replace_idx | array4kb_valid_25; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1082 = 5'h1a == replace_idx | array4kb_valid_26; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1083 = 5'h1b == replace_idx | array4kb_valid_27; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1084 = 5'h1c == replace_idx | array4kb_valid_28; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1085 = 5'h1d == replace_idx | array4kb_valid_29; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1086 = 5'h1e == replace_idx | array4kb_valid_30; // @[TLB.scala 65:31 87:{33,33}]
  wire  _GEN_1087 = 5'h1f == replace_idx | array4kb_valid_31; // @[TLB.scala 65:31 87:{33,33}]
  reg  array2mb_0_flag_d; // @[TLB.scala 98:31]
  reg  array2mb_0_flag_a; // @[TLB.scala 98:31]
  reg  array2mb_0_flag_g; // @[TLB.scala 98:31]
  reg  array2mb_0_flag_u; // @[TLB.scala 98:31]
  reg  array2mb_0_flag_x; // @[TLB.scala 98:31]
  reg  array2mb_0_flag_w; // @[TLB.scala 98:31]
  reg  array2mb_0_flag_r; // @[TLB.scala 98:31]
  reg  array2mb_0_flag_v; // @[TLB.scala 98:31]
  reg [8:0] array2mb_0_vpn2; // @[TLB.scala 98:31]
  reg [8:0] array2mb_0_vpn1; // @[TLB.scala 98:31]
  reg [1:0] array2mb_0_ppn2; // @[TLB.scala 98:31]
  reg [8:0] array2mb_0_ppn1; // @[TLB.scala 98:31]
  reg [15:0] array2mb_0_asid; // @[TLB.scala 98:31]
  reg  array2mb_1_flag_d; // @[TLB.scala 98:31]
  reg  array2mb_1_flag_a; // @[TLB.scala 98:31]
  reg  array2mb_1_flag_g; // @[TLB.scala 98:31]
  reg  array2mb_1_flag_u; // @[TLB.scala 98:31]
  reg  array2mb_1_flag_x; // @[TLB.scala 98:31]
  reg  array2mb_1_flag_w; // @[TLB.scala 98:31]
  reg  array2mb_1_flag_r; // @[TLB.scala 98:31]
  reg  array2mb_1_flag_v; // @[TLB.scala 98:31]
  reg [8:0] array2mb_1_vpn2; // @[TLB.scala 98:31]
  reg [8:0] array2mb_1_vpn1; // @[TLB.scala 98:31]
  reg [1:0] array2mb_1_ppn2; // @[TLB.scala 98:31]
  reg [8:0] array2mb_1_ppn1; // @[TLB.scala 98:31]
  reg [15:0] array2mb_1_asid; // @[TLB.scala 98:31]
  reg  array2mb_2_flag_d; // @[TLB.scala 98:31]
  reg  array2mb_2_flag_a; // @[TLB.scala 98:31]
  reg  array2mb_2_flag_g; // @[TLB.scala 98:31]
  reg  array2mb_2_flag_u; // @[TLB.scala 98:31]
  reg  array2mb_2_flag_x; // @[TLB.scala 98:31]
  reg  array2mb_2_flag_w; // @[TLB.scala 98:31]
  reg  array2mb_2_flag_r; // @[TLB.scala 98:31]
  reg  array2mb_2_flag_v; // @[TLB.scala 98:31]
  reg [8:0] array2mb_2_vpn2; // @[TLB.scala 98:31]
  reg [8:0] array2mb_2_vpn1; // @[TLB.scala 98:31]
  reg [1:0] array2mb_2_ppn2; // @[TLB.scala 98:31]
  reg [8:0] array2mb_2_ppn1; // @[TLB.scala 98:31]
  reg [15:0] array2mb_2_asid; // @[TLB.scala 98:31]
  reg  array2mb_3_flag_d; // @[TLB.scala 98:31]
  reg  array2mb_3_flag_a; // @[TLB.scala 98:31]
  reg  array2mb_3_flag_g; // @[TLB.scala 98:31]
  reg  array2mb_3_flag_u; // @[TLB.scala 98:31]
  reg  array2mb_3_flag_x; // @[TLB.scala 98:31]
  reg  array2mb_3_flag_w; // @[TLB.scala 98:31]
  reg  array2mb_3_flag_r; // @[TLB.scala 98:31]
  reg  array2mb_3_flag_v; // @[TLB.scala 98:31]
  reg [8:0] array2mb_3_vpn2; // @[TLB.scala 98:31]
  reg [8:0] array2mb_3_vpn1; // @[TLB.scala 98:31]
  reg [1:0] array2mb_3_ppn2; // @[TLB.scala 98:31]
  reg [8:0] array2mb_3_ppn1; // @[TLB.scala 98:31]
  reg [15:0] array2mb_3_asid; // @[TLB.scala 98:31]
  reg  array2mb_4_flag_d; // @[TLB.scala 98:31]
  reg  array2mb_4_flag_a; // @[TLB.scala 98:31]
  reg  array2mb_4_flag_g; // @[TLB.scala 98:31]
  reg  array2mb_4_flag_u; // @[TLB.scala 98:31]
  reg  array2mb_4_flag_x; // @[TLB.scala 98:31]
  reg  array2mb_4_flag_w; // @[TLB.scala 98:31]
  reg  array2mb_4_flag_r; // @[TLB.scala 98:31]
  reg  array2mb_4_flag_v; // @[TLB.scala 98:31]
  reg [8:0] array2mb_4_vpn2; // @[TLB.scala 98:31]
  reg [8:0] array2mb_4_vpn1; // @[TLB.scala 98:31]
  reg [1:0] array2mb_4_ppn2; // @[TLB.scala 98:31]
  reg [8:0] array2mb_4_ppn1; // @[TLB.scala 98:31]
  reg [15:0] array2mb_4_asid; // @[TLB.scala 98:31]
  reg  array2mb_5_flag_d; // @[TLB.scala 98:31]
  reg  array2mb_5_flag_a; // @[TLB.scala 98:31]
  reg  array2mb_5_flag_g; // @[TLB.scala 98:31]
  reg  array2mb_5_flag_u; // @[TLB.scala 98:31]
  reg  array2mb_5_flag_x; // @[TLB.scala 98:31]
  reg  array2mb_5_flag_w; // @[TLB.scala 98:31]
  reg  array2mb_5_flag_r; // @[TLB.scala 98:31]
  reg  array2mb_5_flag_v; // @[TLB.scala 98:31]
  reg [8:0] array2mb_5_vpn2; // @[TLB.scala 98:31]
  reg [8:0] array2mb_5_vpn1; // @[TLB.scala 98:31]
  reg [1:0] array2mb_5_ppn2; // @[TLB.scala 98:31]
  reg [8:0] array2mb_5_ppn1; // @[TLB.scala 98:31]
  reg [15:0] array2mb_5_asid; // @[TLB.scala 98:31]
  reg  array2mb_6_flag_d; // @[TLB.scala 98:31]
  reg  array2mb_6_flag_a; // @[TLB.scala 98:31]
  reg  array2mb_6_flag_g; // @[TLB.scala 98:31]
  reg  array2mb_6_flag_u; // @[TLB.scala 98:31]
  reg  array2mb_6_flag_x; // @[TLB.scala 98:31]
  reg  array2mb_6_flag_w; // @[TLB.scala 98:31]
  reg  array2mb_6_flag_r; // @[TLB.scala 98:31]
  reg  array2mb_6_flag_v; // @[TLB.scala 98:31]
  reg [8:0] array2mb_6_vpn2; // @[TLB.scala 98:31]
  reg [8:0] array2mb_6_vpn1; // @[TLB.scala 98:31]
  reg [1:0] array2mb_6_ppn2; // @[TLB.scala 98:31]
  reg [8:0] array2mb_6_ppn1; // @[TLB.scala 98:31]
  reg [15:0] array2mb_6_asid; // @[TLB.scala 98:31]
  reg  array2mb_7_flag_d; // @[TLB.scala 98:31]
  reg  array2mb_7_flag_a; // @[TLB.scala 98:31]
  reg  array2mb_7_flag_g; // @[TLB.scala 98:31]
  reg  array2mb_7_flag_u; // @[TLB.scala 98:31]
  reg  array2mb_7_flag_x; // @[TLB.scala 98:31]
  reg  array2mb_7_flag_w; // @[TLB.scala 98:31]
  reg  array2mb_7_flag_r; // @[TLB.scala 98:31]
  reg  array2mb_7_flag_v; // @[TLB.scala 98:31]
  reg [8:0] array2mb_7_vpn2; // @[TLB.scala 98:31]
  reg [8:0] array2mb_7_vpn1; // @[TLB.scala 98:31]
  reg [1:0] array2mb_7_ppn2; // @[TLB.scala 98:31]
  reg [8:0] array2mb_7_ppn1; // @[TLB.scala 98:31]
  reg [15:0] array2mb_7_asid; // @[TLB.scala 98:31]
  reg  array2mb_valid_0; // @[TLB.scala 99:31]
  reg  array2mb_valid_1; // @[TLB.scala 99:31]
  reg  array2mb_valid_2; // @[TLB.scala 99:31]
  reg  array2mb_valid_3; // @[TLB.scala 99:31]
  reg  array2mb_valid_4; // @[TLB.scala 99:31]
  reg  array2mb_valid_5; // @[TLB.scala 99:31]
  reg  array2mb_valid_6; // @[TLB.scala 99:31]
  reg  array2mb_valid_7; // @[TLB.scala 99:31]
  wire [17:0] _T_138 = {array2mb_0_vpn2,array2mb_0_vpn1}; // @[Cat.scala 33:92]
  wire  _GEN_1664 = array2mb_valid_0 & _T_138 == hi_1 & (array2mb_0_asid == io_satp_asid | array2mb_0_flag_g); // @[TLB.scala 105:77 106:22 102:35]
  wire  _GEN_1666 = array2mb_valid_0 & _T_138 == hi_1 & array2mb_0_flag_d; // @[TLB.scala 105:77 107:22 100:35]
  wire  _GEN_1667 = array2mb_valid_0 & _T_138 == hi_1 & array2mb_0_flag_a; // @[TLB.scala 105:77 107:22 100:35]
  wire  _GEN_1669 = array2mb_valid_0 & _T_138 == hi_1 & array2mb_0_flag_u; // @[TLB.scala 105:77 107:22 100:35]
  wire  _GEN_1670 = array2mb_valid_0 & _T_138 == hi_1 & array2mb_0_flag_x; // @[TLB.scala 105:77 107:22 100:35]
  wire  _GEN_1671 = array2mb_valid_0 & _T_138 == hi_1 & array2mb_0_flag_w; // @[TLB.scala 105:77 107:22 100:35]
  wire  _GEN_1672 = array2mb_valid_0 & _T_138 == hi_1 & array2mb_0_flag_r; // @[TLB.scala 105:77 107:22 100:35]
  wire  _GEN_1673 = array2mb_valid_0 & _T_138 == hi_1 & array2mb_0_flag_v; // @[TLB.scala 105:77 107:22 100:35]
  wire [1:0] _GEN_1676 = array2mb_valid_0 & _T_138 == hi_1 ? array2mb_0_ppn2 : 2'h0; // @[TLB.scala 105:77 107:22 100:35]
  wire [8:0] _GEN_1677 = array2mb_valid_0 & _T_138 == hi_1 ? array2mb_0_ppn1 : 9'h0; // @[TLB.scala 105:77 107:22 100:35]
  wire [17:0] _T_142 = {array2mb_1_vpn2,array2mb_1_vpn1}; // @[Cat.scala 33:92]
  wire  _GEN_1679 = array2mb_valid_1 & _T_142 == hi_1 ? array2mb_1_asid == io_satp_asid | array2mb_1_flag_g : _GEN_1664; // @[TLB.scala 105:77 106:22]
  wire  _GEN_1681 = array2mb_valid_1 & _T_142 == hi_1 ? array2mb_1_flag_d : _GEN_1666; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1682 = array2mb_valid_1 & _T_142 == hi_1 ? array2mb_1_flag_a : _GEN_1667; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1684 = array2mb_valid_1 & _T_142 == hi_1 ? array2mb_1_flag_u : _GEN_1669; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1685 = array2mb_valid_1 & _T_142 == hi_1 ? array2mb_1_flag_x : _GEN_1670; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1686 = array2mb_valid_1 & _T_142 == hi_1 ? array2mb_1_flag_w : _GEN_1671; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1687 = array2mb_valid_1 & _T_142 == hi_1 ? array2mb_1_flag_r : _GEN_1672; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1688 = array2mb_valid_1 & _T_142 == hi_1 ? array2mb_1_flag_v : _GEN_1673; // @[TLB.scala 105:77 107:22]
  wire [1:0] _GEN_1691 = array2mb_valid_1 & _T_142 == hi_1 ? array2mb_1_ppn2 : _GEN_1676; // @[TLB.scala 105:77 107:22]
  wire [8:0] _GEN_1692 = array2mb_valid_1 & _T_142 == hi_1 ? array2mb_1_ppn1 : _GEN_1677; // @[TLB.scala 105:77 107:22]
  wire [17:0] _T_146 = {array2mb_2_vpn2,array2mb_2_vpn1}; // @[Cat.scala 33:92]
  wire  _GEN_1694 = array2mb_valid_2 & _T_146 == hi_1 ? array2mb_2_asid == io_satp_asid | array2mb_2_flag_g : _GEN_1679; // @[TLB.scala 105:77 106:22]
  wire  _GEN_1696 = array2mb_valid_2 & _T_146 == hi_1 ? array2mb_2_flag_d : _GEN_1681; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1697 = array2mb_valid_2 & _T_146 == hi_1 ? array2mb_2_flag_a : _GEN_1682; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1699 = array2mb_valid_2 & _T_146 == hi_1 ? array2mb_2_flag_u : _GEN_1684; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1700 = array2mb_valid_2 & _T_146 == hi_1 ? array2mb_2_flag_x : _GEN_1685; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1701 = array2mb_valid_2 & _T_146 == hi_1 ? array2mb_2_flag_w : _GEN_1686; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1702 = array2mb_valid_2 & _T_146 == hi_1 ? array2mb_2_flag_r : _GEN_1687; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1703 = array2mb_valid_2 & _T_146 == hi_1 ? array2mb_2_flag_v : _GEN_1688; // @[TLB.scala 105:77 107:22]
  wire [1:0] _GEN_1706 = array2mb_valid_2 & _T_146 == hi_1 ? array2mb_2_ppn2 : _GEN_1691; // @[TLB.scala 105:77 107:22]
  wire [8:0] _GEN_1707 = array2mb_valid_2 & _T_146 == hi_1 ? array2mb_2_ppn1 : _GEN_1692; // @[TLB.scala 105:77 107:22]
  wire [17:0] _T_150 = {array2mb_3_vpn2,array2mb_3_vpn1}; // @[Cat.scala 33:92]
  wire  _GEN_1709 = array2mb_valid_3 & _T_150 == hi_1 ? array2mb_3_asid == io_satp_asid | array2mb_3_flag_g : _GEN_1694; // @[TLB.scala 105:77 106:22]
  wire  _GEN_1711 = array2mb_valid_3 & _T_150 == hi_1 ? array2mb_3_flag_d : _GEN_1696; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1712 = array2mb_valid_3 & _T_150 == hi_1 ? array2mb_3_flag_a : _GEN_1697; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1714 = array2mb_valid_3 & _T_150 == hi_1 ? array2mb_3_flag_u : _GEN_1699; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1715 = array2mb_valid_3 & _T_150 == hi_1 ? array2mb_3_flag_x : _GEN_1700; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1716 = array2mb_valid_3 & _T_150 == hi_1 ? array2mb_3_flag_w : _GEN_1701; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1717 = array2mb_valid_3 & _T_150 == hi_1 ? array2mb_3_flag_r : _GEN_1702; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1718 = array2mb_valid_3 & _T_150 == hi_1 ? array2mb_3_flag_v : _GEN_1703; // @[TLB.scala 105:77 107:22]
  wire [1:0] _GEN_1721 = array2mb_valid_3 & _T_150 == hi_1 ? array2mb_3_ppn2 : _GEN_1706; // @[TLB.scala 105:77 107:22]
  wire [8:0] _GEN_1722 = array2mb_valid_3 & _T_150 == hi_1 ? array2mb_3_ppn1 : _GEN_1707; // @[TLB.scala 105:77 107:22]
  wire [17:0] _T_154 = {array2mb_4_vpn2,array2mb_4_vpn1}; // @[Cat.scala 33:92]
  wire  _GEN_1724 = array2mb_valid_4 & _T_154 == hi_1 ? array2mb_4_asid == io_satp_asid | array2mb_4_flag_g : _GEN_1709; // @[TLB.scala 105:77 106:22]
  wire  _GEN_1726 = array2mb_valid_4 & _T_154 == hi_1 ? array2mb_4_flag_d : _GEN_1711; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1727 = array2mb_valid_4 & _T_154 == hi_1 ? array2mb_4_flag_a : _GEN_1712; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1729 = array2mb_valid_4 & _T_154 == hi_1 ? array2mb_4_flag_u : _GEN_1714; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1730 = array2mb_valid_4 & _T_154 == hi_1 ? array2mb_4_flag_x : _GEN_1715; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1731 = array2mb_valid_4 & _T_154 == hi_1 ? array2mb_4_flag_w : _GEN_1716; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1732 = array2mb_valid_4 & _T_154 == hi_1 ? array2mb_4_flag_r : _GEN_1717; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1733 = array2mb_valid_4 & _T_154 == hi_1 ? array2mb_4_flag_v : _GEN_1718; // @[TLB.scala 105:77 107:22]
  wire [1:0] _GEN_1736 = array2mb_valid_4 & _T_154 == hi_1 ? array2mb_4_ppn2 : _GEN_1721; // @[TLB.scala 105:77 107:22]
  wire [8:0] _GEN_1737 = array2mb_valid_4 & _T_154 == hi_1 ? array2mb_4_ppn1 : _GEN_1722; // @[TLB.scala 105:77 107:22]
  wire [17:0] _T_158 = {array2mb_5_vpn2,array2mb_5_vpn1}; // @[Cat.scala 33:92]
  wire  _GEN_1739 = array2mb_valid_5 & _T_158 == hi_1 ? array2mb_5_asid == io_satp_asid | array2mb_5_flag_g : _GEN_1724; // @[TLB.scala 105:77 106:22]
  wire  _GEN_1741 = array2mb_valid_5 & _T_158 == hi_1 ? array2mb_5_flag_d : _GEN_1726; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1742 = array2mb_valid_5 & _T_158 == hi_1 ? array2mb_5_flag_a : _GEN_1727; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1744 = array2mb_valid_5 & _T_158 == hi_1 ? array2mb_5_flag_u : _GEN_1729; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1745 = array2mb_valid_5 & _T_158 == hi_1 ? array2mb_5_flag_x : _GEN_1730; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1746 = array2mb_valid_5 & _T_158 == hi_1 ? array2mb_5_flag_w : _GEN_1731; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1747 = array2mb_valid_5 & _T_158 == hi_1 ? array2mb_5_flag_r : _GEN_1732; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1748 = array2mb_valid_5 & _T_158 == hi_1 ? array2mb_5_flag_v : _GEN_1733; // @[TLB.scala 105:77 107:22]
  wire [1:0] _GEN_1751 = array2mb_valid_5 & _T_158 == hi_1 ? array2mb_5_ppn2 : _GEN_1736; // @[TLB.scala 105:77 107:22]
  wire [8:0] _GEN_1752 = array2mb_valid_5 & _T_158 == hi_1 ? array2mb_5_ppn1 : _GEN_1737; // @[TLB.scala 105:77 107:22]
  wire [17:0] _T_162 = {array2mb_6_vpn2,array2mb_6_vpn1}; // @[Cat.scala 33:92]
  wire  _GEN_1754 = array2mb_valid_6 & _T_162 == hi_1 ? array2mb_6_asid == io_satp_asid | array2mb_6_flag_g : _GEN_1739; // @[TLB.scala 105:77 106:22]
  wire  _GEN_1756 = array2mb_valid_6 & _T_162 == hi_1 ? array2mb_6_flag_d : _GEN_1741; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1757 = array2mb_valid_6 & _T_162 == hi_1 ? array2mb_6_flag_a : _GEN_1742; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1759 = array2mb_valid_6 & _T_162 == hi_1 ? array2mb_6_flag_u : _GEN_1744; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1760 = array2mb_valid_6 & _T_162 == hi_1 ? array2mb_6_flag_x : _GEN_1745; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1761 = array2mb_valid_6 & _T_162 == hi_1 ? array2mb_6_flag_w : _GEN_1746; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1762 = array2mb_valid_6 & _T_162 == hi_1 ? array2mb_6_flag_r : _GEN_1747; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1763 = array2mb_valid_6 & _T_162 == hi_1 ? array2mb_6_flag_v : _GEN_1748; // @[TLB.scala 105:77 107:22]
  wire [1:0] _GEN_1766 = array2mb_valid_6 & _T_162 == hi_1 ? array2mb_6_ppn2 : _GEN_1751; // @[TLB.scala 105:77 107:22]
  wire [8:0] _GEN_1767 = array2mb_valid_6 & _T_162 == hi_1 ? array2mb_6_ppn1 : _GEN_1752; // @[TLB.scala 105:77 107:22]
  wire [17:0] _T_166 = {array2mb_7_vpn2,array2mb_7_vpn1}; // @[Cat.scala 33:92]
  wire  hit2mb = array2mb_valid_7 & _T_166 == hi_1 ? array2mb_7_asid == io_satp_asid | array2mb_7_flag_g : _GEN_1754; // @[TLB.scala 105:77 106:22]
  wire  array2mb_rdata_flag_d = array2mb_valid_7 & _T_166 == hi_1 ? array2mb_7_flag_d : _GEN_1756; // @[TLB.scala 105:77 107:22]
  wire  array2mb_rdata_flag_a = array2mb_valid_7 & _T_166 == hi_1 ? array2mb_7_flag_a : _GEN_1757; // @[TLB.scala 105:77 107:22]
  wire  array2mb_rdata_flag_u = array2mb_valid_7 & _T_166 == hi_1 ? array2mb_7_flag_u : _GEN_1759; // @[TLB.scala 105:77 107:22]
  wire  array2mb_rdata_flag_x = array2mb_valid_7 & _T_166 == hi_1 ? array2mb_7_flag_x : _GEN_1760; // @[TLB.scala 105:77 107:22]
  wire  array2mb_rdata_flag_w = array2mb_valid_7 & _T_166 == hi_1 ? array2mb_7_flag_w : _GEN_1761; // @[TLB.scala 105:77 107:22]
  wire  array2mb_rdata_flag_r = array2mb_valid_7 & _T_166 == hi_1 ? array2mb_7_flag_r : _GEN_1762; // @[TLB.scala 105:77 107:22]
  wire  array2mb_rdata_flag_v = array2mb_valid_7 & _T_166 == hi_1 ? array2mb_7_flag_v : _GEN_1763; // @[TLB.scala 105:77 107:22]
  wire [1:0] array2mb_rdata_ppn2 = array2mb_valid_7 & _T_166 == hi_1 ? array2mb_7_ppn2 : _GEN_1766; // @[TLB.scala 105:77 107:22]
  wire [8:0] array2mb_rdata_ppn1 = array2mb_valid_7 & _T_166 == hi_1 ? array2mb_7_ppn1 : _GEN_1767; // @[TLB.scala 105:77 107:22]
  wire  _GEN_1896 = 3'h0 == replace_idx[2:0] | array2mb_valid_0; // @[TLB.scala 119:{33,33} 99:31]
  wire  _GEN_1897 = 3'h1 == replace_idx[2:0] | array2mb_valid_1; // @[TLB.scala 119:{33,33} 99:31]
  wire  _GEN_1898 = 3'h2 == replace_idx[2:0] | array2mb_valid_2; // @[TLB.scala 119:{33,33} 99:31]
  wire  _GEN_1899 = 3'h3 == replace_idx[2:0] | array2mb_valid_3; // @[TLB.scala 119:{33,33} 99:31]
  wire  _GEN_1900 = 3'h4 == replace_idx[2:0] | array2mb_valid_4; // @[TLB.scala 119:{33,33} 99:31]
  wire  _GEN_1901 = 3'h5 == replace_idx[2:0] | array2mb_valid_5; // @[TLB.scala 119:{33,33} 99:31]
  wire  _GEN_1902 = 3'h6 == replace_idx[2:0] | array2mb_valid_6; // @[TLB.scala 119:{33,33} 99:31]
  wire  _GEN_1903 = 3'h7 == replace_idx[2:0] | array2mb_valid_7; // @[TLB.scala 119:{33,33} 99:31]
  reg  array1gb_0_flag_d; // @[TLB.scala 130:31]
  reg  array1gb_0_flag_a; // @[TLB.scala 130:31]
  reg  array1gb_0_flag_g; // @[TLB.scala 130:31]
  reg  array1gb_0_flag_u; // @[TLB.scala 130:31]
  reg  array1gb_0_flag_x; // @[TLB.scala 130:31]
  reg  array1gb_0_flag_w; // @[TLB.scala 130:31]
  reg  array1gb_0_flag_r; // @[TLB.scala 130:31]
  reg  array1gb_0_flag_v; // @[TLB.scala 130:31]
  reg [8:0] array1gb_0_vpn2; // @[TLB.scala 130:31]
  reg [1:0] array1gb_0_ppn2; // @[TLB.scala 130:31]
  reg [15:0] array1gb_0_asid; // @[TLB.scala 130:31]
  reg  array1gb_1_flag_d; // @[TLB.scala 130:31]
  reg  array1gb_1_flag_a; // @[TLB.scala 130:31]
  reg  array1gb_1_flag_g; // @[TLB.scala 130:31]
  reg  array1gb_1_flag_u; // @[TLB.scala 130:31]
  reg  array1gb_1_flag_x; // @[TLB.scala 130:31]
  reg  array1gb_1_flag_w; // @[TLB.scala 130:31]
  reg  array1gb_1_flag_r; // @[TLB.scala 130:31]
  reg  array1gb_1_flag_v; // @[TLB.scala 130:31]
  reg [8:0] array1gb_1_vpn2; // @[TLB.scala 130:31]
  reg [1:0] array1gb_1_ppn2; // @[TLB.scala 130:31]
  reg [15:0] array1gb_1_asid; // @[TLB.scala 130:31]
  reg  array1gb_2_flag_d; // @[TLB.scala 130:31]
  reg  array1gb_2_flag_a; // @[TLB.scala 130:31]
  reg  array1gb_2_flag_g; // @[TLB.scala 130:31]
  reg  array1gb_2_flag_u; // @[TLB.scala 130:31]
  reg  array1gb_2_flag_x; // @[TLB.scala 130:31]
  reg  array1gb_2_flag_w; // @[TLB.scala 130:31]
  reg  array1gb_2_flag_r; // @[TLB.scala 130:31]
  reg  array1gb_2_flag_v; // @[TLB.scala 130:31]
  reg [8:0] array1gb_2_vpn2; // @[TLB.scala 130:31]
  reg [1:0] array1gb_2_ppn2; // @[TLB.scala 130:31]
  reg [15:0] array1gb_2_asid; // @[TLB.scala 130:31]
  reg  array1gb_3_flag_d; // @[TLB.scala 130:31]
  reg  array1gb_3_flag_a; // @[TLB.scala 130:31]
  reg  array1gb_3_flag_g; // @[TLB.scala 130:31]
  reg  array1gb_3_flag_u; // @[TLB.scala 130:31]
  reg  array1gb_3_flag_x; // @[TLB.scala 130:31]
  reg  array1gb_3_flag_w; // @[TLB.scala 130:31]
  reg  array1gb_3_flag_r; // @[TLB.scala 130:31]
  reg  array1gb_3_flag_v; // @[TLB.scala 130:31]
  reg [8:0] array1gb_3_vpn2; // @[TLB.scala 130:31]
  reg [1:0] array1gb_3_ppn2; // @[TLB.scala 130:31]
  reg [15:0] array1gb_3_asid; // @[TLB.scala 130:31]
  reg  array1gb_valid_0; // @[TLB.scala 131:31]
  reg  array1gb_valid_1; // @[TLB.scala 131:31]
  reg  array1gb_valid_2; // @[TLB.scala 131:31]
  reg  array1gb_valid_3; // @[TLB.scala 131:31]
  wire  _GEN_2032 = array1gb_valid_0 & array1gb_0_vpn2 == io_vaddr_vpn2 & (array1gb_0_asid == io_satp_asid |
    array1gb_0_flag_g); // @[TLB.scala 137:77 138:22 134:35]
  wire  _GEN_2034 = array1gb_valid_0 & array1gb_0_vpn2 == io_vaddr_vpn2 & array1gb_0_flag_d; // @[TLB.scala 137:77 139:22 132:35]
  wire  _GEN_2035 = array1gb_valid_0 & array1gb_0_vpn2 == io_vaddr_vpn2 & array1gb_0_flag_a; // @[TLB.scala 137:77 139:22 132:35]
  wire  _GEN_2037 = array1gb_valid_0 & array1gb_0_vpn2 == io_vaddr_vpn2 & array1gb_0_flag_u; // @[TLB.scala 137:77 139:22 132:35]
  wire  _GEN_2038 = array1gb_valid_0 & array1gb_0_vpn2 == io_vaddr_vpn2 & array1gb_0_flag_x; // @[TLB.scala 137:77 139:22 132:35]
  wire  _GEN_2039 = array1gb_valid_0 & array1gb_0_vpn2 == io_vaddr_vpn2 & array1gb_0_flag_w; // @[TLB.scala 137:77 139:22 132:35]
  wire  _GEN_2040 = array1gb_valid_0 & array1gb_0_vpn2 == io_vaddr_vpn2 & array1gb_0_flag_r; // @[TLB.scala 137:77 139:22 132:35]
  wire  _GEN_2041 = array1gb_valid_0 & array1gb_0_vpn2 == io_vaddr_vpn2 & array1gb_0_flag_v; // @[TLB.scala 137:77 139:22 132:35]
  wire [1:0] _GEN_2043 = array1gb_valid_0 & array1gb_0_vpn2 == io_vaddr_vpn2 ? array1gb_0_ppn2 : 2'h0; // @[TLB.scala 137:77 139:22 132:35]
  wire  _GEN_2045 = array1gb_valid_1 & array1gb_1_vpn2 == io_vaddr_vpn2 ? array1gb_1_asid == io_satp_asid |
    array1gb_1_flag_g : _GEN_2032; // @[TLB.scala 137:77 138:22]
  wire  _GEN_2047 = array1gb_valid_1 & array1gb_1_vpn2 == io_vaddr_vpn2 ? array1gb_1_flag_d : _GEN_2034; // @[TLB.scala 137:77 139:22]
  wire  _GEN_2048 = array1gb_valid_1 & array1gb_1_vpn2 == io_vaddr_vpn2 ? array1gb_1_flag_a : _GEN_2035; // @[TLB.scala 137:77 139:22]
  wire  _GEN_2050 = array1gb_valid_1 & array1gb_1_vpn2 == io_vaddr_vpn2 ? array1gb_1_flag_u : _GEN_2037; // @[TLB.scala 137:77 139:22]
  wire  _GEN_2051 = array1gb_valid_1 & array1gb_1_vpn2 == io_vaddr_vpn2 ? array1gb_1_flag_x : _GEN_2038; // @[TLB.scala 137:77 139:22]
  wire  _GEN_2052 = array1gb_valid_1 & array1gb_1_vpn2 == io_vaddr_vpn2 ? array1gb_1_flag_w : _GEN_2039; // @[TLB.scala 137:77 139:22]
  wire  _GEN_2053 = array1gb_valid_1 & array1gb_1_vpn2 == io_vaddr_vpn2 ? array1gb_1_flag_r : _GEN_2040; // @[TLB.scala 137:77 139:22]
  wire  _GEN_2054 = array1gb_valid_1 & array1gb_1_vpn2 == io_vaddr_vpn2 ? array1gb_1_flag_v : _GEN_2041; // @[TLB.scala 137:77 139:22]
  wire [1:0] _GEN_2056 = array1gb_valid_1 & array1gb_1_vpn2 == io_vaddr_vpn2 ? array1gb_1_ppn2 : _GEN_2043; // @[TLB.scala 137:77 139:22]
  wire  _GEN_2058 = array1gb_valid_2 & array1gb_2_vpn2 == io_vaddr_vpn2 ? array1gb_2_asid == io_satp_asid |
    array1gb_2_flag_g : _GEN_2045; // @[TLB.scala 137:77 138:22]
  wire  _GEN_2060 = array1gb_valid_2 & array1gb_2_vpn2 == io_vaddr_vpn2 ? array1gb_2_flag_d : _GEN_2047; // @[TLB.scala 137:77 139:22]
  wire  _GEN_2061 = array1gb_valid_2 & array1gb_2_vpn2 == io_vaddr_vpn2 ? array1gb_2_flag_a : _GEN_2048; // @[TLB.scala 137:77 139:22]
  wire  _GEN_2063 = array1gb_valid_2 & array1gb_2_vpn2 == io_vaddr_vpn2 ? array1gb_2_flag_u : _GEN_2050; // @[TLB.scala 137:77 139:22]
  wire  _GEN_2064 = array1gb_valid_2 & array1gb_2_vpn2 == io_vaddr_vpn2 ? array1gb_2_flag_x : _GEN_2051; // @[TLB.scala 137:77 139:22]
  wire  _GEN_2065 = array1gb_valid_2 & array1gb_2_vpn2 == io_vaddr_vpn2 ? array1gb_2_flag_w : _GEN_2052; // @[TLB.scala 137:77 139:22]
  wire  _GEN_2066 = array1gb_valid_2 & array1gb_2_vpn2 == io_vaddr_vpn2 ? array1gb_2_flag_r : _GEN_2053; // @[TLB.scala 137:77 139:22]
  wire  _GEN_2067 = array1gb_valid_2 & array1gb_2_vpn2 == io_vaddr_vpn2 ? array1gb_2_flag_v : _GEN_2054; // @[TLB.scala 137:77 139:22]
  wire [1:0] _GEN_2069 = array1gb_valid_2 & array1gb_2_vpn2 == io_vaddr_vpn2 ? array1gb_2_ppn2 : _GEN_2056; // @[TLB.scala 137:77 139:22]
  wire  hit1gb = array1gb_valid_3 & array1gb_3_vpn2 == io_vaddr_vpn2 ? array1gb_3_asid == io_satp_asid |
    array1gb_3_flag_g : _GEN_2058; // @[TLB.scala 137:77 138:22]
  wire  array1gb_rdata_flag_d = array1gb_valid_3 & array1gb_3_vpn2 == io_vaddr_vpn2 ? array1gb_3_flag_d : _GEN_2060; // @[TLB.scala 137:77 139:22]
  wire  array1gb_rdata_flag_a = array1gb_valid_3 & array1gb_3_vpn2 == io_vaddr_vpn2 ? array1gb_3_flag_a : _GEN_2061; // @[TLB.scala 137:77 139:22]
  wire  array1gb_rdata_flag_u = array1gb_valid_3 & array1gb_3_vpn2 == io_vaddr_vpn2 ? array1gb_3_flag_u : _GEN_2063; // @[TLB.scala 137:77 139:22]
  wire  array1gb_rdata_flag_x = array1gb_valid_3 & array1gb_3_vpn2 == io_vaddr_vpn2 ? array1gb_3_flag_x : _GEN_2064; // @[TLB.scala 137:77 139:22]
  wire  array1gb_rdata_flag_w = array1gb_valid_3 & array1gb_3_vpn2 == io_vaddr_vpn2 ? array1gb_3_flag_w : _GEN_2065; // @[TLB.scala 137:77 139:22]
  wire  array1gb_rdata_flag_r = array1gb_valid_3 & array1gb_3_vpn2 == io_vaddr_vpn2 ? array1gb_3_flag_r : _GEN_2066; // @[TLB.scala 137:77 139:22]
  wire  array1gb_rdata_flag_v = array1gb_valid_3 & array1gb_3_vpn2 == io_vaddr_vpn2 ? array1gb_3_flag_v : _GEN_2067; // @[TLB.scala 137:77 139:22]
  wire [1:0] array1gb_rdata_ppn2 = array1gb_valid_3 & array1gb_3_vpn2 == io_vaddr_vpn2 ? array1gb_3_ppn2 : _GEN_2069; // @[TLB.scala 137:77 139:22]
  wire  _GEN_2132 = 2'h0 == replace_idx[1:0] | array1gb_valid_0; // @[TLB.scala 131:31 149:{33,33}]
  wire  _GEN_2133 = 2'h1 == replace_idx[1:0] | array1gb_valid_1; // @[TLB.scala 131:31 149:{33,33}]
  wire  _GEN_2134 = 2'h2 == replace_idx[1:0] | array1gb_valid_2; // @[TLB.scala 131:31 149:{33,33}]
  wire  _GEN_2135 = 2'h3 == replace_idx[1:0] | array1gb_valid_3; // @[TLB.scala 131:31 149:{33,33}]
  wire  _GEN_2193 = hit1gb & array1gb_rdata_flag_d; // @[TLB.scala 158:13 172:22 173:18]
  wire  _GEN_2194 = hit1gb & array1gb_rdata_flag_a; // @[TLB.scala 158:13 172:22 173:18]
  wire  _GEN_2196 = hit1gb & array1gb_rdata_flag_u; // @[TLB.scala 158:13 172:22 173:18]
  wire  _GEN_2197 = hit1gb & array1gb_rdata_flag_x; // @[TLB.scala 158:13 172:22 173:18]
  wire  _GEN_2198 = hit1gb & array1gb_rdata_flag_w; // @[TLB.scala 158:13 172:22 173:18]
  wire  _GEN_2199 = hit1gb & array1gb_rdata_flag_r; // @[TLB.scala 158:13 172:22 173:18]
  wire  _GEN_2200 = hit1gb & array1gb_rdata_flag_v; // @[TLB.scala 158:13 172:22 173:18]
  wire [1:0] _GEN_2203 = hit1gb ? array1gb_rdata_ppn2 : 2'h0; // @[TLB.scala 158:13 172:22 176:18]
  wire [1:0] _GEN_2204 = hit1gb ? 2'h2 : 2'h0; // @[TLB.scala 159:13 172:22 177:18]
  wire  _GEN_2206 = hit2mb ? array2mb_rdata_flag_d : _GEN_2193; // @[TLB.scala 166:22 167:18]
  wire  _GEN_2207 = hit2mb ? array2mb_rdata_flag_a : _GEN_2194; // @[TLB.scala 166:22 167:18]
  wire  _GEN_2209 = hit2mb ? array2mb_rdata_flag_u : _GEN_2196; // @[TLB.scala 166:22 167:18]
  wire  _GEN_2210 = hit2mb ? array2mb_rdata_flag_x : _GEN_2197; // @[TLB.scala 166:22 167:18]
  wire  _GEN_2211 = hit2mb ? array2mb_rdata_flag_w : _GEN_2198; // @[TLB.scala 166:22 167:18]
  wire  _GEN_2212 = hit2mb ? array2mb_rdata_flag_r : _GEN_2199; // @[TLB.scala 166:22 167:18]
  wire  _GEN_2213 = hit2mb ? array2mb_rdata_flag_v : _GEN_2200; // @[TLB.scala 166:22 167:18]
  wire [8:0] _GEN_2215 = hit2mb ? array2mb_rdata_ppn1 : 9'h0; // @[TLB.scala 166:22 169:18]
  wire [1:0] _GEN_2216 = hit2mb ? array2mb_rdata_ppn2 : _GEN_2203; // @[TLB.scala 166:22 170:18]
  wire [1:0] _GEN_2217 = hit2mb ? 2'h1 : _GEN_2204; // @[TLB.scala 166:22 171:18]
  MaxPeriodFibonacciLFSR_1 replace_idx_prng ( // @[PRNG.scala 91:22]
    .clock(replace_idx_prng_clock),
    .reset(replace_idx_prng_reset),
    .io_out_0(replace_idx_prng_io_out_0),
    .io_out_1(replace_idx_prng_io_out_1),
    .io_out_2(replace_idx_prng_io_out_2),
    .io_out_3(replace_idx_prng_io_out_3),
    .io_out_4(replace_idx_prng_io_out_4)
  );
  assign io_rpte_ppn2 = hit4kb ? array4kb_rdata_ppn2 : _GEN_2216; // @[TLB.scala 161:16 165:18]
  assign io_rpte_ppn1 = hit4kb ? array4kb_rdata_ppn1 : _GEN_2215; // @[TLB.scala 161:16 164:18]
  assign io_rpte_ppn0 = hit4kb ? array4kb_rdata_ppn0 : 9'h0; // @[TLB.scala 161:16 163:18]
  assign io_rpte_flag_d = hit4kb ? array4kb_rdata_flag_d : _GEN_2206; // @[TLB.scala 161:16 162:18]
  assign io_rpte_flag_a = hit4kb ? array4kb_rdata_flag_a : _GEN_2207; // @[TLB.scala 161:16 162:18]
  assign io_rpte_flag_u = hit4kb ? array4kb_rdata_flag_u : _GEN_2209; // @[TLB.scala 161:16 162:18]
  assign io_rpte_flag_x = hit4kb ? array4kb_rdata_flag_x : _GEN_2210; // @[TLB.scala 161:16 162:18]
  assign io_rpte_flag_w = hit4kb ? array4kb_rdata_flag_w : _GEN_2211; // @[TLB.scala 161:16 162:18]
  assign io_rpte_flag_r = hit4kb ? array4kb_rdata_flag_r : _GEN_2212; // @[TLB.scala 161:16 162:18]
  assign io_rpte_flag_v = hit4kb ? array4kb_rdata_flag_v : _GEN_2213; // @[TLB.scala 161:16 162:18]
  assign io_rlevel = hit4kb ? 2'h0 : _GEN_2217; // @[TLB.scala 159:13 161:16]
  assign io_hit = hit4kb | hit2mb | hit1gb; // @[TLB.scala 160:33]
  assign replace_idx_prng_clock = clock;
  assign replace_idx_prng_reset = reset;
  always @(posedge clock) begin
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_0_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h0 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_0_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_0_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h0 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_0_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_0_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h0 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_0_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_0_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h0 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_0_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_0_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h0 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_0_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_0_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h0 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_0_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_0_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h0 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_0_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_0_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h0 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_0_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_0_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h0 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_0_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_0_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h0 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_0_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_0_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h0 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_0_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_0_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h0 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_0_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_0_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h0 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_0_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_0_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h0 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_0_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_0_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h0 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_0_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_1_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_1_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_1_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_1_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_1_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_1_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_1_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_1_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_1_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_1_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_1_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_1_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_1_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_1_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_1_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_1_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_1_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_1_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_1_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_1_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_1_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_1_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_1_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_1_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_1_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_1_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_1_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_1_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_1_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_1_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_2_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h2 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_2_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_2_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h2 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_2_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_2_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h2 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_2_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_2_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h2 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_2_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_2_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h2 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_2_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_2_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h2 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_2_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_2_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h2 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_2_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_2_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h2 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_2_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_2_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h2 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_2_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_2_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h2 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_2_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_2_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h2 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_2_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_2_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h2 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_2_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_2_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h2 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_2_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_2_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h2 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_2_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_2_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h2 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_2_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_3_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h3 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_3_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_3_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h3 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_3_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_3_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h3 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_3_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_3_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h3 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_3_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_3_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h3 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_3_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_3_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h3 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_3_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_3_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h3 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_3_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_3_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h3 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_3_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_3_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h3 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_3_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_3_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h3 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_3_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_3_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h3 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_3_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_3_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h3 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_3_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_3_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h3 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_3_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_3_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h3 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_3_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_3_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h3 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_3_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_4_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h4 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_4_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_4_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h4 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_4_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_4_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h4 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_4_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_4_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h4 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_4_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_4_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h4 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_4_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_4_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h4 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_4_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_4_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h4 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_4_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_4_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h4 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_4_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_4_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h4 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_4_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_4_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h4 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_4_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_4_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h4 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_4_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_4_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h4 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_4_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_4_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h4 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_4_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_4_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h4 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_4_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_4_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h4 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_4_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_5_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h5 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_5_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_5_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h5 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_5_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_5_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h5 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_5_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_5_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h5 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_5_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_5_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h5 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_5_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_5_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h5 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_5_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_5_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h5 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_5_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_5_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h5 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_5_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_5_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h5 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_5_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_5_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h5 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_5_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_5_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h5 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_5_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_5_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h5 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_5_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_5_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h5 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_5_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_5_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h5 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_5_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_5_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h5 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_5_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_6_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h6 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_6_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_6_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h6 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_6_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_6_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h6 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_6_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_6_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h6 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_6_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_6_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h6 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_6_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_6_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h6 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_6_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_6_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h6 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_6_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_6_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h6 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_6_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_6_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h6 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_6_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_6_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h6 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_6_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_6_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h6 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_6_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_6_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h6 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_6_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_6_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h6 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_6_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_6_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h6 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_6_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_6_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h6 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_6_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_7_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h7 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_7_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_7_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h7 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_7_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_7_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h7 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_7_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_7_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h7 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_7_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_7_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h7 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_7_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_7_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h7 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_7_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_7_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h7 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_7_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_7_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h7 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_7_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_7_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h7 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_7_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_7_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h7 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_7_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_7_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h7 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_7_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_7_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h7 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_7_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_7_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h7 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_7_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_7_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h7 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_7_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_7_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h7 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_7_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_8_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h8 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_8_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_8_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h8 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_8_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_8_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h8 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_8_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_8_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h8 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_8_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_8_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h8 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_8_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_8_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h8 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_8_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_8_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h8 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_8_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_8_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h8 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_8_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_8_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h8 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_8_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_8_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h8 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_8_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_8_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h8 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_8_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_8_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h8 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_8_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_8_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h8 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_8_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_8_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h8 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_8_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_8_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h8 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_8_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_9_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h9 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_9_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_9_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h9 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_9_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_9_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h9 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_9_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_9_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h9 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_9_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_9_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h9 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_9_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_9_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h9 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_9_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_9_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h9 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_9_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_9_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h9 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_9_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_9_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h9 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_9_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_9_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h9 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_9_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_9_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h9 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_9_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_9_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h9 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_9_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_9_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h9 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_9_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_9_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h9 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_9_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_9_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h9 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_9_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_10_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'ha == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_10_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_10_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'ha == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_10_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_10_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'ha == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_10_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_10_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'ha == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_10_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_10_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'ha == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_10_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_10_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'ha == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_10_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_10_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'ha == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_10_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_10_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'ha == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_10_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_10_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'ha == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_10_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_10_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'ha == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_10_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_10_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'ha == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_10_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_10_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'ha == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_10_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_10_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'ha == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_10_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_10_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'ha == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_10_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_10_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'ha == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_10_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_11_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hb == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_11_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_11_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hb == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_11_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_11_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hb == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_11_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_11_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hb == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_11_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_11_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hb == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_11_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_11_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hb == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_11_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_11_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hb == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_11_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_11_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hb == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_11_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_11_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hb == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_11_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_11_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hb == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_11_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_11_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hb == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_11_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_11_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hb == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_11_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_11_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hb == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_11_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_11_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hb == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_11_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_11_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hb == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_11_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_12_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hc == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_12_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_12_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hc == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_12_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_12_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hc == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_12_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_12_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hc == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_12_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_12_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hc == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_12_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_12_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hc == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_12_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_12_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hc == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_12_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_12_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hc == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_12_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_12_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hc == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_12_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_12_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hc == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_12_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_12_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hc == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_12_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_12_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hc == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_12_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_12_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hc == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_12_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_12_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hc == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_12_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_12_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hc == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_12_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_13_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hd == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_13_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_13_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hd == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_13_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_13_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hd == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_13_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_13_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hd == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_13_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_13_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hd == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_13_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_13_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hd == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_13_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_13_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hd == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_13_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_13_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hd == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_13_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_13_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hd == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_13_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_13_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hd == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_13_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_13_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hd == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_13_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_13_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hd == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_13_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_13_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hd == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_13_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_13_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hd == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_13_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_13_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hd == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_13_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_14_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'he == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_14_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_14_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'he == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_14_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_14_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'he == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_14_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_14_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'he == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_14_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_14_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'he == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_14_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_14_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'he == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_14_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_14_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'he == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_14_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_14_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'he == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_14_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_14_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'he == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_14_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_14_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'he == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_14_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_14_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'he == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_14_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_14_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'he == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_14_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_14_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'he == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_14_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_14_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'he == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_14_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_14_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'he == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_14_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_15_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hf == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_15_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_15_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hf == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_15_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_15_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hf == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_15_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_15_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hf == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_15_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_15_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hf == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_15_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_15_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hf == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_15_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_15_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hf == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_15_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_15_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hf == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_15_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_15_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hf == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_15_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_15_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hf == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_15_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_15_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hf == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_15_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_15_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hf == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_15_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_15_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hf == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_15_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_15_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hf == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_15_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_15_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'hf == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_15_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_16_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h10 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_16_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_16_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h10 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_16_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_16_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h10 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_16_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_16_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h10 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_16_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_16_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h10 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_16_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_16_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h10 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_16_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_16_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h10 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_16_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_16_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h10 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_16_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_16_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h10 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_16_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_16_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h10 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_16_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_16_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h10 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_16_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_16_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h10 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_16_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_16_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h10 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_16_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_16_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h10 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_16_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_16_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h10 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_16_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_17_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h11 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_17_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_17_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h11 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_17_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_17_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h11 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_17_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_17_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h11 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_17_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_17_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h11 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_17_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_17_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h11 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_17_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_17_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h11 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_17_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_17_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h11 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_17_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_17_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h11 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_17_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_17_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h11 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_17_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_17_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h11 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_17_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_17_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h11 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_17_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_17_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h11 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_17_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_17_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h11 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_17_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_17_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h11 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_17_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_18_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h12 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_18_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_18_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h12 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_18_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_18_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h12 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_18_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_18_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h12 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_18_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_18_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h12 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_18_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_18_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h12 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_18_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_18_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h12 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_18_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_18_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h12 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_18_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_18_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h12 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_18_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_18_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h12 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_18_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_18_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h12 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_18_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_18_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h12 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_18_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_18_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h12 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_18_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_18_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h12 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_18_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_18_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h12 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_18_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_19_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h13 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_19_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_19_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h13 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_19_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_19_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h13 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_19_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_19_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h13 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_19_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_19_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h13 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_19_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_19_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h13 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_19_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_19_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h13 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_19_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_19_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h13 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_19_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_19_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h13 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_19_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_19_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h13 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_19_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_19_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h13 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_19_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_19_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h13 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_19_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_19_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h13 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_19_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_19_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h13 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_19_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_19_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h13 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_19_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_20_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h14 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_20_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_20_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h14 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_20_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_20_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h14 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_20_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_20_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h14 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_20_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_20_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h14 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_20_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_20_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h14 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_20_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_20_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h14 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_20_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_20_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h14 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_20_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_20_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h14 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_20_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_20_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h14 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_20_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_20_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h14 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_20_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_20_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h14 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_20_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_20_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h14 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_20_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_20_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h14 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_20_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_20_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h14 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_20_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_21_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h15 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_21_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_21_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h15 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_21_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_21_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h15 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_21_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_21_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h15 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_21_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_21_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h15 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_21_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_21_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h15 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_21_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_21_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h15 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_21_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_21_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h15 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_21_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_21_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h15 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_21_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_21_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h15 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_21_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_21_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h15 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_21_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_21_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h15 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_21_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_21_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h15 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_21_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_21_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h15 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_21_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_21_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h15 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_21_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_22_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h16 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_22_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_22_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h16 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_22_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_22_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h16 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_22_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_22_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h16 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_22_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_22_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h16 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_22_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_22_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h16 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_22_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_22_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h16 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_22_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_22_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h16 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_22_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_22_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h16 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_22_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_22_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h16 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_22_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_22_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h16 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_22_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_22_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h16 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_22_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_22_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h16 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_22_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_22_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h16 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_22_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_22_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h16 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_22_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_23_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h17 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_23_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_23_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h17 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_23_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_23_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h17 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_23_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_23_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h17 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_23_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_23_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h17 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_23_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_23_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h17 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_23_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_23_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h17 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_23_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_23_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h17 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_23_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_23_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h17 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_23_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_23_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h17 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_23_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_23_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h17 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_23_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_23_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h17 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_23_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_23_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h17 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_23_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_23_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h17 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_23_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_23_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h17 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_23_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_24_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h18 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_24_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_24_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h18 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_24_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_24_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h18 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_24_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_24_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h18 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_24_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_24_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h18 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_24_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_24_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h18 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_24_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_24_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h18 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_24_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_24_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h18 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_24_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_24_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h18 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_24_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_24_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h18 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_24_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_24_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h18 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_24_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_24_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h18 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_24_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_24_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h18 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_24_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_24_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h18 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_24_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_24_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h18 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_24_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_25_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h19 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_25_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_25_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h19 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_25_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_25_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h19 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_25_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_25_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h19 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_25_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_25_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h19 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_25_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_25_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h19 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_25_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_25_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h19 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_25_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_25_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h19 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_25_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_25_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h19 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_25_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_25_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h19 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_25_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_25_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h19 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_25_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_25_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h19 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_25_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_25_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h19 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_25_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_25_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h19 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_25_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_25_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h19 == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_25_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_26_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1a == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_26_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_26_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1a == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_26_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_26_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1a == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_26_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_26_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1a == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_26_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_26_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1a == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_26_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_26_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1a == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_26_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_26_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1a == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_26_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_26_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1a == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_26_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_26_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1a == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_26_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_26_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1a == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_26_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_26_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1a == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_26_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_26_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1a == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_26_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_26_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1a == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_26_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_26_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1a == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_26_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_26_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1a == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_26_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_27_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1b == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_27_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_27_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1b == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_27_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_27_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1b == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_27_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_27_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1b == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_27_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_27_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1b == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_27_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_27_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1b == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_27_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_27_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1b == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_27_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_27_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1b == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_27_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_27_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1b == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_27_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_27_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1b == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_27_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_27_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1b == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_27_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_27_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1b == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_27_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_27_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1b == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_27_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_27_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1b == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_27_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_27_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1b == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_27_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_28_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1c == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_28_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_28_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1c == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_28_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_28_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1c == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_28_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_28_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1c == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_28_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_28_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1c == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_28_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_28_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1c == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_28_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_28_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1c == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_28_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_28_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1c == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_28_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_28_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1c == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_28_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_28_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1c == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_28_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_28_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1c == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_28_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_28_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1c == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_28_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_28_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1c == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_28_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_28_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1c == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_28_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_28_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1c == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_28_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_29_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1d == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_29_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_29_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1d == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_29_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_29_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1d == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_29_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_29_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1d == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_29_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_29_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1d == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_29_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_29_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1d == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_29_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_29_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1d == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_29_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_29_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1d == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_29_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_29_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1d == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_29_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_29_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1d == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_29_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_29_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1d == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_29_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_29_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1d == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_29_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_29_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1d == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_29_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_29_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1d == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_29_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_29_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1d == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_29_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_30_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1e == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_30_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_30_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1e == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_30_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_30_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1e == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_30_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_30_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1e == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_30_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_30_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1e == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_30_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_30_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1e == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_30_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_30_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1e == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_30_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_30_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1e == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_30_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_30_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1e == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_30_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_30_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1e == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_30_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_30_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1e == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_30_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_30_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1e == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_30_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_30_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1e == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_30_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_30_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1e == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_30_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_30_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1e == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_30_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_31_flag_d <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1f == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_31_flag_d <= io_wpte_flag_d; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_31_flag_a <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1f == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_31_flag_a <= io_wpte_flag_a; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_31_flag_g <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1f == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_31_flag_g <= io_wpte_flag_g; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_31_flag_u <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1f == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_31_flag_u <= io_wpte_flag_u; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_31_flag_x <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1f == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_31_flag_x <= io_wpte_flag_x; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_31_flag_w <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1f == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_31_flag_w <= io_wpte_flag_w; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_31_flag_r <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1f == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_31_flag_r <= io_wpte_flag_r; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_31_flag_v <= 1'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1f == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_31_flag_v <= io_wpte_flag_v; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_31_vpn2 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1f == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_31_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_31_vpn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1f == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_31_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_31_vpn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1f == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_31_vpn0 <= io_wvaddr_vpn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_31_ppn2 <= 2'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1f == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_31_ppn2 <= io_wpte_ppn2; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_31_ppn1 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1f == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_31_ppn1 <= io_wpte_ppn1; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_31_ppn0 <= 9'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1f == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_31_ppn0 <= io_wpte_ppn0; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 64:31]
      array4kb_31_asid <= 16'h0; // @[TLB.scala 64:31]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      if (5'h1f == replace_idx) begin // @[TLB.scala 86:33]
        array4kb_31_asid <= io_satp_asid; // @[TLB.scala 86:33]
      end
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_0 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_0 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_0 <= _GEN_1056;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_1 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_1 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_1 <= _GEN_1057;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_2 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_2 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_2 <= _GEN_1058;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_3 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_3 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_3 <= _GEN_1059;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_4 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_4 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_4 <= _GEN_1060;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_5 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_5 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_5 <= _GEN_1061;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_6 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_6 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_6 <= _GEN_1062;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_7 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_7 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_7 <= _GEN_1063;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_8 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_8 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_8 <= _GEN_1064;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_9 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_9 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_9 <= _GEN_1065;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_10 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_10 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_10 <= _GEN_1066;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_11 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_11 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_11 <= _GEN_1067;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_12 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_12 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_12 <= _GEN_1068;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_13 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_13 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_13 <= _GEN_1069;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_14 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_14 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_14 <= _GEN_1070;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_15 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_15 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_15 <= _GEN_1071;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_16 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_16 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_16 <= _GEN_1072;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_17 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_17 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_17 <= _GEN_1073;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_18 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_18 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_18 <= _GEN_1074;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_19 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_19 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_19 <= _GEN_1075;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_20 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_20 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_20 <= _GEN_1076;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_21 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_21 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_21 <= _GEN_1077;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_22 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_22 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_22 <= _GEN_1078;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_23 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_23 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_23 <= _GEN_1079;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_24 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_24 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_24 <= _GEN_1080;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_25 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_25 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_25 <= _GEN_1081;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_26 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_26 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_26 <= _GEN_1082;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_27 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_27 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_27 <= _GEN_1083;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_28 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_28 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_28 <= _GEN_1084;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_29 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_29 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_29 <= _GEN_1085;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_30 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_30 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_30 <= _GEN_1086;
    end
    if (reset) begin // @[TLB.scala 65:31]
      array4kb_valid_31 <= 1'h0; // @[TLB.scala 65:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 89:23]
      array4kb_valid_31 <= 1'h0; // @[TLB.scala 91:25]
    end else if (io_wen & io_wlevel == 2'h0) begin // @[TLB.scala 85:39]
      array4kb_valid_31 <= _GEN_1087;
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_0_flag_d <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h0 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_0_flag_d <= io_wpte_flag_d; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_0_flag_a <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h0 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_0_flag_a <= io_wpte_flag_a; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_0_flag_g <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h0 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_0_flag_g <= io_wpte_flag_g; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_0_flag_u <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h0 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_0_flag_u <= io_wpte_flag_u; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_0_flag_x <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h0 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_0_flag_x <= io_wpte_flag_x; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_0_flag_w <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h0 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_0_flag_w <= io_wpte_flag_w; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_0_flag_r <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h0 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_0_flag_r <= io_wpte_flag_r; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_0_flag_v <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h0 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_0_flag_v <= io_wpte_flag_v; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_0_vpn2 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h0 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_0_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_0_vpn1 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h0 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_0_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_0_ppn2 <= 2'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h0 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_0_ppn2 <= io_wpte_ppn2; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_0_ppn1 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h0 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_0_ppn1 <= io_wpte_ppn1; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_0_asid <= 16'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h0 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_0_asid <= io_satp_asid; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_1_flag_d <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h1 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_1_flag_d <= io_wpte_flag_d; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_1_flag_a <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h1 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_1_flag_a <= io_wpte_flag_a; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_1_flag_g <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h1 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_1_flag_g <= io_wpte_flag_g; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_1_flag_u <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h1 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_1_flag_u <= io_wpte_flag_u; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_1_flag_x <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h1 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_1_flag_x <= io_wpte_flag_x; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_1_flag_w <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h1 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_1_flag_w <= io_wpte_flag_w; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_1_flag_r <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h1 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_1_flag_r <= io_wpte_flag_r; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_1_flag_v <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h1 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_1_flag_v <= io_wpte_flag_v; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_1_vpn2 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h1 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_1_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_1_vpn1 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h1 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_1_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_1_ppn2 <= 2'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h1 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_1_ppn2 <= io_wpte_ppn2; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_1_ppn1 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h1 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_1_ppn1 <= io_wpte_ppn1; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_1_asid <= 16'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h1 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_1_asid <= io_satp_asid; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_2_flag_d <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h2 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_2_flag_d <= io_wpte_flag_d; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_2_flag_a <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h2 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_2_flag_a <= io_wpte_flag_a; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_2_flag_g <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h2 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_2_flag_g <= io_wpte_flag_g; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_2_flag_u <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h2 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_2_flag_u <= io_wpte_flag_u; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_2_flag_x <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h2 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_2_flag_x <= io_wpte_flag_x; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_2_flag_w <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h2 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_2_flag_w <= io_wpte_flag_w; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_2_flag_r <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h2 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_2_flag_r <= io_wpte_flag_r; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_2_flag_v <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h2 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_2_flag_v <= io_wpte_flag_v; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_2_vpn2 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h2 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_2_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_2_vpn1 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h2 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_2_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_2_ppn2 <= 2'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h2 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_2_ppn2 <= io_wpte_ppn2; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_2_ppn1 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h2 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_2_ppn1 <= io_wpte_ppn1; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_2_asid <= 16'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h2 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_2_asid <= io_satp_asid; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_3_flag_d <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h3 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_3_flag_d <= io_wpte_flag_d; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_3_flag_a <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h3 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_3_flag_a <= io_wpte_flag_a; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_3_flag_g <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h3 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_3_flag_g <= io_wpte_flag_g; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_3_flag_u <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h3 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_3_flag_u <= io_wpte_flag_u; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_3_flag_x <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h3 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_3_flag_x <= io_wpte_flag_x; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_3_flag_w <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h3 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_3_flag_w <= io_wpte_flag_w; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_3_flag_r <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h3 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_3_flag_r <= io_wpte_flag_r; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_3_flag_v <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h3 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_3_flag_v <= io_wpte_flag_v; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_3_vpn2 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h3 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_3_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_3_vpn1 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h3 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_3_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_3_ppn2 <= 2'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h3 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_3_ppn2 <= io_wpte_ppn2; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_3_ppn1 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h3 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_3_ppn1 <= io_wpte_ppn1; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_3_asid <= 16'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h3 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_3_asid <= io_satp_asid; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_4_flag_d <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h4 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_4_flag_d <= io_wpte_flag_d; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_4_flag_a <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h4 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_4_flag_a <= io_wpte_flag_a; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_4_flag_g <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h4 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_4_flag_g <= io_wpte_flag_g; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_4_flag_u <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h4 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_4_flag_u <= io_wpte_flag_u; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_4_flag_x <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h4 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_4_flag_x <= io_wpte_flag_x; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_4_flag_w <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h4 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_4_flag_w <= io_wpte_flag_w; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_4_flag_r <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h4 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_4_flag_r <= io_wpte_flag_r; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_4_flag_v <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h4 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_4_flag_v <= io_wpte_flag_v; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_4_vpn2 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h4 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_4_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_4_vpn1 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h4 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_4_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_4_ppn2 <= 2'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h4 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_4_ppn2 <= io_wpte_ppn2; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_4_ppn1 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h4 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_4_ppn1 <= io_wpte_ppn1; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_4_asid <= 16'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h4 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_4_asid <= io_satp_asid; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_5_flag_d <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h5 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_5_flag_d <= io_wpte_flag_d; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_5_flag_a <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h5 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_5_flag_a <= io_wpte_flag_a; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_5_flag_g <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h5 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_5_flag_g <= io_wpte_flag_g; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_5_flag_u <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h5 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_5_flag_u <= io_wpte_flag_u; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_5_flag_x <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h5 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_5_flag_x <= io_wpte_flag_x; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_5_flag_w <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h5 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_5_flag_w <= io_wpte_flag_w; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_5_flag_r <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h5 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_5_flag_r <= io_wpte_flag_r; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_5_flag_v <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h5 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_5_flag_v <= io_wpte_flag_v; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_5_vpn2 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h5 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_5_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_5_vpn1 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h5 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_5_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_5_ppn2 <= 2'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h5 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_5_ppn2 <= io_wpte_ppn2; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_5_ppn1 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h5 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_5_ppn1 <= io_wpte_ppn1; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_5_asid <= 16'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h5 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_5_asid <= io_satp_asid; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_6_flag_d <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h6 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_6_flag_d <= io_wpte_flag_d; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_6_flag_a <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h6 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_6_flag_a <= io_wpte_flag_a; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_6_flag_g <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h6 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_6_flag_g <= io_wpte_flag_g; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_6_flag_u <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h6 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_6_flag_u <= io_wpte_flag_u; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_6_flag_x <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h6 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_6_flag_x <= io_wpte_flag_x; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_6_flag_w <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h6 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_6_flag_w <= io_wpte_flag_w; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_6_flag_r <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h6 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_6_flag_r <= io_wpte_flag_r; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_6_flag_v <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h6 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_6_flag_v <= io_wpte_flag_v; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_6_vpn2 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h6 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_6_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_6_vpn1 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h6 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_6_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_6_ppn2 <= 2'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h6 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_6_ppn2 <= io_wpte_ppn2; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_6_ppn1 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h6 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_6_ppn1 <= io_wpte_ppn1; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_6_asid <= 16'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h6 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_6_asid <= io_satp_asid; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_7_flag_d <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h7 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_7_flag_d <= io_wpte_flag_d; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_7_flag_a <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h7 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_7_flag_a <= io_wpte_flag_a; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_7_flag_g <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h7 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_7_flag_g <= io_wpte_flag_g; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_7_flag_u <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h7 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_7_flag_u <= io_wpte_flag_u; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_7_flag_x <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h7 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_7_flag_x <= io_wpte_flag_x; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_7_flag_w <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h7 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_7_flag_w <= io_wpte_flag_w; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_7_flag_r <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h7 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_7_flag_r <= io_wpte_flag_r; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_7_flag_v <= 1'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h7 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_7_flag_v <= io_wpte_flag_v; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_7_vpn2 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h7 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_7_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_7_vpn1 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h7 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_7_vpn1 <= io_wvaddr_vpn1; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_7_ppn2 <= 2'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h7 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_7_ppn2 <= io_wpte_ppn2; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_7_ppn1 <= 9'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h7 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_7_ppn1 <= io_wpte_ppn1; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 98:31]
      array2mb_7_asid <= 16'h0; // @[TLB.scala 98:31]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      if (3'h7 == replace_idx[2:0]) begin // @[TLB.scala 118:33]
        array2mb_7_asid <= io_satp_asid; // @[TLB.scala 118:33]
      end
    end
    if (reset) begin // @[TLB.scala 99:31]
      array2mb_valid_0 <= 1'h0; // @[TLB.scala 99:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 121:23]
      array2mb_valid_0 <= 1'h0; // @[TLB.scala 123:25]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      array2mb_valid_0 <= _GEN_1896;
    end
    if (reset) begin // @[TLB.scala 99:31]
      array2mb_valid_1 <= 1'h0; // @[TLB.scala 99:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 121:23]
      array2mb_valid_1 <= 1'h0; // @[TLB.scala 123:25]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      array2mb_valid_1 <= _GEN_1897;
    end
    if (reset) begin // @[TLB.scala 99:31]
      array2mb_valid_2 <= 1'h0; // @[TLB.scala 99:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 121:23]
      array2mb_valid_2 <= 1'h0; // @[TLB.scala 123:25]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      array2mb_valid_2 <= _GEN_1898;
    end
    if (reset) begin // @[TLB.scala 99:31]
      array2mb_valid_3 <= 1'h0; // @[TLB.scala 99:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 121:23]
      array2mb_valid_3 <= 1'h0; // @[TLB.scala 123:25]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      array2mb_valid_3 <= _GEN_1899;
    end
    if (reset) begin // @[TLB.scala 99:31]
      array2mb_valid_4 <= 1'h0; // @[TLB.scala 99:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 121:23]
      array2mb_valid_4 <= 1'h0; // @[TLB.scala 123:25]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      array2mb_valid_4 <= _GEN_1900;
    end
    if (reset) begin // @[TLB.scala 99:31]
      array2mb_valid_5 <= 1'h0; // @[TLB.scala 99:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 121:23]
      array2mb_valid_5 <= 1'h0; // @[TLB.scala 123:25]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      array2mb_valid_5 <= _GEN_1901;
    end
    if (reset) begin // @[TLB.scala 99:31]
      array2mb_valid_6 <= 1'h0; // @[TLB.scala 99:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 121:23]
      array2mb_valid_6 <= 1'h0; // @[TLB.scala 123:25]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      array2mb_valid_6 <= _GEN_1902;
    end
    if (reset) begin // @[TLB.scala 99:31]
      array2mb_valid_7 <= 1'h0; // @[TLB.scala 99:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 121:23]
      array2mb_valid_7 <= 1'h0; // @[TLB.scala 123:25]
    end else if (io_wen & io_wlevel == 2'h1) begin // @[TLB.scala 117:39]
      array2mb_valid_7 <= _GEN_1903;
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_0_flag_d <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h0 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_0_flag_d <= io_wpte_flag_d; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_0_flag_a <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h0 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_0_flag_a <= io_wpte_flag_a; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_0_flag_g <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h0 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_0_flag_g <= io_wpte_flag_g; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_0_flag_u <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h0 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_0_flag_u <= io_wpte_flag_u; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_0_flag_x <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h0 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_0_flag_x <= io_wpte_flag_x; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_0_flag_w <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h0 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_0_flag_w <= io_wpte_flag_w; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_0_flag_r <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h0 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_0_flag_r <= io_wpte_flag_r; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_0_flag_v <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h0 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_0_flag_v <= io_wpte_flag_v; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_0_vpn2 <= 9'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h0 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_0_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_0_ppn2 <= 2'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h0 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_0_ppn2 <= io_wpte_ppn2; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_0_asid <= 16'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h0 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_0_asid <= io_satp_asid; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_1_flag_d <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h1 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_1_flag_d <= io_wpte_flag_d; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_1_flag_a <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h1 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_1_flag_a <= io_wpte_flag_a; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_1_flag_g <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h1 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_1_flag_g <= io_wpte_flag_g; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_1_flag_u <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h1 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_1_flag_u <= io_wpte_flag_u; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_1_flag_x <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h1 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_1_flag_x <= io_wpte_flag_x; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_1_flag_w <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h1 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_1_flag_w <= io_wpte_flag_w; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_1_flag_r <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h1 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_1_flag_r <= io_wpte_flag_r; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_1_flag_v <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h1 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_1_flag_v <= io_wpte_flag_v; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_1_vpn2 <= 9'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h1 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_1_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_1_ppn2 <= 2'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h1 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_1_ppn2 <= io_wpte_ppn2; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_1_asid <= 16'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h1 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_1_asid <= io_satp_asid; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_2_flag_d <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h2 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_2_flag_d <= io_wpte_flag_d; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_2_flag_a <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h2 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_2_flag_a <= io_wpte_flag_a; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_2_flag_g <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h2 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_2_flag_g <= io_wpte_flag_g; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_2_flag_u <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h2 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_2_flag_u <= io_wpte_flag_u; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_2_flag_x <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h2 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_2_flag_x <= io_wpte_flag_x; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_2_flag_w <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h2 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_2_flag_w <= io_wpte_flag_w; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_2_flag_r <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h2 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_2_flag_r <= io_wpte_flag_r; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_2_flag_v <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h2 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_2_flag_v <= io_wpte_flag_v; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_2_vpn2 <= 9'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h2 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_2_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_2_ppn2 <= 2'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h2 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_2_ppn2 <= io_wpte_ppn2; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_2_asid <= 16'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h2 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_2_asid <= io_satp_asid; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_3_flag_d <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h3 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_3_flag_d <= io_wpte_flag_d; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_3_flag_a <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h3 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_3_flag_a <= io_wpte_flag_a; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_3_flag_g <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h3 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_3_flag_g <= io_wpte_flag_g; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_3_flag_u <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h3 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_3_flag_u <= io_wpte_flag_u; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_3_flag_x <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h3 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_3_flag_x <= io_wpte_flag_x; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_3_flag_w <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h3 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_3_flag_w <= io_wpte_flag_w; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_3_flag_r <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h3 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_3_flag_r <= io_wpte_flag_r; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_3_flag_v <= 1'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h3 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_3_flag_v <= io_wpte_flag_v; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_3_vpn2 <= 9'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h3 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_3_vpn2 <= io_wvaddr_vpn2; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_3_ppn2 <= 2'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h3 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_3_ppn2 <= io_wpte_ppn2; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 130:31]
      array1gb_3_asid <= 16'h0; // @[TLB.scala 130:31]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      if (2'h3 == replace_idx[1:0]) begin // @[TLB.scala 148:33]
        array1gb_3_asid <= io_satp_asid; // @[TLB.scala 148:33]
      end
    end
    if (reset) begin // @[TLB.scala 131:31]
      array1gb_valid_0 <= 1'h0; // @[TLB.scala 131:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 151:23]
      array1gb_valid_0 <= 1'h0; // @[TLB.scala 153:25]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      array1gb_valid_0 <= _GEN_2132;
    end
    if (reset) begin // @[TLB.scala 131:31]
      array1gb_valid_1 <= 1'h0; // @[TLB.scala 131:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 151:23]
      array1gb_valid_1 <= 1'h0; // @[TLB.scala 153:25]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      array1gb_valid_1 <= _GEN_2133;
    end
    if (reset) begin // @[TLB.scala 131:31]
      array1gb_valid_2 <= 1'h0; // @[TLB.scala 131:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 151:23]
      array1gb_valid_2 <= 1'h0; // @[TLB.scala 153:25]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      array1gb_valid_2 <= _GEN_2134;
    end
    if (reset) begin // @[TLB.scala 131:31]
      array1gb_valid_3 <= 1'h0; // @[TLB.scala 131:31]
    end else if (io_sfence_vma) begin // @[TLB.scala 151:23]
      array1gb_valid_3 <= 1'h0; // @[TLB.scala 153:25]
    end else if (io_wen & io_wlevel == 2'h2) begin // @[TLB.scala 147:39]
      array1gb_valid_3 <= _GEN_2135;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_rlevel != 2'h3)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at TLB.scala:48 assert(io.rlevel =/= 3.U)\n"); // @[TLB.scala 48:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~reset & ~(io_rlevel != 2'h3)) begin
          $fatal; // @[TLB.scala 48:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2 & ~(io_wlevel != 2'h3)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at TLB.scala:49 assert(io.wlevel =/= 3.U)\n"); // @[TLB.scala 49:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_2 & ~(io_wlevel != 2'h3)) begin
          $fatal; // @[TLB.scala 49:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  array4kb_0_flag_d = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  array4kb_0_flag_a = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  array4kb_0_flag_g = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  array4kb_0_flag_u = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  array4kb_0_flag_x = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  array4kb_0_flag_w = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  array4kb_0_flag_r = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  array4kb_0_flag_v = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  array4kb_0_vpn2 = _RAND_8[8:0];
  _RAND_9 = {1{`RANDOM}};
  array4kb_0_vpn1 = _RAND_9[8:0];
  _RAND_10 = {1{`RANDOM}};
  array4kb_0_vpn0 = _RAND_10[8:0];
  _RAND_11 = {1{`RANDOM}};
  array4kb_0_ppn2 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  array4kb_0_ppn1 = _RAND_12[8:0];
  _RAND_13 = {1{`RANDOM}};
  array4kb_0_ppn0 = _RAND_13[8:0];
  _RAND_14 = {1{`RANDOM}};
  array4kb_0_asid = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  array4kb_1_flag_d = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  array4kb_1_flag_a = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  array4kb_1_flag_g = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  array4kb_1_flag_u = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  array4kb_1_flag_x = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  array4kb_1_flag_w = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  array4kb_1_flag_r = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  array4kb_1_flag_v = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  array4kb_1_vpn2 = _RAND_23[8:0];
  _RAND_24 = {1{`RANDOM}};
  array4kb_1_vpn1 = _RAND_24[8:0];
  _RAND_25 = {1{`RANDOM}};
  array4kb_1_vpn0 = _RAND_25[8:0];
  _RAND_26 = {1{`RANDOM}};
  array4kb_1_ppn2 = _RAND_26[1:0];
  _RAND_27 = {1{`RANDOM}};
  array4kb_1_ppn1 = _RAND_27[8:0];
  _RAND_28 = {1{`RANDOM}};
  array4kb_1_ppn0 = _RAND_28[8:0];
  _RAND_29 = {1{`RANDOM}};
  array4kb_1_asid = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  array4kb_2_flag_d = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  array4kb_2_flag_a = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  array4kb_2_flag_g = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  array4kb_2_flag_u = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  array4kb_2_flag_x = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  array4kb_2_flag_w = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  array4kb_2_flag_r = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  array4kb_2_flag_v = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  array4kb_2_vpn2 = _RAND_38[8:0];
  _RAND_39 = {1{`RANDOM}};
  array4kb_2_vpn1 = _RAND_39[8:0];
  _RAND_40 = {1{`RANDOM}};
  array4kb_2_vpn0 = _RAND_40[8:0];
  _RAND_41 = {1{`RANDOM}};
  array4kb_2_ppn2 = _RAND_41[1:0];
  _RAND_42 = {1{`RANDOM}};
  array4kb_2_ppn1 = _RAND_42[8:0];
  _RAND_43 = {1{`RANDOM}};
  array4kb_2_ppn0 = _RAND_43[8:0];
  _RAND_44 = {1{`RANDOM}};
  array4kb_2_asid = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  array4kb_3_flag_d = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  array4kb_3_flag_a = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  array4kb_3_flag_g = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  array4kb_3_flag_u = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  array4kb_3_flag_x = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  array4kb_3_flag_w = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  array4kb_3_flag_r = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  array4kb_3_flag_v = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  array4kb_3_vpn2 = _RAND_53[8:0];
  _RAND_54 = {1{`RANDOM}};
  array4kb_3_vpn1 = _RAND_54[8:0];
  _RAND_55 = {1{`RANDOM}};
  array4kb_3_vpn0 = _RAND_55[8:0];
  _RAND_56 = {1{`RANDOM}};
  array4kb_3_ppn2 = _RAND_56[1:0];
  _RAND_57 = {1{`RANDOM}};
  array4kb_3_ppn1 = _RAND_57[8:0];
  _RAND_58 = {1{`RANDOM}};
  array4kb_3_ppn0 = _RAND_58[8:0];
  _RAND_59 = {1{`RANDOM}};
  array4kb_3_asid = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  array4kb_4_flag_d = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  array4kb_4_flag_a = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  array4kb_4_flag_g = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  array4kb_4_flag_u = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  array4kb_4_flag_x = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  array4kb_4_flag_w = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  array4kb_4_flag_r = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  array4kb_4_flag_v = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  array4kb_4_vpn2 = _RAND_68[8:0];
  _RAND_69 = {1{`RANDOM}};
  array4kb_4_vpn1 = _RAND_69[8:0];
  _RAND_70 = {1{`RANDOM}};
  array4kb_4_vpn0 = _RAND_70[8:0];
  _RAND_71 = {1{`RANDOM}};
  array4kb_4_ppn2 = _RAND_71[1:0];
  _RAND_72 = {1{`RANDOM}};
  array4kb_4_ppn1 = _RAND_72[8:0];
  _RAND_73 = {1{`RANDOM}};
  array4kb_4_ppn0 = _RAND_73[8:0];
  _RAND_74 = {1{`RANDOM}};
  array4kb_4_asid = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  array4kb_5_flag_d = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  array4kb_5_flag_a = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  array4kb_5_flag_g = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  array4kb_5_flag_u = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  array4kb_5_flag_x = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  array4kb_5_flag_w = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  array4kb_5_flag_r = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  array4kb_5_flag_v = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  array4kb_5_vpn2 = _RAND_83[8:0];
  _RAND_84 = {1{`RANDOM}};
  array4kb_5_vpn1 = _RAND_84[8:0];
  _RAND_85 = {1{`RANDOM}};
  array4kb_5_vpn0 = _RAND_85[8:0];
  _RAND_86 = {1{`RANDOM}};
  array4kb_5_ppn2 = _RAND_86[1:0];
  _RAND_87 = {1{`RANDOM}};
  array4kb_5_ppn1 = _RAND_87[8:0];
  _RAND_88 = {1{`RANDOM}};
  array4kb_5_ppn0 = _RAND_88[8:0];
  _RAND_89 = {1{`RANDOM}};
  array4kb_5_asid = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  array4kb_6_flag_d = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  array4kb_6_flag_a = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  array4kb_6_flag_g = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  array4kb_6_flag_u = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  array4kb_6_flag_x = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  array4kb_6_flag_w = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  array4kb_6_flag_r = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  array4kb_6_flag_v = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  array4kb_6_vpn2 = _RAND_98[8:0];
  _RAND_99 = {1{`RANDOM}};
  array4kb_6_vpn1 = _RAND_99[8:0];
  _RAND_100 = {1{`RANDOM}};
  array4kb_6_vpn0 = _RAND_100[8:0];
  _RAND_101 = {1{`RANDOM}};
  array4kb_6_ppn2 = _RAND_101[1:0];
  _RAND_102 = {1{`RANDOM}};
  array4kb_6_ppn1 = _RAND_102[8:0];
  _RAND_103 = {1{`RANDOM}};
  array4kb_6_ppn0 = _RAND_103[8:0];
  _RAND_104 = {1{`RANDOM}};
  array4kb_6_asid = _RAND_104[15:0];
  _RAND_105 = {1{`RANDOM}};
  array4kb_7_flag_d = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  array4kb_7_flag_a = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  array4kb_7_flag_g = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  array4kb_7_flag_u = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  array4kb_7_flag_x = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  array4kb_7_flag_w = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  array4kb_7_flag_r = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  array4kb_7_flag_v = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  array4kb_7_vpn2 = _RAND_113[8:0];
  _RAND_114 = {1{`RANDOM}};
  array4kb_7_vpn1 = _RAND_114[8:0];
  _RAND_115 = {1{`RANDOM}};
  array4kb_7_vpn0 = _RAND_115[8:0];
  _RAND_116 = {1{`RANDOM}};
  array4kb_7_ppn2 = _RAND_116[1:0];
  _RAND_117 = {1{`RANDOM}};
  array4kb_7_ppn1 = _RAND_117[8:0];
  _RAND_118 = {1{`RANDOM}};
  array4kb_7_ppn0 = _RAND_118[8:0];
  _RAND_119 = {1{`RANDOM}};
  array4kb_7_asid = _RAND_119[15:0];
  _RAND_120 = {1{`RANDOM}};
  array4kb_8_flag_d = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  array4kb_8_flag_a = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  array4kb_8_flag_g = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  array4kb_8_flag_u = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  array4kb_8_flag_x = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  array4kb_8_flag_w = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  array4kb_8_flag_r = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  array4kb_8_flag_v = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  array4kb_8_vpn2 = _RAND_128[8:0];
  _RAND_129 = {1{`RANDOM}};
  array4kb_8_vpn1 = _RAND_129[8:0];
  _RAND_130 = {1{`RANDOM}};
  array4kb_8_vpn0 = _RAND_130[8:0];
  _RAND_131 = {1{`RANDOM}};
  array4kb_8_ppn2 = _RAND_131[1:0];
  _RAND_132 = {1{`RANDOM}};
  array4kb_8_ppn1 = _RAND_132[8:0];
  _RAND_133 = {1{`RANDOM}};
  array4kb_8_ppn0 = _RAND_133[8:0];
  _RAND_134 = {1{`RANDOM}};
  array4kb_8_asid = _RAND_134[15:0];
  _RAND_135 = {1{`RANDOM}};
  array4kb_9_flag_d = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  array4kb_9_flag_a = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  array4kb_9_flag_g = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  array4kb_9_flag_u = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  array4kb_9_flag_x = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  array4kb_9_flag_w = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  array4kb_9_flag_r = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  array4kb_9_flag_v = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  array4kb_9_vpn2 = _RAND_143[8:0];
  _RAND_144 = {1{`RANDOM}};
  array4kb_9_vpn1 = _RAND_144[8:0];
  _RAND_145 = {1{`RANDOM}};
  array4kb_9_vpn0 = _RAND_145[8:0];
  _RAND_146 = {1{`RANDOM}};
  array4kb_9_ppn2 = _RAND_146[1:0];
  _RAND_147 = {1{`RANDOM}};
  array4kb_9_ppn1 = _RAND_147[8:0];
  _RAND_148 = {1{`RANDOM}};
  array4kb_9_ppn0 = _RAND_148[8:0];
  _RAND_149 = {1{`RANDOM}};
  array4kb_9_asid = _RAND_149[15:0];
  _RAND_150 = {1{`RANDOM}};
  array4kb_10_flag_d = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  array4kb_10_flag_a = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  array4kb_10_flag_g = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  array4kb_10_flag_u = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  array4kb_10_flag_x = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  array4kb_10_flag_w = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  array4kb_10_flag_r = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  array4kb_10_flag_v = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  array4kb_10_vpn2 = _RAND_158[8:0];
  _RAND_159 = {1{`RANDOM}};
  array4kb_10_vpn1 = _RAND_159[8:0];
  _RAND_160 = {1{`RANDOM}};
  array4kb_10_vpn0 = _RAND_160[8:0];
  _RAND_161 = {1{`RANDOM}};
  array4kb_10_ppn2 = _RAND_161[1:0];
  _RAND_162 = {1{`RANDOM}};
  array4kb_10_ppn1 = _RAND_162[8:0];
  _RAND_163 = {1{`RANDOM}};
  array4kb_10_ppn0 = _RAND_163[8:0];
  _RAND_164 = {1{`RANDOM}};
  array4kb_10_asid = _RAND_164[15:0];
  _RAND_165 = {1{`RANDOM}};
  array4kb_11_flag_d = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  array4kb_11_flag_a = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  array4kb_11_flag_g = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  array4kb_11_flag_u = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  array4kb_11_flag_x = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  array4kb_11_flag_w = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  array4kb_11_flag_r = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  array4kb_11_flag_v = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  array4kb_11_vpn2 = _RAND_173[8:0];
  _RAND_174 = {1{`RANDOM}};
  array4kb_11_vpn1 = _RAND_174[8:0];
  _RAND_175 = {1{`RANDOM}};
  array4kb_11_vpn0 = _RAND_175[8:0];
  _RAND_176 = {1{`RANDOM}};
  array4kb_11_ppn2 = _RAND_176[1:0];
  _RAND_177 = {1{`RANDOM}};
  array4kb_11_ppn1 = _RAND_177[8:0];
  _RAND_178 = {1{`RANDOM}};
  array4kb_11_ppn0 = _RAND_178[8:0];
  _RAND_179 = {1{`RANDOM}};
  array4kb_11_asid = _RAND_179[15:0];
  _RAND_180 = {1{`RANDOM}};
  array4kb_12_flag_d = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  array4kb_12_flag_a = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  array4kb_12_flag_g = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  array4kb_12_flag_u = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  array4kb_12_flag_x = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  array4kb_12_flag_w = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  array4kb_12_flag_r = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  array4kb_12_flag_v = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  array4kb_12_vpn2 = _RAND_188[8:0];
  _RAND_189 = {1{`RANDOM}};
  array4kb_12_vpn1 = _RAND_189[8:0];
  _RAND_190 = {1{`RANDOM}};
  array4kb_12_vpn0 = _RAND_190[8:0];
  _RAND_191 = {1{`RANDOM}};
  array4kb_12_ppn2 = _RAND_191[1:0];
  _RAND_192 = {1{`RANDOM}};
  array4kb_12_ppn1 = _RAND_192[8:0];
  _RAND_193 = {1{`RANDOM}};
  array4kb_12_ppn0 = _RAND_193[8:0];
  _RAND_194 = {1{`RANDOM}};
  array4kb_12_asid = _RAND_194[15:0];
  _RAND_195 = {1{`RANDOM}};
  array4kb_13_flag_d = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  array4kb_13_flag_a = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  array4kb_13_flag_g = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  array4kb_13_flag_u = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  array4kb_13_flag_x = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  array4kb_13_flag_w = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  array4kb_13_flag_r = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  array4kb_13_flag_v = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  array4kb_13_vpn2 = _RAND_203[8:0];
  _RAND_204 = {1{`RANDOM}};
  array4kb_13_vpn1 = _RAND_204[8:0];
  _RAND_205 = {1{`RANDOM}};
  array4kb_13_vpn0 = _RAND_205[8:0];
  _RAND_206 = {1{`RANDOM}};
  array4kb_13_ppn2 = _RAND_206[1:0];
  _RAND_207 = {1{`RANDOM}};
  array4kb_13_ppn1 = _RAND_207[8:0];
  _RAND_208 = {1{`RANDOM}};
  array4kb_13_ppn0 = _RAND_208[8:0];
  _RAND_209 = {1{`RANDOM}};
  array4kb_13_asid = _RAND_209[15:0];
  _RAND_210 = {1{`RANDOM}};
  array4kb_14_flag_d = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  array4kb_14_flag_a = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  array4kb_14_flag_g = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  array4kb_14_flag_u = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  array4kb_14_flag_x = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  array4kb_14_flag_w = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  array4kb_14_flag_r = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  array4kb_14_flag_v = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  array4kb_14_vpn2 = _RAND_218[8:0];
  _RAND_219 = {1{`RANDOM}};
  array4kb_14_vpn1 = _RAND_219[8:0];
  _RAND_220 = {1{`RANDOM}};
  array4kb_14_vpn0 = _RAND_220[8:0];
  _RAND_221 = {1{`RANDOM}};
  array4kb_14_ppn2 = _RAND_221[1:0];
  _RAND_222 = {1{`RANDOM}};
  array4kb_14_ppn1 = _RAND_222[8:0];
  _RAND_223 = {1{`RANDOM}};
  array4kb_14_ppn0 = _RAND_223[8:0];
  _RAND_224 = {1{`RANDOM}};
  array4kb_14_asid = _RAND_224[15:0];
  _RAND_225 = {1{`RANDOM}};
  array4kb_15_flag_d = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  array4kb_15_flag_a = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  array4kb_15_flag_g = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  array4kb_15_flag_u = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  array4kb_15_flag_x = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  array4kb_15_flag_w = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  array4kb_15_flag_r = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  array4kb_15_flag_v = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  array4kb_15_vpn2 = _RAND_233[8:0];
  _RAND_234 = {1{`RANDOM}};
  array4kb_15_vpn1 = _RAND_234[8:0];
  _RAND_235 = {1{`RANDOM}};
  array4kb_15_vpn0 = _RAND_235[8:0];
  _RAND_236 = {1{`RANDOM}};
  array4kb_15_ppn2 = _RAND_236[1:0];
  _RAND_237 = {1{`RANDOM}};
  array4kb_15_ppn1 = _RAND_237[8:0];
  _RAND_238 = {1{`RANDOM}};
  array4kb_15_ppn0 = _RAND_238[8:0];
  _RAND_239 = {1{`RANDOM}};
  array4kb_15_asid = _RAND_239[15:0];
  _RAND_240 = {1{`RANDOM}};
  array4kb_16_flag_d = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  array4kb_16_flag_a = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  array4kb_16_flag_g = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  array4kb_16_flag_u = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  array4kb_16_flag_x = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  array4kb_16_flag_w = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  array4kb_16_flag_r = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  array4kb_16_flag_v = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  array4kb_16_vpn2 = _RAND_248[8:0];
  _RAND_249 = {1{`RANDOM}};
  array4kb_16_vpn1 = _RAND_249[8:0];
  _RAND_250 = {1{`RANDOM}};
  array4kb_16_vpn0 = _RAND_250[8:0];
  _RAND_251 = {1{`RANDOM}};
  array4kb_16_ppn2 = _RAND_251[1:0];
  _RAND_252 = {1{`RANDOM}};
  array4kb_16_ppn1 = _RAND_252[8:0];
  _RAND_253 = {1{`RANDOM}};
  array4kb_16_ppn0 = _RAND_253[8:0];
  _RAND_254 = {1{`RANDOM}};
  array4kb_16_asid = _RAND_254[15:0];
  _RAND_255 = {1{`RANDOM}};
  array4kb_17_flag_d = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  array4kb_17_flag_a = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  array4kb_17_flag_g = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  array4kb_17_flag_u = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  array4kb_17_flag_x = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  array4kb_17_flag_w = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  array4kb_17_flag_r = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  array4kb_17_flag_v = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  array4kb_17_vpn2 = _RAND_263[8:0];
  _RAND_264 = {1{`RANDOM}};
  array4kb_17_vpn1 = _RAND_264[8:0];
  _RAND_265 = {1{`RANDOM}};
  array4kb_17_vpn0 = _RAND_265[8:0];
  _RAND_266 = {1{`RANDOM}};
  array4kb_17_ppn2 = _RAND_266[1:0];
  _RAND_267 = {1{`RANDOM}};
  array4kb_17_ppn1 = _RAND_267[8:0];
  _RAND_268 = {1{`RANDOM}};
  array4kb_17_ppn0 = _RAND_268[8:0];
  _RAND_269 = {1{`RANDOM}};
  array4kb_17_asid = _RAND_269[15:0];
  _RAND_270 = {1{`RANDOM}};
  array4kb_18_flag_d = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  array4kb_18_flag_a = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  array4kb_18_flag_g = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  array4kb_18_flag_u = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  array4kb_18_flag_x = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  array4kb_18_flag_w = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  array4kb_18_flag_r = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  array4kb_18_flag_v = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  array4kb_18_vpn2 = _RAND_278[8:0];
  _RAND_279 = {1{`RANDOM}};
  array4kb_18_vpn1 = _RAND_279[8:0];
  _RAND_280 = {1{`RANDOM}};
  array4kb_18_vpn0 = _RAND_280[8:0];
  _RAND_281 = {1{`RANDOM}};
  array4kb_18_ppn2 = _RAND_281[1:0];
  _RAND_282 = {1{`RANDOM}};
  array4kb_18_ppn1 = _RAND_282[8:0];
  _RAND_283 = {1{`RANDOM}};
  array4kb_18_ppn0 = _RAND_283[8:0];
  _RAND_284 = {1{`RANDOM}};
  array4kb_18_asid = _RAND_284[15:0];
  _RAND_285 = {1{`RANDOM}};
  array4kb_19_flag_d = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  array4kb_19_flag_a = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  array4kb_19_flag_g = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  array4kb_19_flag_u = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  array4kb_19_flag_x = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  array4kb_19_flag_w = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  array4kb_19_flag_r = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  array4kb_19_flag_v = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  array4kb_19_vpn2 = _RAND_293[8:0];
  _RAND_294 = {1{`RANDOM}};
  array4kb_19_vpn1 = _RAND_294[8:0];
  _RAND_295 = {1{`RANDOM}};
  array4kb_19_vpn0 = _RAND_295[8:0];
  _RAND_296 = {1{`RANDOM}};
  array4kb_19_ppn2 = _RAND_296[1:0];
  _RAND_297 = {1{`RANDOM}};
  array4kb_19_ppn1 = _RAND_297[8:0];
  _RAND_298 = {1{`RANDOM}};
  array4kb_19_ppn0 = _RAND_298[8:0];
  _RAND_299 = {1{`RANDOM}};
  array4kb_19_asid = _RAND_299[15:0];
  _RAND_300 = {1{`RANDOM}};
  array4kb_20_flag_d = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  array4kb_20_flag_a = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  array4kb_20_flag_g = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  array4kb_20_flag_u = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  array4kb_20_flag_x = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  array4kb_20_flag_w = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  array4kb_20_flag_r = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  array4kb_20_flag_v = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  array4kb_20_vpn2 = _RAND_308[8:0];
  _RAND_309 = {1{`RANDOM}};
  array4kb_20_vpn1 = _RAND_309[8:0];
  _RAND_310 = {1{`RANDOM}};
  array4kb_20_vpn0 = _RAND_310[8:0];
  _RAND_311 = {1{`RANDOM}};
  array4kb_20_ppn2 = _RAND_311[1:0];
  _RAND_312 = {1{`RANDOM}};
  array4kb_20_ppn1 = _RAND_312[8:0];
  _RAND_313 = {1{`RANDOM}};
  array4kb_20_ppn0 = _RAND_313[8:0];
  _RAND_314 = {1{`RANDOM}};
  array4kb_20_asid = _RAND_314[15:0];
  _RAND_315 = {1{`RANDOM}};
  array4kb_21_flag_d = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  array4kb_21_flag_a = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  array4kb_21_flag_g = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  array4kb_21_flag_u = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  array4kb_21_flag_x = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  array4kb_21_flag_w = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  array4kb_21_flag_r = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  array4kb_21_flag_v = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  array4kb_21_vpn2 = _RAND_323[8:0];
  _RAND_324 = {1{`RANDOM}};
  array4kb_21_vpn1 = _RAND_324[8:0];
  _RAND_325 = {1{`RANDOM}};
  array4kb_21_vpn0 = _RAND_325[8:0];
  _RAND_326 = {1{`RANDOM}};
  array4kb_21_ppn2 = _RAND_326[1:0];
  _RAND_327 = {1{`RANDOM}};
  array4kb_21_ppn1 = _RAND_327[8:0];
  _RAND_328 = {1{`RANDOM}};
  array4kb_21_ppn0 = _RAND_328[8:0];
  _RAND_329 = {1{`RANDOM}};
  array4kb_21_asid = _RAND_329[15:0];
  _RAND_330 = {1{`RANDOM}};
  array4kb_22_flag_d = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  array4kb_22_flag_a = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  array4kb_22_flag_g = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  array4kb_22_flag_u = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  array4kb_22_flag_x = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  array4kb_22_flag_w = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  array4kb_22_flag_r = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  array4kb_22_flag_v = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  array4kb_22_vpn2 = _RAND_338[8:0];
  _RAND_339 = {1{`RANDOM}};
  array4kb_22_vpn1 = _RAND_339[8:0];
  _RAND_340 = {1{`RANDOM}};
  array4kb_22_vpn0 = _RAND_340[8:0];
  _RAND_341 = {1{`RANDOM}};
  array4kb_22_ppn2 = _RAND_341[1:0];
  _RAND_342 = {1{`RANDOM}};
  array4kb_22_ppn1 = _RAND_342[8:0];
  _RAND_343 = {1{`RANDOM}};
  array4kb_22_ppn0 = _RAND_343[8:0];
  _RAND_344 = {1{`RANDOM}};
  array4kb_22_asid = _RAND_344[15:0];
  _RAND_345 = {1{`RANDOM}};
  array4kb_23_flag_d = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  array4kb_23_flag_a = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  array4kb_23_flag_g = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  array4kb_23_flag_u = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  array4kb_23_flag_x = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  array4kb_23_flag_w = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  array4kb_23_flag_r = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  array4kb_23_flag_v = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  array4kb_23_vpn2 = _RAND_353[8:0];
  _RAND_354 = {1{`RANDOM}};
  array4kb_23_vpn1 = _RAND_354[8:0];
  _RAND_355 = {1{`RANDOM}};
  array4kb_23_vpn0 = _RAND_355[8:0];
  _RAND_356 = {1{`RANDOM}};
  array4kb_23_ppn2 = _RAND_356[1:0];
  _RAND_357 = {1{`RANDOM}};
  array4kb_23_ppn1 = _RAND_357[8:0];
  _RAND_358 = {1{`RANDOM}};
  array4kb_23_ppn0 = _RAND_358[8:0];
  _RAND_359 = {1{`RANDOM}};
  array4kb_23_asid = _RAND_359[15:0];
  _RAND_360 = {1{`RANDOM}};
  array4kb_24_flag_d = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  array4kb_24_flag_a = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  array4kb_24_flag_g = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  array4kb_24_flag_u = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  array4kb_24_flag_x = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  array4kb_24_flag_w = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  array4kb_24_flag_r = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  array4kb_24_flag_v = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  array4kb_24_vpn2 = _RAND_368[8:0];
  _RAND_369 = {1{`RANDOM}};
  array4kb_24_vpn1 = _RAND_369[8:0];
  _RAND_370 = {1{`RANDOM}};
  array4kb_24_vpn0 = _RAND_370[8:0];
  _RAND_371 = {1{`RANDOM}};
  array4kb_24_ppn2 = _RAND_371[1:0];
  _RAND_372 = {1{`RANDOM}};
  array4kb_24_ppn1 = _RAND_372[8:0];
  _RAND_373 = {1{`RANDOM}};
  array4kb_24_ppn0 = _RAND_373[8:0];
  _RAND_374 = {1{`RANDOM}};
  array4kb_24_asid = _RAND_374[15:0];
  _RAND_375 = {1{`RANDOM}};
  array4kb_25_flag_d = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  array4kb_25_flag_a = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  array4kb_25_flag_g = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  array4kb_25_flag_u = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  array4kb_25_flag_x = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  array4kb_25_flag_w = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  array4kb_25_flag_r = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  array4kb_25_flag_v = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  array4kb_25_vpn2 = _RAND_383[8:0];
  _RAND_384 = {1{`RANDOM}};
  array4kb_25_vpn1 = _RAND_384[8:0];
  _RAND_385 = {1{`RANDOM}};
  array4kb_25_vpn0 = _RAND_385[8:0];
  _RAND_386 = {1{`RANDOM}};
  array4kb_25_ppn2 = _RAND_386[1:0];
  _RAND_387 = {1{`RANDOM}};
  array4kb_25_ppn1 = _RAND_387[8:0];
  _RAND_388 = {1{`RANDOM}};
  array4kb_25_ppn0 = _RAND_388[8:0];
  _RAND_389 = {1{`RANDOM}};
  array4kb_25_asid = _RAND_389[15:0];
  _RAND_390 = {1{`RANDOM}};
  array4kb_26_flag_d = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  array4kb_26_flag_a = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  array4kb_26_flag_g = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  array4kb_26_flag_u = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  array4kb_26_flag_x = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  array4kb_26_flag_w = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  array4kb_26_flag_r = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  array4kb_26_flag_v = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  array4kb_26_vpn2 = _RAND_398[8:0];
  _RAND_399 = {1{`RANDOM}};
  array4kb_26_vpn1 = _RAND_399[8:0];
  _RAND_400 = {1{`RANDOM}};
  array4kb_26_vpn0 = _RAND_400[8:0];
  _RAND_401 = {1{`RANDOM}};
  array4kb_26_ppn2 = _RAND_401[1:0];
  _RAND_402 = {1{`RANDOM}};
  array4kb_26_ppn1 = _RAND_402[8:0];
  _RAND_403 = {1{`RANDOM}};
  array4kb_26_ppn0 = _RAND_403[8:0];
  _RAND_404 = {1{`RANDOM}};
  array4kb_26_asid = _RAND_404[15:0];
  _RAND_405 = {1{`RANDOM}};
  array4kb_27_flag_d = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  array4kb_27_flag_a = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  array4kb_27_flag_g = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  array4kb_27_flag_u = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  array4kb_27_flag_x = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  array4kb_27_flag_w = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  array4kb_27_flag_r = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  array4kb_27_flag_v = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  array4kb_27_vpn2 = _RAND_413[8:0];
  _RAND_414 = {1{`RANDOM}};
  array4kb_27_vpn1 = _RAND_414[8:0];
  _RAND_415 = {1{`RANDOM}};
  array4kb_27_vpn0 = _RAND_415[8:0];
  _RAND_416 = {1{`RANDOM}};
  array4kb_27_ppn2 = _RAND_416[1:0];
  _RAND_417 = {1{`RANDOM}};
  array4kb_27_ppn1 = _RAND_417[8:0];
  _RAND_418 = {1{`RANDOM}};
  array4kb_27_ppn0 = _RAND_418[8:0];
  _RAND_419 = {1{`RANDOM}};
  array4kb_27_asid = _RAND_419[15:0];
  _RAND_420 = {1{`RANDOM}};
  array4kb_28_flag_d = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  array4kb_28_flag_a = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  array4kb_28_flag_g = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  array4kb_28_flag_u = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  array4kb_28_flag_x = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  array4kb_28_flag_w = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  array4kb_28_flag_r = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  array4kb_28_flag_v = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  array4kb_28_vpn2 = _RAND_428[8:0];
  _RAND_429 = {1{`RANDOM}};
  array4kb_28_vpn1 = _RAND_429[8:0];
  _RAND_430 = {1{`RANDOM}};
  array4kb_28_vpn0 = _RAND_430[8:0];
  _RAND_431 = {1{`RANDOM}};
  array4kb_28_ppn2 = _RAND_431[1:0];
  _RAND_432 = {1{`RANDOM}};
  array4kb_28_ppn1 = _RAND_432[8:0];
  _RAND_433 = {1{`RANDOM}};
  array4kb_28_ppn0 = _RAND_433[8:0];
  _RAND_434 = {1{`RANDOM}};
  array4kb_28_asid = _RAND_434[15:0];
  _RAND_435 = {1{`RANDOM}};
  array4kb_29_flag_d = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  array4kb_29_flag_a = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  array4kb_29_flag_g = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  array4kb_29_flag_u = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  array4kb_29_flag_x = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  array4kb_29_flag_w = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  array4kb_29_flag_r = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  array4kb_29_flag_v = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  array4kb_29_vpn2 = _RAND_443[8:0];
  _RAND_444 = {1{`RANDOM}};
  array4kb_29_vpn1 = _RAND_444[8:0];
  _RAND_445 = {1{`RANDOM}};
  array4kb_29_vpn0 = _RAND_445[8:0];
  _RAND_446 = {1{`RANDOM}};
  array4kb_29_ppn2 = _RAND_446[1:0];
  _RAND_447 = {1{`RANDOM}};
  array4kb_29_ppn1 = _RAND_447[8:0];
  _RAND_448 = {1{`RANDOM}};
  array4kb_29_ppn0 = _RAND_448[8:0];
  _RAND_449 = {1{`RANDOM}};
  array4kb_29_asid = _RAND_449[15:0];
  _RAND_450 = {1{`RANDOM}};
  array4kb_30_flag_d = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  array4kb_30_flag_a = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  array4kb_30_flag_g = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  array4kb_30_flag_u = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  array4kb_30_flag_x = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  array4kb_30_flag_w = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  array4kb_30_flag_r = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  array4kb_30_flag_v = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  array4kb_30_vpn2 = _RAND_458[8:0];
  _RAND_459 = {1{`RANDOM}};
  array4kb_30_vpn1 = _RAND_459[8:0];
  _RAND_460 = {1{`RANDOM}};
  array4kb_30_vpn0 = _RAND_460[8:0];
  _RAND_461 = {1{`RANDOM}};
  array4kb_30_ppn2 = _RAND_461[1:0];
  _RAND_462 = {1{`RANDOM}};
  array4kb_30_ppn1 = _RAND_462[8:0];
  _RAND_463 = {1{`RANDOM}};
  array4kb_30_ppn0 = _RAND_463[8:0];
  _RAND_464 = {1{`RANDOM}};
  array4kb_30_asid = _RAND_464[15:0];
  _RAND_465 = {1{`RANDOM}};
  array4kb_31_flag_d = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  array4kb_31_flag_a = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  array4kb_31_flag_g = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  array4kb_31_flag_u = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  array4kb_31_flag_x = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  array4kb_31_flag_w = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  array4kb_31_flag_r = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  array4kb_31_flag_v = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  array4kb_31_vpn2 = _RAND_473[8:0];
  _RAND_474 = {1{`RANDOM}};
  array4kb_31_vpn1 = _RAND_474[8:0];
  _RAND_475 = {1{`RANDOM}};
  array4kb_31_vpn0 = _RAND_475[8:0];
  _RAND_476 = {1{`RANDOM}};
  array4kb_31_ppn2 = _RAND_476[1:0];
  _RAND_477 = {1{`RANDOM}};
  array4kb_31_ppn1 = _RAND_477[8:0];
  _RAND_478 = {1{`RANDOM}};
  array4kb_31_ppn0 = _RAND_478[8:0];
  _RAND_479 = {1{`RANDOM}};
  array4kb_31_asid = _RAND_479[15:0];
  _RAND_480 = {1{`RANDOM}};
  array4kb_valid_0 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  array4kb_valid_1 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  array4kb_valid_2 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  array4kb_valid_3 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  array4kb_valid_4 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  array4kb_valid_5 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  array4kb_valid_6 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  array4kb_valid_7 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  array4kb_valid_8 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  array4kb_valid_9 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  array4kb_valid_10 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  array4kb_valid_11 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  array4kb_valid_12 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  array4kb_valid_13 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  array4kb_valid_14 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  array4kb_valid_15 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  array4kb_valid_16 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  array4kb_valid_17 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  array4kb_valid_18 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  array4kb_valid_19 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  array4kb_valid_20 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  array4kb_valid_21 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  array4kb_valid_22 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  array4kb_valid_23 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  array4kb_valid_24 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  array4kb_valid_25 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  array4kb_valid_26 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  array4kb_valid_27 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  array4kb_valid_28 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  array4kb_valid_29 = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  array4kb_valid_30 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  array4kb_valid_31 = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  array2mb_0_flag_d = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  array2mb_0_flag_a = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  array2mb_0_flag_g = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  array2mb_0_flag_u = _RAND_515[0:0];
  _RAND_516 = {1{`RANDOM}};
  array2mb_0_flag_x = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  array2mb_0_flag_w = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  array2mb_0_flag_r = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  array2mb_0_flag_v = _RAND_519[0:0];
  _RAND_520 = {1{`RANDOM}};
  array2mb_0_vpn2 = _RAND_520[8:0];
  _RAND_521 = {1{`RANDOM}};
  array2mb_0_vpn1 = _RAND_521[8:0];
  _RAND_522 = {1{`RANDOM}};
  array2mb_0_ppn2 = _RAND_522[1:0];
  _RAND_523 = {1{`RANDOM}};
  array2mb_0_ppn1 = _RAND_523[8:0];
  _RAND_524 = {1{`RANDOM}};
  array2mb_0_asid = _RAND_524[15:0];
  _RAND_525 = {1{`RANDOM}};
  array2mb_1_flag_d = _RAND_525[0:0];
  _RAND_526 = {1{`RANDOM}};
  array2mb_1_flag_a = _RAND_526[0:0];
  _RAND_527 = {1{`RANDOM}};
  array2mb_1_flag_g = _RAND_527[0:0];
  _RAND_528 = {1{`RANDOM}};
  array2mb_1_flag_u = _RAND_528[0:0];
  _RAND_529 = {1{`RANDOM}};
  array2mb_1_flag_x = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  array2mb_1_flag_w = _RAND_530[0:0];
  _RAND_531 = {1{`RANDOM}};
  array2mb_1_flag_r = _RAND_531[0:0];
  _RAND_532 = {1{`RANDOM}};
  array2mb_1_flag_v = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  array2mb_1_vpn2 = _RAND_533[8:0];
  _RAND_534 = {1{`RANDOM}};
  array2mb_1_vpn1 = _RAND_534[8:0];
  _RAND_535 = {1{`RANDOM}};
  array2mb_1_ppn2 = _RAND_535[1:0];
  _RAND_536 = {1{`RANDOM}};
  array2mb_1_ppn1 = _RAND_536[8:0];
  _RAND_537 = {1{`RANDOM}};
  array2mb_1_asid = _RAND_537[15:0];
  _RAND_538 = {1{`RANDOM}};
  array2mb_2_flag_d = _RAND_538[0:0];
  _RAND_539 = {1{`RANDOM}};
  array2mb_2_flag_a = _RAND_539[0:0];
  _RAND_540 = {1{`RANDOM}};
  array2mb_2_flag_g = _RAND_540[0:0];
  _RAND_541 = {1{`RANDOM}};
  array2mb_2_flag_u = _RAND_541[0:0];
  _RAND_542 = {1{`RANDOM}};
  array2mb_2_flag_x = _RAND_542[0:0];
  _RAND_543 = {1{`RANDOM}};
  array2mb_2_flag_w = _RAND_543[0:0];
  _RAND_544 = {1{`RANDOM}};
  array2mb_2_flag_r = _RAND_544[0:0];
  _RAND_545 = {1{`RANDOM}};
  array2mb_2_flag_v = _RAND_545[0:0];
  _RAND_546 = {1{`RANDOM}};
  array2mb_2_vpn2 = _RAND_546[8:0];
  _RAND_547 = {1{`RANDOM}};
  array2mb_2_vpn1 = _RAND_547[8:0];
  _RAND_548 = {1{`RANDOM}};
  array2mb_2_ppn2 = _RAND_548[1:0];
  _RAND_549 = {1{`RANDOM}};
  array2mb_2_ppn1 = _RAND_549[8:0];
  _RAND_550 = {1{`RANDOM}};
  array2mb_2_asid = _RAND_550[15:0];
  _RAND_551 = {1{`RANDOM}};
  array2mb_3_flag_d = _RAND_551[0:0];
  _RAND_552 = {1{`RANDOM}};
  array2mb_3_flag_a = _RAND_552[0:0];
  _RAND_553 = {1{`RANDOM}};
  array2mb_3_flag_g = _RAND_553[0:0];
  _RAND_554 = {1{`RANDOM}};
  array2mb_3_flag_u = _RAND_554[0:0];
  _RAND_555 = {1{`RANDOM}};
  array2mb_3_flag_x = _RAND_555[0:0];
  _RAND_556 = {1{`RANDOM}};
  array2mb_3_flag_w = _RAND_556[0:0];
  _RAND_557 = {1{`RANDOM}};
  array2mb_3_flag_r = _RAND_557[0:0];
  _RAND_558 = {1{`RANDOM}};
  array2mb_3_flag_v = _RAND_558[0:0];
  _RAND_559 = {1{`RANDOM}};
  array2mb_3_vpn2 = _RAND_559[8:0];
  _RAND_560 = {1{`RANDOM}};
  array2mb_3_vpn1 = _RAND_560[8:0];
  _RAND_561 = {1{`RANDOM}};
  array2mb_3_ppn2 = _RAND_561[1:0];
  _RAND_562 = {1{`RANDOM}};
  array2mb_3_ppn1 = _RAND_562[8:0];
  _RAND_563 = {1{`RANDOM}};
  array2mb_3_asid = _RAND_563[15:0];
  _RAND_564 = {1{`RANDOM}};
  array2mb_4_flag_d = _RAND_564[0:0];
  _RAND_565 = {1{`RANDOM}};
  array2mb_4_flag_a = _RAND_565[0:0];
  _RAND_566 = {1{`RANDOM}};
  array2mb_4_flag_g = _RAND_566[0:0];
  _RAND_567 = {1{`RANDOM}};
  array2mb_4_flag_u = _RAND_567[0:0];
  _RAND_568 = {1{`RANDOM}};
  array2mb_4_flag_x = _RAND_568[0:0];
  _RAND_569 = {1{`RANDOM}};
  array2mb_4_flag_w = _RAND_569[0:0];
  _RAND_570 = {1{`RANDOM}};
  array2mb_4_flag_r = _RAND_570[0:0];
  _RAND_571 = {1{`RANDOM}};
  array2mb_4_flag_v = _RAND_571[0:0];
  _RAND_572 = {1{`RANDOM}};
  array2mb_4_vpn2 = _RAND_572[8:0];
  _RAND_573 = {1{`RANDOM}};
  array2mb_4_vpn1 = _RAND_573[8:0];
  _RAND_574 = {1{`RANDOM}};
  array2mb_4_ppn2 = _RAND_574[1:0];
  _RAND_575 = {1{`RANDOM}};
  array2mb_4_ppn1 = _RAND_575[8:0];
  _RAND_576 = {1{`RANDOM}};
  array2mb_4_asid = _RAND_576[15:0];
  _RAND_577 = {1{`RANDOM}};
  array2mb_5_flag_d = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  array2mb_5_flag_a = _RAND_578[0:0];
  _RAND_579 = {1{`RANDOM}};
  array2mb_5_flag_g = _RAND_579[0:0];
  _RAND_580 = {1{`RANDOM}};
  array2mb_5_flag_u = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  array2mb_5_flag_x = _RAND_581[0:0];
  _RAND_582 = {1{`RANDOM}};
  array2mb_5_flag_w = _RAND_582[0:0];
  _RAND_583 = {1{`RANDOM}};
  array2mb_5_flag_r = _RAND_583[0:0];
  _RAND_584 = {1{`RANDOM}};
  array2mb_5_flag_v = _RAND_584[0:0];
  _RAND_585 = {1{`RANDOM}};
  array2mb_5_vpn2 = _RAND_585[8:0];
  _RAND_586 = {1{`RANDOM}};
  array2mb_5_vpn1 = _RAND_586[8:0];
  _RAND_587 = {1{`RANDOM}};
  array2mb_5_ppn2 = _RAND_587[1:0];
  _RAND_588 = {1{`RANDOM}};
  array2mb_5_ppn1 = _RAND_588[8:0];
  _RAND_589 = {1{`RANDOM}};
  array2mb_5_asid = _RAND_589[15:0];
  _RAND_590 = {1{`RANDOM}};
  array2mb_6_flag_d = _RAND_590[0:0];
  _RAND_591 = {1{`RANDOM}};
  array2mb_6_flag_a = _RAND_591[0:0];
  _RAND_592 = {1{`RANDOM}};
  array2mb_6_flag_g = _RAND_592[0:0];
  _RAND_593 = {1{`RANDOM}};
  array2mb_6_flag_u = _RAND_593[0:0];
  _RAND_594 = {1{`RANDOM}};
  array2mb_6_flag_x = _RAND_594[0:0];
  _RAND_595 = {1{`RANDOM}};
  array2mb_6_flag_w = _RAND_595[0:0];
  _RAND_596 = {1{`RANDOM}};
  array2mb_6_flag_r = _RAND_596[0:0];
  _RAND_597 = {1{`RANDOM}};
  array2mb_6_flag_v = _RAND_597[0:0];
  _RAND_598 = {1{`RANDOM}};
  array2mb_6_vpn2 = _RAND_598[8:0];
  _RAND_599 = {1{`RANDOM}};
  array2mb_6_vpn1 = _RAND_599[8:0];
  _RAND_600 = {1{`RANDOM}};
  array2mb_6_ppn2 = _RAND_600[1:0];
  _RAND_601 = {1{`RANDOM}};
  array2mb_6_ppn1 = _RAND_601[8:0];
  _RAND_602 = {1{`RANDOM}};
  array2mb_6_asid = _RAND_602[15:0];
  _RAND_603 = {1{`RANDOM}};
  array2mb_7_flag_d = _RAND_603[0:0];
  _RAND_604 = {1{`RANDOM}};
  array2mb_7_flag_a = _RAND_604[0:0];
  _RAND_605 = {1{`RANDOM}};
  array2mb_7_flag_g = _RAND_605[0:0];
  _RAND_606 = {1{`RANDOM}};
  array2mb_7_flag_u = _RAND_606[0:0];
  _RAND_607 = {1{`RANDOM}};
  array2mb_7_flag_x = _RAND_607[0:0];
  _RAND_608 = {1{`RANDOM}};
  array2mb_7_flag_w = _RAND_608[0:0];
  _RAND_609 = {1{`RANDOM}};
  array2mb_7_flag_r = _RAND_609[0:0];
  _RAND_610 = {1{`RANDOM}};
  array2mb_7_flag_v = _RAND_610[0:0];
  _RAND_611 = {1{`RANDOM}};
  array2mb_7_vpn2 = _RAND_611[8:0];
  _RAND_612 = {1{`RANDOM}};
  array2mb_7_vpn1 = _RAND_612[8:0];
  _RAND_613 = {1{`RANDOM}};
  array2mb_7_ppn2 = _RAND_613[1:0];
  _RAND_614 = {1{`RANDOM}};
  array2mb_7_ppn1 = _RAND_614[8:0];
  _RAND_615 = {1{`RANDOM}};
  array2mb_7_asid = _RAND_615[15:0];
  _RAND_616 = {1{`RANDOM}};
  array2mb_valid_0 = _RAND_616[0:0];
  _RAND_617 = {1{`RANDOM}};
  array2mb_valid_1 = _RAND_617[0:0];
  _RAND_618 = {1{`RANDOM}};
  array2mb_valid_2 = _RAND_618[0:0];
  _RAND_619 = {1{`RANDOM}};
  array2mb_valid_3 = _RAND_619[0:0];
  _RAND_620 = {1{`RANDOM}};
  array2mb_valid_4 = _RAND_620[0:0];
  _RAND_621 = {1{`RANDOM}};
  array2mb_valid_5 = _RAND_621[0:0];
  _RAND_622 = {1{`RANDOM}};
  array2mb_valid_6 = _RAND_622[0:0];
  _RAND_623 = {1{`RANDOM}};
  array2mb_valid_7 = _RAND_623[0:0];
  _RAND_624 = {1{`RANDOM}};
  array1gb_0_flag_d = _RAND_624[0:0];
  _RAND_625 = {1{`RANDOM}};
  array1gb_0_flag_a = _RAND_625[0:0];
  _RAND_626 = {1{`RANDOM}};
  array1gb_0_flag_g = _RAND_626[0:0];
  _RAND_627 = {1{`RANDOM}};
  array1gb_0_flag_u = _RAND_627[0:0];
  _RAND_628 = {1{`RANDOM}};
  array1gb_0_flag_x = _RAND_628[0:0];
  _RAND_629 = {1{`RANDOM}};
  array1gb_0_flag_w = _RAND_629[0:0];
  _RAND_630 = {1{`RANDOM}};
  array1gb_0_flag_r = _RAND_630[0:0];
  _RAND_631 = {1{`RANDOM}};
  array1gb_0_flag_v = _RAND_631[0:0];
  _RAND_632 = {1{`RANDOM}};
  array1gb_0_vpn2 = _RAND_632[8:0];
  _RAND_633 = {1{`RANDOM}};
  array1gb_0_ppn2 = _RAND_633[1:0];
  _RAND_634 = {1{`RANDOM}};
  array1gb_0_asid = _RAND_634[15:0];
  _RAND_635 = {1{`RANDOM}};
  array1gb_1_flag_d = _RAND_635[0:0];
  _RAND_636 = {1{`RANDOM}};
  array1gb_1_flag_a = _RAND_636[0:0];
  _RAND_637 = {1{`RANDOM}};
  array1gb_1_flag_g = _RAND_637[0:0];
  _RAND_638 = {1{`RANDOM}};
  array1gb_1_flag_u = _RAND_638[0:0];
  _RAND_639 = {1{`RANDOM}};
  array1gb_1_flag_x = _RAND_639[0:0];
  _RAND_640 = {1{`RANDOM}};
  array1gb_1_flag_w = _RAND_640[0:0];
  _RAND_641 = {1{`RANDOM}};
  array1gb_1_flag_r = _RAND_641[0:0];
  _RAND_642 = {1{`RANDOM}};
  array1gb_1_flag_v = _RAND_642[0:0];
  _RAND_643 = {1{`RANDOM}};
  array1gb_1_vpn2 = _RAND_643[8:0];
  _RAND_644 = {1{`RANDOM}};
  array1gb_1_ppn2 = _RAND_644[1:0];
  _RAND_645 = {1{`RANDOM}};
  array1gb_1_asid = _RAND_645[15:0];
  _RAND_646 = {1{`RANDOM}};
  array1gb_2_flag_d = _RAND_646[0:0];
  _RAND_647 = {1{`RANDOM}};
  array1gb_2_flag_a = _RAND_647[0:0];
  _RAND_648 = {1{`RANDOM}};
  array1gb_2_flag_g = _RAND_648[0:0];
  _RAND_649 = {1{`RANDOM}};
  array1gb_2_flag_u = _RAND_649[0:0];
  _RAND_650 = {1{`RANDOM}};
  array1gb_2_flag_x = _RAND_650[0:0];
  _RAND_651 = {1{`RANDOM}};
  array1gb_2_flag_w = _RAND_651[0:0];
  _RAND_652 = {1{`RANDOM}};
  array1gb_2_flag_r = _RAND_652[0:0];
  _RAND_653 = {1{`RANDOM}};
  array1gb_2_flag_v = _RAND_653[0:0];
  _RAND_654 = {1{`RANDOM}};
  array1gb_2_vpn2 = _RAND_654[8:0];
  _RAND_655 = {1{`RANDOM}};
  array1gb_2_ppn2 = _RAND_655[1:0];
  _RAND_656 = {1{`RANDOM}};
  array1gb_2_asid = _RAND_656[15:0];
  _RAND_657 = {1{`RANDOM}};
  array1gb_3_flag_d = _RAND_657[0:0];
  _RAND_658 = {1{`RANDOM}};
  array1gb_3_flag_a = _RAND_658[0:0];
  _RAND_659 = {1{`RANDOM}};
  array1gb_3_flag_g = _RAND_659[0:0];
  _RAND_660 = {1{`RANDOM}};
  array1gb_3_flag_u = _RAND_660[0:0];
  _RAND_661 = {1{`RANDOM}};
  array1gb_3_flag_x = _RAND_661[0:0];
  _RAND_662 = {1{`RANDOM}};
  array1gb_3_flag_w = _RAND_662[0:0];
  _RAND_663 = {1{`RANDOM}};
  array1gb_3_flag_r = _RAND_663[0:0];
  _RAND_664 = {1{`RANDOM}};
  array1gb_3_flag_v = _RAND_664[0:0];
  _RAND_665 = {1{`RANDOM}};
  array1gb_3_vpn2 = _RAND_665[8:0];
  _RAND_666 = {1{`RANDOM}};
  array1gb_3_ppn2 = _RAND_666[1:0];
  _RAND_667 = {1{`RANDOM}};
  array1gb_3_asid = _RAND_667[15:0];
  _RAND_668 = {1{`RANDOM}};
  array1gb_valid_0 = _RAND_668[0:0];
  _RAND_669 = {1{`RANDOM}};
  array1gb_valid_1 = _RAND_669[0:0];
  _RAND_670 = {1{`RANDOM}};
  array1gb_valid_2 = _RAND_670[0:0];
  _RAND_671 = {1{`RANDOM}};
  array1gb_valid_3 = _RAND_671[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CachePortProxy(
  input         clock,
  input         reset,
  input  [1:0]  io_prv,
  input         io_sv39_en,
  input  [15:0] io_satp_asid,
  input  [43:0] io_satp_ppn,
  input         io_sfence_vma,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [38:0] io_in_req_bits_addr,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [63:0] io_in_resp_bits_rdata,
  output        io_in_resp_bits_page_fault,
  output        io_in_resp_bits_access_fault,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [38:0] io_out_req_bits_addr,
  output        io_out_resp_ready,
  input         io_out_resp_valid,
  input  [63:0] io_out_resp_bits_rdata,
  input         io_ptw_req_ready,
  output        io_ptw_req_valid,
  output [38:0] io_ptw_req_bits_addr,
  output        io_ptw_resp_ready,
  input         io_ptw_resp_valid,
  input  [63:0] io_ptw_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  wire  tlb_clock; // @[CachePortProxy.scala 28:19]
  wire  tlb_reset; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_sfence_vma; // @[CachePortProxy.scala 28:19]
  wire [8:0] tlb_io_vaddr_vpn2; // @[CachePortProxy.scala 28:19]
  wire [8:0] tlb_io_vaddr_vpn1; // @[CachePortProxy.scala 28:19]
  wire [8:0] tlb_io_vaddr_vpn0; // @[CachePortProxy.scala 28:19]
  wire [1:0] tlb_io_rpte_ppn2; // @[CachePortProxy.scala 28:19]
  wire [8:0] tlb_io_rpte_ppn1; // @[CachePortProxy.scala 28:19]
  wire [8:0] tlb_io_rpte_ppn0; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_rpte_flag_d; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_rpte_flag_a; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_rpte_flag_u; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_rpte_flag_x; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_rpte_flag_w; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_rpte_flag_r; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_rpte_flag_v; // @[CachePortProxy.scala 28:19]
  wire [1:0] tlb_io_rlevel; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_hit; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_wen; // @[CachePortProxy.scala 28:19]
  wire [8:0] tlb_io_wvaddr_vpn2; // @[CachePortProxy.scala 28:19]
  wire [8:0] tlb_io_wvaddr_vpn1; // @[CachePortProxy.scala 28:19]
  wire [8:0] tlb_io_wvaddr_vpn0; // @[CachePortProxy.scala 28:19]
  wire [1:0] tlb_io_wpte_ppn2; // @[CachePortProxy.scala 28:19]
  wire [8:0] tlb_io_wpte_ppn1; // @[CachePortProxy.scala 28:19]
  wire [8:0] tlb_io_wpte_ppn0; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_wpte_flag_d; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_wpte_flag_a; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_wpte_flag_g; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_wpte_flag_u; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_wpte_flag_x; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_wpte_flag_w; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_wpte_flag_r; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_wpte_flag_v; // @[CachePortProxy.scala 28:19]
  wire [1:0] tlb_io_wlevel; // @[CachePortProxy.scala 28:19]
  wire [15:0] tlb_io_satp_asid; // @[CachePortProxy.scala 28:19]
  reg [2:0] state; // @[CachePortProxy.scala 21:93]
  wire  _in_req_bits_T = state == 3'h0; // @[CachePortProxy.scala 24:54]
  reg [38:0] in_req_bits_r_addr; // @[Reg.scala 35:20]
  wire [38:0] _GEN_0 = _in_req_bits_T ? io_in_req_bits_addr : in_req_bits_r_addr; // @[Reg.scala 36:18 35:20 36:22]
  wire [11:0] in_vaddr_offset = _GEN_0[11:0]; // @[CachePortProxy.scala 25:46]
  wire [8:0] in_vaddr_vpn0 = _GEN_0[20:12]; // @[CachePortProxy.scala 25:46]
  wire [8:0] in_vaddr_vpn1 = _GEN_0[29:21]; // @[CachePortProxy.scala 25:46]
  wire [8:0] in_vaddr_vpn2 = _GEN_0[38:30]; // @[CachePortProxy.scala 25:46]
  wire  _atp_en_T_1 = io_prv != 2'h3 & io_sv39_en; // @[CachePortProxy.scala 38:48]
  reg  atp_en_r; // @[Reg.scala 35:20]
  wire  _GEN_7 = _in_req_bits_T ? _atp_en_T_1 : atp_en_r; // @[Reg.scala 36:18 35:20 36:22]
  wire  in_addr_invalid = io_in_req_bits_addr < 39'h10000; // @[CachePortProxy.scala 42:34]
  wire  _access_fault_T_3 = ~_GEN_7; // @[CachePortProxy.scala 43:73]
  wire  access_fault = ~io_in_req_bits_addr[31] & (io_prv == 2'h3 | ~_GEN_7) & in_addr_invalid; // @[CachePortProxy.scala 43:82]
  reg [1:0] ptw_level; // @[CachePortProxy.scala 46:29]
  wire  ptw_pte_flag_v = io_ptw_resp_bits_rdata[0]; // @[CachePortProxy.scala 47:53]
  wire  ptw_pte_flag_r = io_ptw_resp_bits_rdata[1]; // @[CachePortProxy.scala 47:53]
  wire  ptw_pte_flag_w = io_ptw_resp_bits_rdata[2]; // @[CachePortProxy.scala 47:53]
  wire  ptw_pte_flag_x = io_ptw_resp_bits_rdata[3]; // @[CachePortProxy.scala 47:53]
  wire  ptw_pte_flag_u = io_ptw_resp_bits_rdata[4]; // @[CachePortProxy.scala 47:53]
  wire  ptw_pte_flag_g = io_ptw_resp_bits_rdata[5]; // @[CachePortProxy.scala 47:53]
  wire  ptw_pte_flag_a = io_ptw_resp_bits_rdata[6]; // @[CachePortProxy.scala 47:53]
  wire  ptw_pte_flag_d = io_ptw_resp_bits_rdata[7]; // @[CachePortProxy.scala 47:53]
  wire [8:0] ptw_pte_ppn0 = io_ptw_resp_bits_rdata[18:10]; // @[CachePortProxy.scala 47:53]
  wire [8:0] ptw_pte_ppn1 = io_ptw_resp_bits_rdata[27:19]; // @[CachePortProxy.scala 47:53]
  wire [1:0] ptw_pte_ppn2 = io_ptw_resp_bits_rdata[29:28]; // @[CachePortProxy.scala 47:53]
  wire  _ptw_pte_reg_T = io_ptw_resp_ready & io_ptw_resp_valid; // @[Decoupled.scala 51:35]
  reg [1:0] ptw_pte_reg_ppn2; // @[Reg.scala 35:20]
  reg [8:0] ptw_pte_reg_ppn1; // @[Reg.scala 35:20]
  reg [8:0] ptw_pte_reg_ppn0; // @[Reg.scala 35:20]
  reg  ptw_pte_reg_flag_d; // @[Reg.scala 35:20]
  reg  ptw_pte_reg_flag_a; // @[Reg.scala 35:20]
  reg  ptw_pte_reg_flag_g; // @[Reg.scala 35:20]
  reg  ptw_pte_reg_flag_u; // @[Reg.scala 35:20]
  reg  ptw_pte_reg_flag_x; // @[Reg.scala 35:20]
  reg  ptw_pte_reg_flag_w; // @[Reg.scala 35:20]
  reg  ptw_pte_reg_flag_r; // @[Reg.scala 35:20]
  reg  ptw_pte_reg_flag_v; // @[Reg.scala 35:20]
  wire  _ptw_complete_T_4 = ptw_pte_flag_r | ptw_pte_flag_x; // @[CachePortProxy.scala 7:37]
  wire  ptw_complete = ~ptw_pte_flag_v | ~ptw_pte_flag_r & ptw_pte_flag_w | _ptw_complete_T_4 | ptw_level == 2'h0; // @[CachePortProxy.scala 49:96]
  wire  _T_1 = io_in_req_ready & io_in_req_valid; // @[Decoupled.scala 51:35]
  wire  _T_2 = ~tlb_io_hit; // @[CachePortProxy.scala 55:24]
  wire [2:0] _GEN_20 = _GEN_7 & ~tlb_io_hit ? 3'h1 : state; // @[CachePortProxy.scala 55:37 56:17 21:93]
  wire [2:0] _GEN_21 = _T_1 ? _GEN_20 : state; // @[CachePortProxy.scala 54:28 21:93]
  wire  _T_7 = io_ptw_req_ready & io_ptw_req_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _ptw_level_T_1 = ptw_level - 2'h1; // @[CachePortProxy.scala 77:34]
  wire [2:0] _GEN_25 = ptw_complete ? 3'h3 : 3'h1; // @[CachePortProxy.scala 73:28 74:17 76:21]
  wire [1:0] _GEN_26 = ptw_complete ? ptw_level : _ptw_level_T_1; // @[CachePortProxy.scala 73:28 46:29 77:21]
  wire [2:0] _GEN_27 = _ptw_pte_reg_T ? _GEN_25 : state; // @[CachePortProxy.scala 72:30 21:93]
  wire [1:0] _GEN_28 = _ptw_pte_reg_T ? _GEN_26 : ptw_level; // @[CachePortProxy.scala 46:29 72:30]
  wire  _T_11 = io_out_req_ready & io_out_req_valid; // @[Decoupled.scala 51:35]
  wire  pte_flag_v = _in_req_bits_T ? tlb_io_rpte_flag_v : ptw_pte_reg_flag_v; // @[CachePortProxy.scala 117:18]
  wire  pte_flag_r = _in_req_bits_T ? tlb_io_rpte_flag_r : ptw_pte_reg_flag_r; // @[CachePortProxy.scala 117:18]
  wire  pte_flag_w = _in_req_bits_T ? tlb_io_rpte_flag_w : ptw_pte_reg_flag_w; // @[CachePortProxy.scala 117:18]
  wire  pf1 = ~pte_flag_v | ~pte_flag_r & pte_flag_w; // @[CachePortProxy.scala 132:20]
  wire  pte_flag_x = _in_req_bits_T ? tlb_io_rpte_flag_x : ptw_pte_reg_flag_x; // @[CachePortProxy.scala 117:18]
  wire  _T_19 = pte_flag_r | pte_flag_x; // @[CachePortProxy.scala 7:37]
  wire  pte_flag_a = _in_req_bits_T ? tlb_io_rpte_flag_a : ptw_pte_reg_flag_a; // @[CachePortProxy.scala 117:18]
  wire  _T_20 = ~pte_flag_a; // @[CachePortProxy.scala 136:10]
  wire  pf2 = _T_19 & _T_20; // @[CachePortProxy.scala 135:21 128:24]
  reg [1:0] prv_r; // @[Reg.scala 35:20]
  wire [1:0] prv = _in_req_bits_T ? io_prv : prv_r; // @[Utils.scala 50:8]
  wire  pte_flag_u = _in_req_bits_T ? tlb_io_rpte_flag_u : ptw_pte_reg_flag_u; // @[CachePortProxy.scala 117:18]
  wire  _T_23 = prv == 2'h0 & ~pte_flag_u; // @[CachePortProxy.scala 139:26]
  wire  pf3 = _T_19 & _T_23; // @[CachePortProxy.scala 135:21 129:24]
  wire  _T_24 = ~pte_flag_x; // @[CachePortProxy.scala 143:12]
  wire  pf4 = _T_19 & _T_24; // @[CachePortProxy.scala 135:21 130:24]
  wire  _T_25 = state == 3'h3; // @[CachePortProxy.scala 152:16]
  wire [8:0] pte_ppn1 = _in_req_bits_T ? tlb_io_rpte_ppn1 : ptw_pte_reg_ppn1; // @[CachePortProxy.scala 117:18]
  wire [8:0] pte_ppn0 = _in_req_bits_T ? tlb_io_rpte_ppn0 : ptw_pte_reg_ppn0; // @[CachePortProxy.scala 117:18]
  wire [17:0] _T_27 = {pte_ppn1,pte_ppn0}; // @[Cat.scala 33:92]
  wire  _T_33 = ptw_level == 2'h2 & _T_27 != 18'h0 | ptw_level == 2'h1 & pte_ppn0 != 9'h0; // @[CachePortProxy.scala 153:67]
  wire  _GEN_45 = state == 3'h3 & _T_33; // @[CachePortProxy.scala 131:24 152:36]
  wire  pf5 = _T_19 & _GEN_45; // @[CachePortProxy.scala 135:21 131:24]
  wire  page_fault = pf1 | pf2 | pf3 | pf4 | pf5; // @[CachePortProxy.scala 158:42]
  wire [2:0] _GEN_29 = _T_11 | page_fault ? 3'h0 : state; // @[CachePortProxy.scala 82:43 83:15 21:93]
  wire  _T_14 = io_in_resp_ready & io_in_resp_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_30 = _T_14 ? 3'h0 : state; // @[CachePortProxy.scala 87:29 88:15 21:93]
  wire [2:0] _GEN_31 = 3'h4 == state ? _GEN_30 : state; // @[CachePortProxy.scala 52:17 21:93]
  wire [2:0] _GEN_32 = 3'h3 == state ? _GEN_29 : _GEN_31; // @[CachePortProxy.scala 52:17]
  wire [55:0] _l2_addr_T = {io_satp_ppn,in_vaddr_vpn2,3'h0}; // @[Cat.scala 33:92]
  wire [31:0] l1_addr = {ptw_pte_reg_ppn2,ptw_pte_reg_ppn1,ptw_pte_reg_ppn0,in_vaddr_vpn1,3'h0}; // @[Cat.scala 33:92]
  wire [31:0] l0_addr = {ptw_pte_reg_ppn2,ptw_pte_reg_ppn1,ptw_pte_reg_ppn0,in_vaddr_vpn0,3'h0}; // @[Cat.scala 33:92]
  wire [31:0] l2_addr = _l2_addr_T[31:0]; // @[CachePortProxy.scala 94:21 98:11]
  wire [31:0] _io_ptw_req_bits_addr_T_1 = 2'h2 == ptw_level ? l2_addr : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] _io_ptw_req_bits_addr_T_3 = 2'h1 == ptw_level ? l1_addr : _io_ptw_req_bits_addr_T_1; // @[Mux.scala 81:58]
  wire [31:0] _io_ptw_req_bits_addr_T_5 = 2'h0 == ptw_level ? l0_addr : _io_ptw_req_bits_addr_T_3; // @[Mux.scala 81:58]
  wire [1:0] pte_ppn2 = _in_req_bits_T ? tlb_io_rpte_ppn2 : ptw_pte_reg_ppn2; // @[CachePortProxy.scala 117:18]
  wire [1:0] level = _in_req_bits_T ? tlb_io_rlevel : ptw_level; // @[CachePortProxy.scala 118:18]
  wire  _tlb_io_wen_T_1 = ~page_fault; // @[CachePortProxy.scala 121:50]
  wire  _tlb_io_wen_T_2 = _T_25 & ~page_fault; // @[CachePortProxy.scala 121:47]
  wire [8:0] paddr_ppn0 = level > 2'h0 ? in_vaddr_vpn0 : pte_ppn0; // @[CachePortProxy.scala 163:22]
  wire [8:0] paddr_ppn1 = level > 2'h1 ? in_vaddr_vpn1 : pte_ppn1; // @[CachePortProxy.scala 164:22]
  wire [31:0] _io_out_req_bits_addr_T = {pte_ppn2,paddr_ppn1,paddr_ppn0,in_vaddr_offset}; // @[CachePortProxy.scala 173:43]
  wire [38:0] _io_out_req_bits_addr_WIRE = {{7'd0}, _io_out_req_bits_addr_T}; // @[CachePortProxy.scala 173:{43,43}]
  wire  _page_fault_reg_T_7 = page_fault & _GEN_7 & (_in_req_bits_T & tlb_io_hit & _T_1 | _T_25); // @[CachePortProxy.scala 178:26]
  reg  page_fault_reg; // @[Utils.scala 36:20]
  wire  _GEN_51 = _page_fault_reg_T_7 | page_fault_reg; // @[Utils.scala 41:19 36:20 41:23]
  TLB tlb ( // @[CachePortProxy.scala 28:19]
    .clock(tlb_clock),
    .reset(tlb_reset),
    .io_sfence_vma(tlb_io_sfence_vma),
    .io_vaddr_vpn2(tlb_io_vaddr_vpn2),
    .io_vaddr_vpn1(tlb_io_vaddr_vpn1),
    .io_vaddr_vpn0(tlb_io_vaddr_vpn0),
    .io_rpte_ppn2(tlb_io_rpte_ppn2),
    .io_rpte_ppn1(tlb_io_rpte_ppn1),
    .io_rpte_ppn0(tlb_io_rpte_ppn0),
    .io_rpte_flag_d(tlb_io_rpte_flag_d),
    .io_rpte_flag_a(tlb_io_rpte_flag_a),
    .io_rpte_flag_u(tlb_io_rpte_flag_u),
    .io_rpte_flag_x(tlb_io_rpte_flag_x),
    .io_rpte_flag_w(tlb_io_rpte_flag_w),
    .io_rpte_flag_r(tlb_io_rpte_flag_r),
    .io_rpte_flag_v(tlb_io_rpte_flag_v),
    .io_rlevel(tlb_io_rlevel),
    .io_hit(tlb_io_hit),
    .io_wen(tlb_io_wen),
    .io_wvaddr_vpn2(tlb_io_wvaddr_vpn2),
    .io_wvaddr_vpn1(tlb_io_wvaddr_vpn1),
    .io_wvaddr_vpn0(tlb_io_wvaddr_vpn0),
    .io_wpte_ppn2(tlb_io_wpte_ppn2),
    .io_wpte_ppn1(tlb_io_wpte_ppn1),
    .io_wpte_ppn0(tlb_io_wpte_ppn0),
    .io_wpte_flag_d(tlb_io_wpte_flag_d),
    .io_wpte_flag_a(tlb_io_wpte_flag_a),
    .io_wpte_flag_g(tlb_io_wpte_flag_g),
    .io_wpte_flag_u(tlb_io_wpte_flag_u),
    .io_wpte_flag_x(tlb_io_wpte_flag_x),
    .io_wpte_flag_w(tlb_io_wpte_flag_w),
    .io_wpte_flag_r(tlb_io_wpte_flag_r),
    .io_wpte_flag_v(tlb_io_wpte_flag_v),
    .io_wlevel(tlb_io_wlevel),
    .io_satp_asid(tlb_io_satp_asid)
  );
  assign io_in_req_ready = _in_req_bits_T & (io_out_req_ready | access_fault | _GEN_7 & (_T_2 | page_fault)); // @[CachePortProxy.scala 168:41]
  assign io_in_resp_valid = io_out_resp_valid | io_in_resp_bits_page_fault | io_in_resp_bits_access_fault; // @[CachePortProxy.scala 185:83]
  assign io_in_resp_bits_rdata = io_out_resp_bits_rdata; // @[CachePortProxy.scala 181:32]
  assign io_in_resp_bits_page_fault = page_fault_reg; // @[CachePortProxy.scala 182:32]
  assign io_in_resp_bits_access_fault = state == 3'h4; // @[CachePortProxy.scala 183:42]
  assign io_out_req_valid = _in_req_bits_T & (tlb_io_hit & _tlb_io_wen_T_1 | _access_fault_T_3 & ~access_fault) &
    io_in_req_valid | _tlb_io_wen_T_2; // @[CachePortProxy.scala 169:126]
  assign io_out_req_bits_addr = _GEN_7 ? _io_out_req_bits_addr_WIRE : _GEN_0; // @[CachePortProxy.scala 172:16 171:19 173:26]
  assign io_out_resp_ready = io_in_resp_ready; // @[CachePortProxy.scala 186:32]
  assign io_ptw_req_valid = state == 3'h1; // @[CachePortProxy.scala 113:31]
  assign io_ptw_req_bits_addr = {{7'd0}, _io_ptw_req_bits_addr_T_5}; // @[CachePortProxy.scala 104:24]
  assign io_ptw_resp_ready = state == 3'h2; // @[CachePortProxy.scala 114:31]
  assign tlb_clock = clock;
  assign tlb_reset = reset;
  assign tlb_io_sfence_vma = io_sfence_vma; // @[CachePortProxy.scala 31:21]
  assign tlb_io_vaddr_vpn2 = io_in_req_bits_addr[38:30]; // @[CachePortProxy.scala 32:52]
  assign tlb_io_vaddr_vpn1 = io_in_req_bits_addr[29:21]; // @[CachePortProxy.scala 32:52]
  assign tlb_io_vaddr_vpn0 = io_in_req_bits_addr[20:12]; // @[CachePortProxy.scala 32:52]
  assign tlb_io_wen = _T_25 & ~page_fault; // @[CachePortProxy.scala 121:47]
  assign tlb_io_wvaddr_vpn2 = _GEN_0[38:30]; // @[CachePortProxy.scala 25:46]
  assign tlb_io_wvaddr_vpn1 = _GEN_0[29:21]; // @[CachePortProxy.scala 25:46]
  assign tlb_io_wvaddr_vpn0 = _GEN_0[20:12]; // @[CachePortProxy.scala 25:46]
  assign tlb_io_wpte_ppn2 = ptw_pte_reg_ppn2; // @[CachePortProxy.scala 123:17]
  assign tlb_io_wpte_ppn1 = ptw_pte_reg_ppn1; // @[CachePortProxy.scala 123:17]
  assign tlb_io_wpte_ppn0 = ptw_pte_reg_ppn0; // @[CachePortProxy.scala 123:17]
  assign tlb_io_wpte_flag_d = ptw_pte_reg_flag_d; // @[CachePortProxy.scala 123:17]
  assign tlb_io_wpte_flag_a = ptw_pte_reg_flag_a; // @[CachePortProxy.scala 123:17]
  assign tlb_io_wpte_flag_g = ptw_pte_reg_flag_g; // @[CachePortProxy.scala 123:17]
  assign tlb_io_wpte_flag_u = ptw_pte_reg_flag_u; // @[CachePortProxy.scala 123:17]
  assign tlb_io_wpte_flag_x = ptw_pte_reg_flag_x; // @[CachePortProxy.scala 123:17]
  assign tlb_io_wpte_flag_w = ptw_pte_reg_flag_w; // @[CachePortProxy.scala 123:17]
  assign tlb_io_wpte_flag_r = ptw_pte_reg_flag_r; // @[CachePortProxy.scala 123:17]
  assign tlb_io_wpte_flag_v = ptw_pte_reg_flag_v; // @[CachePortProxy.scala 123:17]
  assign tlb_io_wlevel = ptw_level; // @[CachePortProxy.scala 124:17]
  assign tlb_io_satp_asid = io_satp_asid; // @[CachePortProxy.scala 30:21]
  always @(posedge clock) begin
    if (reset) begin // @[CachePortProxy.scala 21:93]
      state <= 3'h0; // @[CachePortProxy.scala 21:93]
    end else if (3'h0 == state) begin // @[CachePortProxy.scala 52:17]
      if (io_in_req_valid) begin // @[CachePortProxy.scala 59:29]
        if (_access_fault_T_3 & access_fault) begin // @[CachePortProxy.scala 60:39]
          state <= 3'h4; // @[CachePortProxy.scala 61:17]
        end else begin
          state <= _GEN_21;
        end
      end else begin
        state <= _GEN_21;
      end
    end else if (3'h1 == state) begin // @[CachePortProxy.scala 52:17]
      if (_T_7) begin // @[CachePortProxy.scala 67:29]
        state <= 3'h2; // @[CachePortProxy.scala 68:15]
      end
    end else if (3'h2 == state) begin // @[CachePortProxy.scala 52:17]
      state <= _GEN_27;
    end else begin
      state <= _GEN_32;
    end
    if (reset) begin // @[Reg.scala 35:20]
      in_req_bits_r_addr <= 39'h0; // @[Reg.scala 35:20]
    end else if (_in_req_bits_T) begin // @[Reg.scala 36:18]
      in_req_bits_r_addr <= io_in_req_bits_addr; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      atp_en_r <= 1'h0; // @[Reg.scala 35:20]
    end else if (_in_req_bits_T) begin // @[Reg.scala 36:18]
      atp_en_r <= _atp_en_T_1; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[CachePortProxy.scala 46:29]
      ptw_level <= 2'h0; // @[CachePortProxy.scala 46:29]
    end else if (3'h0 == state) begin // @[CachePortProxy.scala 52:17]
      ptw_level <= 2'h2; // @[CachePortProxy.scala 64:17]
    end else if (!(3'h1 == state)) begin // @[CachePortProxy.scala 52:17]
      if (3'h2 == state) begin // @[CachePortProxy.scala 52:17]
        ptw_level <= _GEN_28;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      ptw_pte_reg_ppn2 <= 2'h0; // @[Reg.scala 35:20]
    end else if (_ptw_pte_reg_T) begin // @[Reg.scala 36:18]
      ptw_pte_reg_ppn2 <= ptw_pte_ppn2; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ptw_pte_reg_ppn1 <= 9'h0; // @[Reg.scala 35:20]
    end else if (_ptw_pte_reg_T) begin // @[Reg.scala 36:18]
      ptw_pte_reg_ppn1 <= ptw_pte_ppn1; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ptw_pte_reg_ppn0 <= 9'h0; // @[Reg.scala 35:20]
    end else if (_ptw_pte_reg_T) begin // @[Reg.scala 36:18]
      ptw_pte_reg_ppn0 <= ptw_pte_ppn0; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ptw_pte_reg_flag_d <= 1'h0; // @[Reg.scala 35:20]
    end else if (_ptw_pte_reg_T) begin // @[Reg.scala 36:18]
      ptw_pte_reg_flag_d <= ptw_pte_flag_d; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ptw_pte_reg_flag_a <= 1'h0; // @[Reg.scala 35:20]
    end else if (_ptw_pte_reg_T) begin // @[Reg.scala 36:18]
      ptw_pte_reg_flag_a <= ptw_pte_flag_a; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ptw_pte_reg_flag_g <= 1'h0; // @[Reg.scala 35:20]
    end else if (_ptw_pte_reg_T) begin // @[Reg.scala 36:18]
      ptw_pte_reg_flag_g <= ptw_pte_flag_g; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ptw_pte_reg_flag_u <= 1'h0; // @[Reg.scala 35:20]
    end else if (_ptw_pte_reg_T) begin // @[Reg.scala 36:18]
      ptw_pte_reg_flag_u <= ptw_pte_flag_u; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ptw_pte_reg_flag_x <= 1'h0; // @[Reg.scala 35:20]
    end else if (_ptw_pte_reg_T) begin // @[Reg.scala 36:18]
      ptw_pte_reg_flag_x <= ptw_pte_flag_x; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ptw_pte_reg_flag_w <= 1'h0; // @[Reg.scala 35:20]
    end else if (_ptw_pte_reg_T) begin // @[Reg.scala 36:18]
      ptw_pte_reg_flag_w <= ptw_pte_flag_w; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ptw_pte_reg_flag_r <= 1'h0; // @[Reg.scala 35:20]
    end else if (_ptw_pte_reg_T) begin // @[Reg.scala 36:18]
      ptw_pte_reg_flag_r <= ptw_pte_flag_r; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ptw_pte_reg_flag_v <= 1'h0; // @[Reg.scala 35:20]
    end else if (_ptw_pte_reg_T) begin // @[Reg.scala 36:18]
      ptw_pte_reg_flag_v <= ptw_pte_flag_v; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      prv_r <= 2'h0; // @[Reg.scala 35:20]
    end else if (_in_req_bits_T) begin // @[Utils.scala 50:8]
      prv_r <= io_prv;
    end
    if (reset) begin // @[Utils.scala 36:20]
      page_fault_reg <= 1'h0; // @[Utils.scala 36:20]
    end else if (_T_14) begin // @[Utils.scala 42:18]
      page_fault_reg <= 1'h0; // @[Utils.scala 42:22]
    end else begin
      page_fault_reg <= _GEN_51;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {2{`RANDOM}};
  in_req_bits_r_addr = _RAND_1[38:0];
  _RAND_2 = {1{`RANDOM}};
  atp_en_r = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  ptw_level = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  ptw_pte_reg_ppn2 = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  ptw_pte_reg_ppn1 = _RAND_5[8:0];
  _RAND_6 = {1{`RANDOM}};
  ptw_pte_reg_ppn0 = _RAND_6[8:0];
  _RAND_7 = {1{`RANDOM}};
  ptw_pte_reg_flag_d = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  ptw_pte_reg_flag_a = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  ptw_pte_reg_flag_g = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  ptw_pte_reg_flag_u = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  ptw_pte_reg_flag_x = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  ptw_pte_reg_flag_w = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  ptw_pte_reg_flag_r = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  ptw_pte_reg_flag_v = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  prv_r = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  page_fault_reg = _RAND_16[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_2(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [63:0] io_enq_bits_pc,
  input  [31:0] io_enq_bits_instr,
  input         io_enq_bits_page_fault,
  input         io_enq_bits_access_fault,
  input  [63:0] io_enq_bits_bp_npc,
  input         io_deq_ready,
  output        io_deq_valid,
  output [63:0] io_deq_bits_pc,
  output [31:0] io_deq_bits_instr,
  output        io_deq_bits_page_fault,
  output        io_deq_bits_access_fault,
  output [63:0] io_deq_bits_bp_npc,
  input         io_flush
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] ram_pc [0:3]; // @[Decoupled.scala 273:95]
  wire  ram_pc_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire [1:0] ram_pc_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [63:0] ram_pc_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [63:0] ram_pc_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_pc_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_pc_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_pc_MPORT_en; // @[Decoupled.scala 273:95]
  reg [31:0] ram_instr [0:3]; // @[Decoupled.scala 273:95]
  wire  ram_instr_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire [1:0] ram_instr_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [31:0] ram_instr_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [31:0] ram_instr_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_instr_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_instr_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_instr_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_page_fault [0:3]; // @[Decoupled.scala 273:95]
  wire  ram_page_fault_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire [1:0] ram_page_fault_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_page_fault_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_page_fault_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_page_fault_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_page_fault_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_page_fault_MPORT_en; // @[Decoupled.scala 273:95]
  reg  ram_access_fault [0:3]; // @[Decoupled.scala 273:95]
  wire  ram_access_fault_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire [1:0] ram_access_fault_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_access_fault_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire  ram_access_fault_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_access_fault_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_access_fault_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_access_fault_MPORT_en; // @[Decoupled.scala 273:95]
  reg [63:0] ram_bp_npc [0:3]; // @[Decoupled.scala 273:95]
  wire  ram_bp_npc_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire [1:0] ram_bp_npc_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [63:0] ram_bp_npc_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [63:0] ram_bp_npc_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_bp_npc_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_bp_npc_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_bp_npc_MPORT_en; // @[Decoupled.scala 273:95]
  reg [1:0] enq_ptr_value; // @[Counter.scala 61:40]
  reg [1:0] deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _value_T_1 = enq_ptr_value + 2'h1; // @[Counter.scala 77:24]
  wire [1:0] _value_T_3 = deq_ptr_value + 2'h1; // @[Counter.scala 77:24]
  assign ram_pc_io_deq_bits_MPORT_en = 1'h1;
  assign ram_pc_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_pc_io_deq_bits_MPORT_data = ram_pc[ram_pc_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_pc_MPORT_data = io_enq_bits_pc;
  assign ram_pc_MPORT_addr = enq_ptr_value;
  assign ram_pc_MPORT_mask = 1'h1;
  assign ram_pc_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_instr_io_deq_bits_MPORT_en = 1'h1;
  assign ram_instr_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_instr_io_deq_bits_MPORT_data = ram_instr[ram_instr_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_instr_MPORT_data = io_enq_bits_instr;
  assign ram_instr_MPORT_addr = enq_ptr_value;
  assign ram_instr_MPORT_mask = 1'h1;
  assign ram_instr_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_page_fault_io_deq_bits_MPORT_en = 1'h1;
  assign ram_page_fault_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_page_fault_io_deq_bits_MPORT_data = ram_page_fault[ram_page_fault_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_page_fault_MPORT_data = io_enq_bits_page_fault;
  assign ram_page_fault_MPORT_addr = enq_ptr_value;
  assign ram_page_fault_MPORT_mask = 1'h1;
  assign ram_page_fault_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_access_fault_io_deq_bits_MPORT_en = 1'h1;
  assign ram_access_fault_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_access_fault_io_deq_bits_MPORT_data = ram_access_fault[ram_access_fault_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_access_fault_MPORT_data = io_enq_bits_access_fault;
  assign ram_access_fault_MPORT_addr = enq_ptr_value;
  assign ram_access_fault_MPORT_mask = 1'h1;
  assign ram_access_fault_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_bp_npc_io_deq_bits_MPORT_en = 1'h1;
  assign ram_bp_npc_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_bp_npc_io_deq_bits_MPORT_data = ram_bp_npc[ram_bp_npc_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_bp_npc_MPORT_data = io_enq_bits_bp_npc;
  assign ram_bp_npc_MPORT_addr = enq_ptr_value;
  assign ram_bp_npc_MPORT_mask = 1'h1;
  assign ram_bp_npc_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = io_deq_ready | ~full; // @[Decoupled.scala 303:16 323:{24,39}]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits_pc = ram_pc_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_instr = ram_instr_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_page_fault = ram_page_fault_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_access_fault = ram_access_fault_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  assign io_deq_bits_bp_npc = ram_bp_npc_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  always @(posedge clock) begin
    if (ram_pc_MPORT_en & ram_pc_MPORT_mask) begin
      ram_pc[ram_pc_MPORT_addr] <= ram_pc_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_instr_MPORT_en & ram_instr_MPORT_mask) begin
      ram_instr[ram_instr_MPORT_addr] <= ram_instr_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_page_fault_MPORT_en & ram_page_fault_MPORT_mask) begin
      ram_page_fault[ram_page_fault_MPORT_addr] <= ram_page_fault_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_access_fault_MPORT_en & ram_access_fault_MPORT_mask) begin
      ram_access_fault[ram_access_fault_MPORT_addr] <= ram_access_fault_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (ram_bp_npc_MPORT_en & ram_bp_npc_MPORT_mask) begin
      ram_bp_npc[ram_bp_npc_MPORT_addr] <= ram_bp_npc_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 2'h0; // @[Counter.scala 61:40]
    end else if (io_flush) begin // @[Decoupled.scala 296:15]
      enq_ptr_value <= 2'h0; // @[Counter.scala 98:11]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 2'h0; // @[Counter.scala 61:40]
    end else if (io_flush) begin // @[Decoupled.scala 296:15]
      deq_ptr_value <= 2'h0; // @[Counter.scala 98:11]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (io_flush) begin // @[Decoupled.scala 296:15]
      maybe_full <= 1'h0; // @[Decoupled.scala 299:16]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_pc[initvar] = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_instr[initvar] = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_page_fault[initvar] = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_access_fault[initvar] = _RAND_3[0:0];
  _RAND_4 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_bp_npc[initvar] = _RAND_4[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  enq_ptr_value = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  deq_ptr_value = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  maybe_full = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Decode(
  input  [63:0] io_in_pc,
  input  [31:0] io_in_instr,
  input         io_in_valid,
  input         io_in_page_fault,
  input         io_in_access_fault,
  output        io_out_valid,
  output [2:0]  io_out_exc,
  output [63:0] io_out_pc,
  output [63:0] io_out_npc,
  output [31:0] io_out_instr,
  output [2:0]  io_out_fu,
  output [3:0]  io_out_alu_op,
  output [1:0]  io_out_jmp_op,
  output [3:0]  io_out_mdu_op,
  output [4:0]  io_out_lsu_op,
  output [1:0]  io_out_mem_len,
  output [1:0]  io_out_csr_op,
  output [2:0]  io_out_sys_op,
  output [1:0]  io_out_rs1_src,
  output [1:0]  io_out_rs2_src,
  output [4:0]  io_out_rs1_index,
  output [4:0]  io_out_rs2_index,
  output [4:0]  io_out_rd_index,
  output        io_out_rd_wen,
  output [31:0] io_out_imm,
  output        io_out_dw
);
  wire [63:0] uop_npc = io_in_pc + 64'h4; // @[Decode.scala 16:29]
  wire [4:0] uop_rs1_index = io_in_instr[19:15]; // @[Decode.scala 18:25]
  wire [4:0] uop_rs2_index = io_in_instr[24:20]; // @[Decode.scala 19:25]
  wire [4:0] uop_rd_index = io_in_instr[11:7]; // @[Decode.scala 20:25]
  wire [31:0] decode_result_invInputs = ~io_in_instr; // @[pla.scala 78:21]
  wire  decode_result_andMatrixInput_0 = decode_result_invInputs[2]; // @[pla.scala 91:29]
  wire  decode_result_andMatrixInput_1 = decode_result_invInputs[5]; // @[pla.scala 91:29]
  wire [1:0] _decode_result_T = {decode_result_andMatrixInput_0,decode_result_andMatrixInput_1}; // @[Cat.scala 33:92]
  wire  _decode_result_T_1 = &_decode_result_T; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_1_1 = decode_result_invInputs[4]; // @[pla.scala 91:29]
  wire [2:0] _decode_result_T_2 = {decode_result_andMatrixInput_0,decode_result_andMatrixInput_1_1,
    decode_result_andMatrixInput_1}; // @[Cat.scala 33:92]
  wire  _decode_result_T_3 = &_decode_result_T_2; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_1_2 = decode_result_invInputs[6]; // @[pla.scala 91:29]
  wire [1:0] _decode_result_T_4 = {decode_result_andMatrixInput_0,decode_result_andMatrixInput_1_2}; // @[Cat.scala 33:92]
  wire  _decode_result_T_5 = &_decode_result_T_4; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_0_3 = io_in_instr[0]; // @[pla.scala 90:45]
  wire  decode_result_andMatrixInput_1_3 = io_in_instr[1]; // @[pla.scala 90:45]
  wire  decode_result_andMatrixInput_3 = decode_result_invInputs[3]; // @[pla.scala 91:29]
  wire  decode_result_andMatrixInput_6 = decode_result_invInputs[12]; // @[pla.scala 91:29]
  wire [6:0] _decode_result_T_6 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3,decode_result_andMatrixInput_1,
    decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_6}; // @[Cat.scala 33:92]
  wire  _decode_result_T_7 = &_decode_result_T_6; // @[pla.scala 98:74]
  wire [7:0] _decode_result_T_8 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3,decode_result_andMatrixInput_1_1,
    decode_result_andMatrixInput_1,decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_6}; // @[Cat.scala 33:92]
  wire  _decode_result_T_9 = &_decode_result_T_8; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_7_1 = decode_result_invInputs[13]; // @[pla.scala 91:29]
  wire [7:0] _decode_result_T_10 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3,decode_result_andMatrixInput_1_1,
    decode_result_andMatrixInput_1,decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_7_1}; // @[Cat.scala 33:92]
  wire  _decode_result_T_11 = &_decode_result_T_10; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_6_3 = decode_result_invInputs[14]; // @[pla.scala 91:29]
  wire [6:0] _decode_result_T_12 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3,decode_result_andMatrixInput_1_1,
    decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_6_3}; // @[Cat.scala 33:92]
  wire  _decode_result_T_13 = &_decode_result_T_12; // @[pla.scala 98:74]
  wire [7:0] _decode_result_T_14 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3,decode_result_andMatrixInput_1_1,
    decode_result_andMatrixInput_1,decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_6_3}; // @[Cat.scala 33:92]
  wire  _decode_result_T_15 = &_decode_result_T_14; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_8 = decode_result_invInputs[25]; // @[pla.scala 91:29]
  wire  decode_result_andMatrixInput_9 = decode_result_invInputs[26]; // @[pla.scala 91:29]
  wire  decode_result_andMatrixInput_10 = decode_result_invInputs[27]; // @[pla.scala 91:29]
  wire  decode_result_andMatrixInput_11 = decode_result_invInputs[28]; // @[pla.scala 91:29]
  wire  decode_result_andMatrixInput_12 = decode_result_invInputs[29]; // @[pla.scala 91:29]
  wire  decode_result_andMatrixInput_13 = decode_result_invInputs[31]; // @[pla.scala 91:29]
  wire [6:0] decode_result_lo_5 = {decode_result_andMatrixInput_6_3,decode_result_andMatrixInput_8,
    decode_result_andMatrixInput_9,decode_result_andMatrixInput_10,decode_result_andMatrixInput_11,
    decode_result_andMatrixInput_12,decode_result_andMatrixInput_13}; // @[Cat.scala 33:92]
  wire [13:0] _decode_result_T_16 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3,decode_result_andMatrixInput_1_2,
    decode_result_andMatrixInput_6,decode_result_andMatrixInput_7_1,decode_result_lo_5}; // @[Cat.scala 33:92]
  wire  _decode_result_T_17 = &_decode_result_T_16; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_0_9 = io_in_instr[2]; // @[pla.scala 90:45]
  wire [2:0] _decode_result_T_18 = {decode_result_andMatrixInput_0_9,decode_result_andMatrixInput_3,
    decode_result_andMatrixInput_1_1}; // @[Cat.scala 33:92]
  wire  _decode_result_T_19 = &_decode_result_T_18; // @[pla.scala 98:74]
  wire [2:0] _decode_result_T_20 = {decode_result_andMatrixInput_0_9,decode_result_andMatrixInput_3,
    decode_result_andMatrixInput_1}; // @[Cat.scala 33:92]
  wire  _decode_result_T_21 = &_decode_result_T_20; // @[pla.scala 98:74]
  wire [2:0] _decode_result_T_22 = {decode_result_andMatrixInput_0_9,decode_result_andMatrixInput_1_1,
    decode_result_andMatrixInput_1}; // @[Cat.scala 33:92]
  wire  _decode_result_T_23 = &_decode_result_T_22; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_1_12 = io_in_instr[3]; // @[pla.scala 90:45]
  wire [1:0] _decode_result_T_24 = {decode_result_andMatrixInput_0,decode_result_andMatrixInput_1_12}; // @[Cat.scala 33:92]
  wire  _decode_result_T_25 = &_decode_result_T_24; // @[pla.scala 98:74]
  wire [8:0] _decode_result_T_26 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0_9,decode_result_andMatrixInput_1_12,decode_result_andMatrixInput_1_1,
    decode_result_andMatrixInput_1,decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_7_1,
    decode_result_andMatrixInput_6_3}; // @[Cat.scala 33:92]
  wire  _decode_result_T_27 = &_decode_result_T_26; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_3_7 = io_in_instr[4]; // @[pla.scala 90:45]
  wire [8:0] _decode_result_T_28 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3_7,decode_result_andMatrixInput_1,
    decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_6,decode_result_andMatrixInput_7_1,
    decode_result_andMatrixInput_6_3}; // @[Cat.scala 33:92]
  wire  _decode_result_T_29 = &_decode_result_T_28; // @[pla.scala 98:74]
  wire [13:0] _decode_result_T_30 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3_7,decode_result_andMatrixInput_1_2,
    decode_result_andMatrixInput_6,decode_result_andMatrixInput_7_1,decode_result_lo_5}; // @[Cat.scala 33:92]
  wire  _decode_result_T_31 = &_decode_result_T_30; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_9_2 = decode_result_invInputs[30]; // @[pla.scala 91:29]
  wire [4:0] decode_result_lo_9 = {decode_result_andMatrixInput_10,decode_result_andMatrixInput_11,
    decode_result_andMatrixInput_12,decode_result_andMatrixInput_9_2,decode_result_andMatrixInput_13}; // @[Cat.scala 33:92]
  wire [10:0] _decode_result_T_32 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_3,decode_result_andMatrixInput_3_7,decode_result_andMatrixInput_1_2,
    decode_result_andMatrixInput_9,decode_result_lo_9}; // @[Cat.scala 33:92]
  wire  _decode_result_T_33 = &_decode_result_T_32; // @[pla.scala 98:74]
  wire [1:0] _decode_result_T_34 = {decode_result_andMatrixInput_0_9,decode_result_andMatrixInput_3_7}; // @[Cat.scala 33:92]
  wire  _decode_result_T_35 = &_decode_result_T_34; // @[pla.scala 98:74]
  wire [5:0] _decode_result_T_36 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0_9,decode_result_andMatrixInput_3,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_1_2}; // @[Cat.scala 33:92]
  wire  _decode_result_T_37 = &_decode_result_T_36; // @[pla.scala 98:74]
  wire [9:0] _decode_result_T_38 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_1_12,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_1,decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_6,
    decode_result_andMatrixInput_7_1,decode_result_andMatrixInput_6_3}; // @[Cat.scala 33:92]
  wire  _decode_result_T_39 = &_decode_result_T_38; // @[pla.scala 98:74]
  wire [14:0] _decode_result_T_40 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_1_12,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_6,decode_result_andMatrixInput_7_1,decode_result_lo_5}
    ; // @[Cat.scala 33:92]
  wire  _decode_result_T_41 = &_decode_result_T_40; // @[pla.scala 98:74]
  wire [6:0] decode_result_lo_13 = {decode_result_andMatrixInput_6_3,decode_result_andMatrixInput_9,
    decode_result_andMatrixInput_10,decode_result_andMatrixInput_11,decode_result_andMatrixInput_12,
    decode_result_andMatrixInput_9_2,decode_result_andMatrixInput_13}; // @[Cat.scala 33:92]
  wire [14:0] _decode_result_T_42 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_1_12,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_6,decode_result_andMatrixInput_7_1,decode_result_lo_13
    }; // @[Cat.scala 33:92]
  wire  _decode_result_T_43 = &_decode_result_T_42; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_2_18 = io_in_instr[5]; // @[pla.scala 90:45]
  wire [3:0] _decode_result_T_44 = {decode_result_andMatrixInput_0,decode_result_andMatrixInput_1_1,
    decode_result_andMatrixInput_2_18,decode_result_andMatrixInput_1_2}; // @[Cat.scala 33:92]
  wire  _decode_result_T_45 = &_decode_result_T_44; // @[pla.scala 98:74]
  wire [4:0] _decode_result_T_46 = {decode_result_andMatrixInput_0_9,decode_result_andMatrixInput_1_12,
    decode_result_andMatrixInput_2_18,decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_11}; // @[Cat.scala 33:92]
  wire  _decode_result_T_47 = &_decode_result_T_46; // @[pla.scala 98:74]
  wire [8:0] _decode_result_T_48 = {decode_result_andMatrixInput_0_9,decode_result_andMatrixInput_1_12,
    decode_result_andMatrixInput_2_18,decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_10,
    decode_result_andMatrixInput_11,decode_result_andMatrixInput_12,decode_result_andMatrixInput_9_2,
    decode_result_andMatrixInput_13}; // @[Cat.scala 33:92]
  wire  _decode_result_T_49 = &_decode_result_T_48; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_3_17 = io_in_instr[6]; // @[pla.scala 90:45]
  wire [4:0] _decode_result_T_50 = {decode_result_andMatrixInput_0,decode_result_andMatrixInput_3,
    decode_result_andMatrixInput_1_1,decode_result_andMatrixInput_3_17,decode_result_andMatrixInput_6_3}; // @[Cat.scala 33:92]
  wire  _decode_result_T_51 = &_decode_result_T_50; // @[pla.scala 98:74]
  wire [2:0] _decode_result_T_52 = {decode_result_andMatrixInput_0_9,decode_result_andMatrixInput_1_12,
    decode_result_andMatrixInput_3_17}; // @[Cat.scala 33:92]
  wire  _decode_result_T_53 = &_decode_result_T_52; // @[pla.scala 98:74]
  wire [1:0] _decode_result_T_54 = {decode_result_andMatrixInput_3_7,decode_result_andMatrixInput_3_17}; // @[Cat.scala 33:92]
  wire  _decode_result_T_55 = &_decode_result_T_54; // @[pla.scala 98:74]
  wire [7:0] _decode_result_T_56 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3,decode_result_andMatrixInput_1_1,
    decode_result_andMatrixInput_2_18,decode_result_andMatrixInput_3_17,decode_result_andMatrixInput_7_1}; // @[Cat.scala 33:92]
  wire  _decode_result_T_57 = &_decode_result_T_56; // @[pla.scala 98:74]
  wire [8:0] _decode_result_T_58 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_3,decode_result_andMatrixInput_1_1,decode_result_andMatrixInput_2_18,
    decode_result_andMatrixInput_3_17,decode_result_andMatrixInput_6,decode_result_andMatrixInput_7_1,
    decode_result_andMatrixInput_6_3}; // @[Cat.scala 33:92]
  wire  _decode_result_T_59 = &_decode_result_T_58; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_5_17 = decode_result_invInputs[7]; // @[pla.scala 91:29]
  wire  decode_result_andMatrixInput_6_16 = decode_result_invInputs[8]; // @[pla.scala 91:29]
  wire  decode_result_andMatrixInput_7_14 = decode_result_invInputs[9]; // @[pla.scala 91:29]
  wire  decode_result_andMatrixInput_8_10 = decode_result_invInputs[10]; // @[pla.scala 91:29]
  wire  decode_result_andMatrixInput_9_6 = decode_result_invInputs[11]; // @[pla.scala 91:29]
  wire  decode_result_andMatrixInput_13_4 = decode_result_invInputs[15]; // @[pla.scala 91:29]
  wire  decode_result_andMatrixInput_14_2 = decode_result_invInputs[16]; // @[pla.scala 91:29]
  wire  decode_result_andMatrixInput_15 = decode_result_invInputs[17]; // @[pla.scala 91:29]
  wire  decode_result_andMatrixInput_16 = decode_result_invInputs[18]; // @[pla.scala 91:29]
  wire  decode_result_andMatrixInput_17 = decode_result_invInputs[19]; // @[pla.scala 91:29]
  wire  decode_result_andMatrixInput_18 = decode_result_invInputs[20]; // @[pla.scala 91:29]
  wire  decode_result_andMatrixInput_19 = decode_result_invInputs[21]; // @[pla.scala 91:29]
  wire  decode_result_andMatrixInput_20 = decode_result_invInputs[22]; // @[pla.scala 91:29]
  wire  decode_result_andMatrixInput_21 = decode_result_invInputs[23]; // @[pla.scala 91:29]
  wire  decode_result_andMatrixInput_22 = decode_result_invInputs[24]; // @[pla.scala 91:29]
  wire [6:0] decode_result_lo_lo_14 = {decode_result_andMatrixInput_8,decode_result_andMatrixInput_9,
    decode_result_andMatrixInput_10,decode_result_andMatrixInput_11,decode_result_andMatrixInput_12,
    decode_result_andMatrixInput_9_2,decode_result_andMatrixInput_13}; // @[Cat.scala 33:92]
  wire [14:0] decode_result_lo_20 = {decode_result_andMatrixInput_15,decode_result_andMatrixInput_16,
    decode_result_andMatrixInput_17,decode_result_andMatrixInput_18,decode_result_andMatrixInput_19,
    decode_result_andMatrixInput_20,decode_result_andMatrixInput_21,decode_result_andMatrixInput_22,
    decode_result_lo_lo_14}; // @[Cat.scala 33:92]
  wire [6:0] decode_result_hi_lo_16 = {decode_result_andMatrixInput_8_10,decode_result_andMatrixInput_9_6,
    decode_result_andMatrixInput_6,decode_result_andMatrixInput_7_1,decode_result_andMatrixInput_6_3,
    decode_result_andMatrixInput_13_4,decode_result_andMatrixInput_14_2}; // @[Cat.scala 33:92]
  wire [29:0] _decode_result_T_60 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_1_1,decode_result_andMatrixInput_2_18,decode_result_andMatrixInput_3_17,
    decode_result_andMatrixInput_5_17,decode_result_andMatrixInput_6_16,decode_result_andMatrixInput_7_14,
    decode_result_hi_lo_16,decode_result_lo_20}; // @[Cat.scala 33:92]
  wire  _decode_result_T_61 = &_decode_result_T_60; // @[pla.scala 98:74]
  wire [8:0] _decode_result_T_62 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0_9,decode_result_andMatrixInput_1_1,decode_result_andMatrixInput_2_18,
    decode_result_andMatrixInput_3_17,decode_result_andMatrixInput_6,decode_result_andMatrixInput_7_1,
    decode_result_andMatrixInput_6_3}; // @[Cat.scala 33:92]
  wire  _decode_result_T_63 = &_decode_result_T_62; // @[pla.scala 98:74]
  wire [6:0] _decode_result_T_64 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0_9,decode_result_andMatrixInput_1_12,decode_result_andMatrixInput_1_1,
    decode_result_andMatrixInput_2_18,decode_result_andMatrixInput_3_17}; // @[Cat.scala 33:92]
  wire  _decode_result_T_65 = &_decode_result_T_64; // @[pla.scala 98:74]
  wire [14:0] decode_result_lo_23 = {decode_result_andMatrixInput_14_2,decode_result_andMatrixInput_15,
    decode_result_andMatrixInput_16,decode_result_andMatrixInput_17,decode_result_andMatrixInput_19,
    decode_result_andMatrixInput_20,decode_result_andMatrixInput_21,decode_result_andMatrixInput_22,
    decode_result_lo_lo_14}; // @[Cat.scala 33:92]
  wire [7:0] decode_result_hi_lo_19 = {decode_result_andMatrixInput_6_16,decode_result_andMatrixInput_7_14,
    decode_result_andMatrixInput_8_10,decode_result_andMatrixInput_9_6,decode_result_andMatrixInput_6,
    decode_result_andMatrixInput_7_1,decode_result_andMatrixInput_6_3,decode_result_andMatrixInput_13_4}; // @[Cat.scala 33:92]
  wire [30:0] _decode_result_T_66 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_2_18,decode_result_andMatrixInput_3_17,decode_result_andMatrixInput_5_17,
    decode_result_hi_lo_19,decode_result_lo_23}; // @[Cat.scala 33:92]
  wire  _decode_result_T_67 = &_decode_result_T_66; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_0_34 = io_in_instr[12]; // @[pla.scala 90:45]
  wire  _decode_result_T_68 = &decode_result_andMatrixInput_0_34; // @[pla.scala 98:74]
  wire [3:0] _decode_result_T_69 = {decode_result_andMatrixInput_0_9,decode_result_andMatrixInput_1_12,
    decode_result_andMatrixInput_1,decode_result_andMatrixInput_0_34}; // @[Cat.scala 33:92]
  wire  _decode_result_T_70 = &_decode_result_T_69; // @[pla.scala 98:74]
  wire [3:0] _decode_result_T_71 = {decode_result_andMatrixInput_0,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_0_34,decode_result_andMatrixInput_7_1}; // @[Cat.scala 33:92]
  wire  _decode_result_T_72 = &_decode_result_T_71; // @[pla.scala 98:74]
  wire [13:0] _decode_result_T_73 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3_7,decode_result_andMatrixInput_1_2,
    decode_result_andMatrixInput_0_34,decode_result_andMatrixInput_7_1,decode_result_lo_lo_14}; // @[Cat.scala 33:92]
  wire  _decode_result_T_74 = &_decode_result_T_73; // @[pla.scala 98:74]
  wire [14:0] _decode_result_T_75 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_1_12,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_0_34,decode_result_andMatrixInput_7_1,
    decode_result_lo_lo_14}; // @[Cat.scala 33:92]
  wire  _decode_result_T_76 = &_decode_result_T_75; // @[pla.scala 98:74]
  wire [2:0] _decode_result_T_77 = {decode_result_andMatrixInput_0,decode_result_andMatrixInput_3_17,
    decode_result_andMatrixInput_0_34}; // @[Cat.scala 33:92]
  wire  _decode_result_T_78 = &_decode_result_T_77; // @[pla.scala 98:74]
  wire [2:0] _decode_result_T_79 = {decode_result_andMatrixInput_3_7,decode_result_andMatrixInput_3_17,
    decode_result_andMatrixInput_0_34}; // @[Cat.scala 33:92]
  wire  _decode_result_T_80 = &_decode_result_T_79; // @[pla.scala 98:74]
  wire [7:0] _decode_result_T_81 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3,decode_result_andMatrixInput_2_18,
    decode_result_andMatrixInput_3_17,decode_result_andMatrixInput_0_34,decode_result_andMatrixInput_7_1}; // @[Cat.scala 33:92]
  wire  _decode_result_T_82 = &_decode_result_T_81; // @[pla.scala 98:74]
  wire [7:0] _decode_result_T_83 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_2_18,decode_result_andMatrixInput_3_17,decode_result_andMatrixInput_0_34}; // @[Cat.scala 33:92]
  wire  _decode_result_T_84 = &_decode_result_T_83; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_1_42 = io_in_instr[13]; // @[pla.scala 90:45]
  wire [1:0] _decode_result_T_85 = {decode_result_andMatrixInput_0,decode_result_andMatrixInput_1_42}; // @[Cat.scala 33:92]
  wire  _decode_result_T_86 = &_decode_result_T_85; // @[pla.scala 98:74]
  wire [3:0] _decode_result_T_87 = {decode_result_andMatrixInput_0,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_1_42,decode_result_andMatrixInput_6_3}; // @[Cat.scala 33:92]
  wire  _decode_result_T_88 = &_decode_result_T_87; // @[pla.scala 98:74]
  wire [6:0] _decode_result_T_89 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_3,decode_result_andMatrixInput_3_7,decode_result_andMatrixInput_1,
    decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_1_42}; // @[Cat.scala 33:92]
  wire  _decode_result_T_90 = &_decode_result_T_89; // @[pla.scala 98:74]
  wire [9:0] _decode_result_T_91 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0_9,decode_result_andMatrixInput_1_12,decode_result_andMatrixInput_1_1,
    decode_result_andMatrixInput_2_18,decode_result_andMatrixInput_1_42,decode_result_andMatrixInput_6_3,
    decode_result_andMatrixInput_10,decode_result_andMatrixInput_11}; // @[Cat.scala 33:92]
  wire  _decode_result_T_92 = &_decode_result_T_91; // @[pla.scala 98:74]
  wire [4:0] decode_result_lo_33 = {decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_1_42,
    decode_result_andMatrixInput_6_3,decode_result_andMatrixInput_10,decode_result_andMatrixInput_11}; // @[Cat.scala 33:92]
  wire [10:0] _decode_result_T_93 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0_9,decode_result_andMatrixInput_1_12,decode_result_andMatrixInput_1_1,
    decode_result_andMatrixInput_2_18,decode_result_lo_33}; // @[Cat.scala 33:92]
  wire  _decode_result_T_94 = &_decode_result_T_93; // @[pla.scala 98:74]
  wire [7:0] decode_result_lo_34 = {decode_result_andMatrixInput_18,decode_result_andMatrixInput_19,
    decode_result_andMatrixInput_20,decode_result_andMatrixInput_21,decode_result_andMatrixInput_22,
    decode_result_andMatrixInput_12,decode_result_andMatrixInput_9_2,decode_result_andMatrixInput_13}; // @[Cat.scala 33:92]
  wire [15:0] _decode_result_T_95 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0_9,decode_result_andMatrixInput_1_12,decode_result_andMatrixInput_1_1,
    decode_result_andMatrixInput_2_18,decode_result_andMatrixInput_1_42,decode_result_andMatrixInput_6_3,
    decode_result_lo_34}; // @[Cat.scala 33:92]
  wire  _decode_result_T_96 = &_decode_result_T_95; // @[pla.scala 98:74]
  wire [16:0] _decode_result_T_97 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0_9,decode_result_andMatrixInput_1_12,decode_result_andMatrixInput_1_1,
    decode_result_andMatrixInput_2_18,decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_1_42,
    decode_result_andMatrixInput_6_3,decode_result_lo_34}; // @[Cat.scala 33:92]
  wire  _decode_result_T_98 = &_decode_result_T_97; // @[pla.scala 98:74]
  wire [2:0] _decode_result_T_99 = {decode_result_andMatrixInput_3_7,decode_result_andMatrixInput_3_17,
    decode_result_andMatrixInput_1_42}; // @[Cat.scala 33:92]
  wire  _decode_result_T_100 = &_decode_result_T_99; // @[pla.scala 98:74]
  wire [7:0] _decode_result_T_101 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_2_18,decode_result_andMatrixInput_3_17,decode_result_andMatrixInput_1_42}; // @[Cat.scala 33:92]
  wire  _decode_result_T_102 = &_decode_result_T_101; // @[pla.scala 98:74]
  wire [3:0] _decode_result_T_103 = {decode_result_andMatrixInput_0,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_0_34,decode_result_andMatrixInput_1_42}; // @[Cat.scala 33:92]
  wire  _decode_result_T_104 = &_decode_result_T_103; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_2_46 = io_in_instr[14]; // @[pla.scala 90:45]
  wire [2:0] _decode_result_T_105 = {decode_result_andMatrixInput_1_1,decode_result_andMatrixInput_1,
    decode_result_andMatrixInput_2_46}; // @[Cat.scala 33:92]
  wire  _decode_result_T_106 = &_decode_result_T_105; // @[pla.scala 98:74]
  wire [3:0] _decode_result_T_107 = {decode_result_andMatrixInput_0,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_6,decode_result_andMatrixInput_2_46}; // @[Cat.scala 33:92]
  wire  _decode_result_T_108 = &_decode_result_T_107; // @[pla.scala 98:74]
  wire [3:0] _decode_result_T_109 = {decode_result_andMatrixInput_0,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_2_46,decode_result_andMatrixInput_9_2}; // @[Cat.scala 33:92]
  wire  _decode_result_T_110 = &_decode_result_T_109; // @[pla.scala 98:74]
  wire [5:0] decode_result_lo_40 = {decode_result_andMatrixInput_2_46,decode_result_andMatrixInput_9,
    decode_result_andMatrixInput_10,decode_result_andMatrixInput_11,decode_result_andMatrixInput_12,
    decode_result_andMatrixInput_13}; // @[Cat.scala 33:92]
  wire [11:0] _decode_result_T_111 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_3,decode_result_andMatrixInput_3_7,decode_result_andMatrixInput_1,
    decode_result_andMatrixInput_1_2,decode_result_lo_40}; // @[Cat.scala 33:92]
  wire  _decode_result_T_112 = &_decode_result_T_111; // @[pla.scala 98:74]
  wire [3:0] _decode_result_T_113 = {decode_result_andMatrixInput_0,decode_result_andMatrixInput_1_1,
    decode_result_andMatrixInput_2_18,decode_result_andMatrixInput_2_46}; // @[Cat.scala 33:92]
  wire  _decode_result_T_114 = &_decode_result_T_113; // @[pla.scala 98:74]
  wire [2:0] _decode_result_T_115 = {decode_result_andMatrixInput_3_7,decode_result_andMatrixInput_3_17,
    decode_result_andMatrixInput_2_46}; // @[Cat.scala 33:92]
  wire  _decode_result_T_116 = &_decode_result_T_115; // @[pla.scala 98:74]
  wire [7:0] _decode_result_T_117 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3,decode_result_andMatrixInput_1_1,
    decode_result_andMatrixInput_2_18,decode_result_andMatrixInput_3_17,decode_result_andMatrixInput_2_46}; // @[Cat.scala 33:92]
  wire  _decode_result_T_118 = &_decode_result_T_117; // @[pla.scala 98:74]
  wire [3:0] _decode_result_T_119 = {decode_result_andMatrixInput_0,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_0_34,decode_result_andMatrixInput_2_46}; // @[Cat.scala 33:92]
  wire  _decode_result_T_120 = &_decode_result_T_119; // @[pla.scala 98:74]
  wire [6:0] decode_result_lo_44 = {decode_result_andMatrixInput_2_46,decode_result_andMatrixInput_8,
    decode_result_andMatrixInput_9,decode_result_andMatrixInput_10,decode_result_andMatrixInput_11,
    decode_result_andMatrixInput_12,decode_result_andMatrixInput_13}; // @[Cat.scala 33:92]
  wire [13:0] _decode_result_T_121 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3_7,decode_result_andMatrixInput_1_2,
    decode_result_andMatrixInput_0_34,decode_result_andMatrixInput_7_1,decode_result_lo_44}; // @[Cat.scala 33:92]
  wire  _decode_result_T_122 = &_decode_result_T_121; // @[pla.scala 98:74]
  wire [14:0] _decode_result_T_123 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_1_12,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_0_34,decode_result_andMatrixInput_7_1,
    decode_result_lo_44}; // @[Cat.scala 33:92]
  wire  _decode_result_T_124 = &_decode_result_T_123; // @[pla.scala 98:74]
  wire [3:0] _decode_result_T_125 = {decode_result_andMatrixInput_0,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_1_42,decode_result_andMatrixInput_2_46}; // @[Cat.scala 33:92]
  wire  _decode_result_T_126 = &_decode_result_T_125; // @[pla.scala 98:74]
  wire [3:0] _decode_result_T_127 = {decode_result_andMatrixInput_0,decode_result_andMatrixInput_2_18,
    decode_result_andMatrixInput_1_42,decode_result_andMatrixInput_2_46}; // @[Cat.scala 33:92]
  wire  _decode_result_T_128 = &_decode_result_T_127; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_20_2 = io_in_instr[20]; // @[pla.scala 90:45]
  wire [7:0] decode_result_lo_lo_30 = {decode_result_andMatrixInput_22,decode_result_andMatrixInput_8,
    decode_result_andMatrixInput_9,decode_result_andMatrixInput_10,decode_result_andMatrixInput_11,
    decode_result_andMatrixInput_12,decode_result_andMatrixInput_9_2,decode_result_andMatrixInput_13}; // @[Cat.scala 33:92]
  wire [15:0] decode_result_lo_48 = {decode_result_andMatrixInput_14_2,decode_result_andMatrixInput_15,
    decode_result_andMatrixInput_16,decode_result_andMatrixInput_17,decode_result_andMatrixInput_20_2,
    decode_result_andMatrixInput_19,decode_result_andMatrixInput_20,decode_result_andMatrixInput_21,
    decode_result_lo_lo_30}; // @[Cat.scala 33:92]
  wire [31:0] _decode_result_T_129 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_2_18,decode_result_andMatrixInput_3_17,decode_result_andMatrixInput_5_17,
    decode_result_hi_lo_19,decode_result_lo_48}; // @[Cat.scala 33:92]
  wire  _decode_result_T_130 = &_decode_result_T_129; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_4_38 = io_in_instr[21]; // @[pla.scala 90:45]
  wire [5:0] _decode_result_T_131 = {decode_result_andMatrixInput_3_7,decode_result_andMatrixInput_3_17,
    decode_result_andMatrixInput_6,decode_result_andMatrixInput_7_1,decode_result_andMatrixInput_4_38,
    decode_result_andMatrixInput_12}; // @[Cat.scala 33:92]
  wire  _decode_result_T_132 = &_decode_result_T_131; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_7_31 = io_in_instr[25]; // @[pla.scala 90:45]
  wire [6:0] decode_result_lo_50 = {decode_result_andMatrixInput_7_31,decode_result_andMatrixInput_9,
    decode_result_andMatrixInput_10,decode_result_andMatrixInput_11,decode_result_andMatrixInput_12,
    decode_result_andMatrixInput_9_2,decode_result_andMatrixInput_13}; // @[Cat.scala 33:92]
  wire [13:0] _decode_result_T_133 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_2_18,decode_result_andMatrixInput_1_2,decode_result_lo_50}; // @[Cat.scala 33:92]
  wire  _decode_result_T_134 = &_decode_result_T_133; // @[pla.scala 98:74]
  wire [14:0] _decode_result_T_135 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3_7,decode_result_andMatrixInput_2_18,
    decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_6,decode_result_andMatrixInput_7_1,decode_result_lo_50
    }; // @[Cat.scala 33:92]
  wire  _decode_result_T_136 = &_decode_result_T_135; // @[pla.scala 98:74]
  wire [4:0] _decode_result_T_137 = {decode_result_andMatrixInput_3_7,decode_result_andMatrixInput_3_17,
    decode_result_andMatrixInput_6,decode_result_andMatrixInput_7_1,decode_result_andMatrixInput_7_31}; // @[Cat.scala 33:92]
  wire  _decode_result_T_138 = &_decode_result_T_137; // @[pla.scala 98:74]
  wire [13:0] _decode_result_T_139 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3_7,decode_result_andMatrixInput_2_18,
    decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_2_46,decode_result_lo_50}; // @[Cat.scala 33:92]
  wire  _decode_result_T_140 = &_decode_result_T_139; // @[pla.scala 98:74]
  wire [14:0] _decode_result_T_141 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_1_12,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_2_18,decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_2_46,
    decode_result_lo_50}; // @[Cat.scala 33:92]
  wire  _decode_result_T_142 = &_decode_result_T_141; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_3_55 = io_in_instr[27]; // @[pla.scala 90:45]
  wire [3:0] _decode_result_T_143 = {decode_result_andMatrixInput_1_12,decode_result_andMatrixInput_2_18,
    decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_3_55}; // @[Cat.scala 33:92]
  wire  _decode_result_T_144 = &_decode_result_T_143; // @[pla.scala 98:74]
  wire [4:0] _decode_result_T_145 = {decode_result_andMatrixInput_1_12,decode_result_andMatrixInput_2_18,
    decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_3_55,decode_result_andMatrixInput_11}; // @[Cat.scala 33:92]
  wire  _decode_result_T_146 = &_decode_result_T_145; // @[pla.scala 98:74]
  wire [5:0] decode_result_lo_57 = {decode_result_andMatrixInput_1_42,decode_result_andMatrixInput_6_3,
    decode_result_andMatrixInput_3_55,decode_result_andMatrixInput_12,decode_result_andMatrixInput_9_2,
    decode_result_andMatrixInput_13}; // @[Cat.scala 33:92]
  wire [11:0] _decode_result_T_147 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0_9,decode_result_andMatrixInput_1_12,decode_result_andMatrixInput_1_1,
    decode_result_andMatrixInput_2_18,decode_result_lo_57}; // @[Cat.scala 33:92]
  wire  _decode_result_T_148 = &_decode_result_T_147; // @[pla.scala 98:74]
  wire [12:0] _decode_result_T_149 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0_9,decode_result_andMatrixInput_1_12,decode_result_andMatrixInput_1_1,
    decode_result_andMatrixInput_2_18,decode_result_andMatrixInput_1_2,decode_result_lo_57}; // @[Cat.scala 33:92]
  wire  _decode_result_T_150 = &_decode_result_T_149; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_4_47 = io_in_instr[28]; // @[pla.scala 90:45]
  wire [4:0] _decode_result_T_151 = {decode_result_andMatrixInput_1_12,decode_result_andMatrixInput_2_18,
    decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_10,decode_result_andMatrixInput_4_47}; // @[Cat.scala 33:92]
  wire  _decode_result_T_152 = &_decode_result_T_151; // @[pla.scala 98:74]
  wire [6:0] decode_result_lo_lo_37 = {decode_result_andMatrixInput_22,decode_result_andMatrixInput_8,
    decode_result_andMatrixInput_9,decode_result_andMatrixInput_10,decode_result_andMatrixInput_4_47,
    decode_result_andMatrixInput_9_2,decode_result_andMatrixInput_13}; // @[Cat.scala 33:92]
  wire [13:0] decode_result_lo_60 = {decode_result_andMatrixInput_15,decode_result_andMatrixInput_16,
    decode_result_andMatrixInput_17,decode_result_andMatrixInput_18,decode_result_andMatrixInput_4_38,
    decode_result_andMatrixInput_20,decode_result_andMatrixInput_21,decode_result_lo_lo_37}; // @[Cat.scala 33:92]
  wire [6:0] decode_result_hi_lo_41 = {decode_result_andMatrixInput_6_16,decode_result_andMatrixInput_7_14,
    decode_result_andMatrixInput_8_10,decode_result_andMatrixInput_9_6,decode_result_andMatrixInput_6_3,
    decode_result_andMatrixInput_13_4,decode_result_andMatrixInput_14_2}; // @[Cat.scala 33:92]
  wire [28:0] _decode_result_T_153 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_2_18,decode_result_andMatrixInput_3_17,decode_result_andMatrixInput_5_17,
    decode_result_hi_lo_41,decode_result_lo_60}; // @[Cat.scala 33:92]
  wire  _decode_result_T_154 = &_decode_result_T_153; // @[pla.scala 98:74]
  wire [14:0] decode_result_lo_61 = {decode_result_andMatrixInput_14_2,decode_result_andMatrixInput_15,
    decode_result_andMatrixInput_16,decode_result_andMatrixInput_17,decode_result_andMatrixInput_18,
    decode_result_andMatrixInput_4_38,decode_result_andMatrixInput_20,decode_result_andMatrixInput_21,
    decode_result_lo_lo_37}; // @[Cat.scala 33:92]
  wire [30:0] _decode_result_T_155 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_2_18,decode_result_andMatrixInput_3_17,decode_result_andMatrixInput_5_17,
    decode_result_hi_lo_19,decode_result_lo_61}; // @[Cat.scala 33:92]
  wire  _decode_result_T_156 = &_decode_result_T_155; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_20_5 = io_in_instr[22]; // @[pla.scala 90:45]
  wire [6:0] decode_result_lo_lo_39 = {decode_result_andMatrixInput_22,decode_result_andMatrixInput_9,
    decode_result_andMatrixInput_10,decode_result_andMatrixInput_4_47,decode_result_andMatrixInput_12,
    decode_result_andMatrixInput_9_2,decode_result_andMatrixInput_13}; // @[Cat.scala 33:92]
  wire [13:0] decode_result_lo_62 = {decode_result_andMatrixInput_15,decode_result_andMatrixInput_16,
    decode_result_andMatrixInput_17,decode_result_andMatrixInput_20_2,decode_result_andMatrixInput_19,
    decode_result_andMatrixInput_20_5,decode_result_andMatrixInput_21,decode_result_lo_lo_39}; // @[Cat.scala 33:92]
  wire [28:0] _decode_result_T_157 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_2_18,decode_result_andMatrixInput_3_17,decode_result_andMatrixInput_5_17,
    decode_result_hi_lo_41,decode_result_lo_62}; // @[Cat.scala 33:92]
  wire  _decode_result_T_158 = &_decode_result_T_157; // @[pla.scala 98:74]
  wire [4:0] decode_result_lo_lo_40 = {decode_result_andMatrixInput_10,decode_result_andMatrixInput_4_47,
    decode_result_andMatrixInput_12,decode_result_andMatrixInput_9_2,decode_result_andMatrixInput_13}; // @[Cat.scala 33:92]
  wire [9:0] decode_result_lo_63 = {decode_result_andMatrixInput_8_10,decode_result_andMatrixInput_9_6,
    decode_result_andMatrixInput_6_3,decode_result_andMatrixInput_7_31,decode_result_andMatrixInput_9,
    decode_result_andMatrixInput_10,decode_result_andMatrixInput_4_47,decode_result_andMatrixInput_12,
    decode_result_andMatrixInput_9_2,decode_result_andMatrixInput_13}; // @[Cat.scala 33:92]
  wire [9:0] decode_result_hi_73 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_2_18,decode_result_andMatrixInput_3_17,decode_result_andMatrixInput_5_17,
    decode_result_andMatrixInput_6_16,decode_result_andMatrixInput_7_14}; // @[Cat.scala 33:92]
  wire [19:0] _decode_result_T_159 = {decode_result_hi_73,decode_result_lo_63}; // @[Cat.scala 33:92]
  wire  _decode_result_T_160 = &_decode_result_T_159; // @[pla.scala 98:74]
  wire [10:0] decode_result_lo_64 = {decode_result_andMatrixInput_9_6,decode_result_andMatrixInput_6,
    decode_result_andMatrixInput_7_1,decode_result_andMatrixInput_6_3,decode_result_andMatrixInput_7_31,
    decode_result_andMatrixInput_9,decode_result_lo_lo_40}; // @[Cat.scala 33:92]
  wire [4:0] decode_result_hi_lo_45 = {decode_result_andMatrixInput_3_17,decode_result_andMatrixInput_5_17,
    decode_result_andMatrixInput_6_16,decode_result_andMatrixInput_7_14,decode_result_andMatrixInput_8_10}; // @[Cat.scala 33:92]
  wire [21:0] _decode_result_T_161 = {decode_result_andMatrixInput_0_3,decode_result_andMatrixInput_1_3,
    decode_result_andMatrixInput_0,decode_result_andMatrixInput_3,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_2_18,decode_result_hi_lo_45,decode_result_lo_64}; // @[Cat.scala 33:92]
  wire  _decode_result_T_162 = &_decode_result_T_161; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_3_65 = io_in_instr[29]; // @[pla.scala 90:45]
  wire [4:0] _decode_result_T_163 = {decode_result_andMatrixInput_1_12,decode_result_andMatrixInput_2_18,
    decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_3_65,decode_result_andMatrixInput_13}; // @[Cat.scala 33:92]
  wire  _decode_result_T_164 = &_decode_result_T_163; // @[pla.scala 98:74]
  wire [4:0] _decode_result_T_165 = {decode_result_andMatrixInput_3_7,decode_result_andMatrixInput_3_17,
    decode_result_andMatrixInput_6,decode_result_andMatrixInput_7_1,decode_result_andMatrixInput_3_65}; // @[Cat.scala 33:92]
  wire  _decode_result_T_166 = &_decode_result_T_165; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_3_67 = io_in_instr[30]; // @[pla.scala 90:45]
  wire [3:0] _decode_result_T_167 = {decode_result_andMatrixInput_0,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_2_18,decode_result_andMatrixInput_3_67}; // @[Cat.scala 33:92]
  wire  _decode_result_T_168 = &_decode_result_T_167; // @[pla.scala 98:74]
  wire [4:0] _decode_result_T_169 = {decode_result_andMatrixInput_0,decode_result_andMatrixInput_3_7,
    decode_result_andMatrixInput_0_34,decode_result_andMatrixInput_7_1,decode_result_andMatrixInput_3_67}; // @[Cat.scala 33:92]
  wire  _decode_result_T_170 = &_decode_result_T_169; // @[pla.scala 98:74]
  wire [5:0] _decode_result_T_171 = {decode_result_andMatrixInput_1_12,decode_result_andMatrixInput_1_2,
    decode_result_andMatrixInput_1_42,decode_result_andMatrixInput_12,decode_result_andMatrixInput_3_67,
    decode_result_andMatrixInput_13}; // @[Cat.scala 33:92]
  wire  _decode_result_T_172 = &_decode_result_T_171; // @[pla.scala 98:74]
  wire [4:0] _decode_result_T_173 = {decode_result_andMatrixInput_1_12,decode_result_andMatrixInput_2_18,
    decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_3_65,decode_result_andMatrixInput_3_67}; // @[Cat.scala 33:92]
  wire  _decode_result_T_174 = &_decode_result_T_173; // @[pla.scala 98:74]
  wire  decode_result_andMatrixInput_4_58 = io_in_instr[31]; // @[pla.scala 90:45]
  wire [4:0] _decode_result_T_175 = {decode_result_andMatrixInput_1_12,decode_result_andMatrixInput_2_18,
    decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_3_65,decode_result_andMatrixInput_4_58}; // @[Cat.scala 33:92]
  wire  _decode_result_T_176 = &_decode_result_T_175; // @[pla.scala 98:74]
  wire [4:0] _decode_result_T_177 = {decode_result_andMatrixInput_1_12,decode_result_andMatrixInput_2_18,
    decode_result_andMatrixInput_1_2,decode_result_andMatrixInput_3_67,decode_result_andMatrixInput_4_58}; // @[Cat.scala 33:92]
  wire  _decode_result_T_178 = &_decode_result_T_177; // @[pla.scala 98:74]
  wire [5:0] _decode_result_orMatrixOutputs_T = {_decode_result_T_39,_decode_result_T_41,_decode_result_T_43,
    _decode_result_T_76,_decode_result_T_124,_decode_result_T_142}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_1 = |_decode_result_orMatrixOutputs_T; // @[pla.scala 114:39]
  wire [2:0] _decode_result_orMatrixOutputs_T_2 = {_decode_result_T_35,_decode_result_T_45,_decode_result_T_55}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_3 = |_decode_result_orMatrixOutputs_T_2; // @[pla.scala 114:39]
  wire [2:0] _decode_result_orMatrixOutputs_T_4 = {_decode_result_T_35,_decode_result_T_51,_decode_result_T_114}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_5 = |_decode_result_orMatrixOutputs_T_4; // @[pla.scala 114:39]
  wire [1:0] _decode_result_orMatrixOutputs_T_6 = {_decode_result_T_53,_decode_result_T_55}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_7 = |_decode_result_orMatrixOutputs_T_6; // @[pla.scala 114:39]
  wire [9:0] decode_result_orMatrixOutputs_lo_1 = {_decode_result_T_84,_decode_result_T_90,_decode_result_T_94,
    _decode_result_T_98,_decode_result_T_102,_decode_result_T_112,_decode_result_T_122,_decode_result_T_136,
    _decode_result_T_140,_decode_result_T_150}; // @[Cat.scala 33:92]
  wire [9:0] decode_result_orMatrixOutputs_hi_3 = {_decode_result_T_7,_decode_result_T_11,_decode_result_T_15,
    _decode_result_T_29,_decode_result_T_31,_decode_result_T_33,_decode_result_T_37,_decode_result_T_63,
    _decode_result_T_65,_decode_result_T_74}; // @[Cat.scala 33:92]
  wire [19:0] _decode_result_orMatrixOutputs_T_8 = {decode_result_orMatrixOutputs_hi_3,
    decode_result_orMatrixOutputs_lo_1}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_9 = |_decode_result_orMatrixOutputs_T_8; // @[pla.scala 114:39]
  wire [4:0] _decode_result_orMatrixOutputs_T_10 = {_decode_result_T_1,_decode_result_T_19,_decode_result_T_35,
    _decode_result_T_45,_decode_result_T_53}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_11 = |_decode_result_orMatrixOutputs_T_10; // @[pla.scala 114:39]
  wire [6:0] _decode_result_orMatrixOutputs_T_12 = {_decode_result_T_5,_decode_result_T_19,_decode_result_T_25,
    _decode_result_T_35,_decode_result_T_51,_decode_result_T_53,_decode_result_T_114}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_13 = |_decode_result_orMatrixOutputs_T_12; // @[pla.scala 114:39]
  wire [2:0] _decode_result_orMatrixOutputs_T_14 = {_decode_result_T_21,_decode_result_T_53,_decode_result_T_116}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_15 = |_decode_result_orMatrixOutputs_T_14; // @[pla.scala 114:39]
  wire [9:0] _decode_result_orMatrixOutputs_T_16 = {_decode_result_T_5,_decode_result_T_19,_decode_result_T_25,
    _decode_result_T_47,_decode_result_T_51,_decode_result_T_72,_decode_result_T_86,_decode_result_T_114,
    _decode_result_T_144,_decode_result_T_152}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_17 = |_decode_result_orMatrixOutputs_T_16; // @[pla.scala 114:39]
  wire [1:0] _decode_result_orMatrixOutputs_T_18 = {_decode_result_T_70,_decode_result_T_166}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_19 = |_decode_result_orMatrixOutputs_T_18; // @[pla.scala 114:39]
  wire [1:0] _decode_result_orMatrixOutputs_T_20 = {_decode_result_T_132,_decode_result_T_138}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_21 = |_decode_result_orMatrixOutputs_T_20; // @[pla.scala 114:39]
  wire [1:0] _decode_result_orMatrixOutputs_T_22 = {_decode_result_T_23,_decode_result_T_138}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_23 = |_decode_result_orMatrixOutputs_T_22; // @[pla.scala 114:39]
  wire  _decode_result_orMatrixOutputs_T_24 = |_decode_result_T_80; // @[pla.scala 114:39]
  wire  _decode_result_orMatrixOutputs_T_25 = |_decode_result_T_100; // @[pla.scala 114:39]
  wire  _decode_result_orMatrixOutputs_T_26 = |_decode_result_T_68; // @[pla.scala 114:39]
  wire [3:0] _decode_result_orMatrixOutputs_T_27 = {_decode_result_T_47,_decode_result_T_86,_decode_result_T_144,
    _decode_result_T_152}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_28 = |_decode_result_orMatrixOutputs_T_27; // @[pla.scala 114:39]
  wire [3:0] _decode_result_orMatrixOutputs_T_29 = {_decode_result_T_45,_decode_result_T_144,_decode_result_T_172,
    _decode_result_T_176}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_30 = |_decode_result_orMatrixOutputs_T_29; // @[pla.scala 114:39]
  wire [4:0] _decode_result_orMatrixOutputs_T_31 = {_decode_result_T_3,_decode_result_T_146,_decode_result_T_152,
    _decode_result_T_174,_decode_result_T_178}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_32 = |_decode_result_orMatrixOutputs_T_31; // @[pla.scala 114:39]
  wire [1:0] _decode_result_orMatrixOutputs_T_33 = {_decode_result_T_49,_decode_result_T_106}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_34 = |_decode_result_orMatrixOutputs_T_33; // @[pla.scala 114:39]
  wire [3:0] _decode_result_orMatrixOutputs_T_35 = {_decode_result_T_144,_decode_result_T_152,_decode_result_T_164,
    _decode_result_T_172}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_36 = |_decode_result_orMatrixOutputs_T_35; // @[pla.scala 114:39]
  wire  _decode_result_orMatrixOutputs_T_37 = |_decode_result_T_47; // @[pla.scala 114:39]
  wire [1:0] _decode_result_orMatrixOutputs_T_38 = {_decode_result_T_72,_decode_result_T_104}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_39 = |_decode_result_orMatrixOutputs_T_38; // @[pla.scala 114:39]
  wire  _decode_result_orMatrixOutputs_T_40 = |_decode_result_T_86; // @[pla.scala 114:39]
  wire  _decode_result_orMatrixOutputs_T_41 = |_decode_result_T_110; // @[pla.scala 114:39]
  wire [2:0] _decode_result_orMatrixOutputs_T_42 = {_decode_result_T_19,_decode_result_T_51,_decode_result_T_114}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_43 = |_decode_result_orMatrixOutputs_T_42; // @[pla.scala 114:39]
  wire [1:0] _decode_result_orMatrixOutputs_T_44 = {_decode_result_T_19,_decode_result_T_53}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_45 = |_decode_result_orMatrixOutputs_T_44; // @[pla.scala 114:39]
  wire [2:0] _decode_result_orMatrixOutputs_T_46 = {_decode_result_T_72,_decode_result_T_78,_decode_result_T_120}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_47 = |_decode_result_orMatrixOutputs_T_46; // @[pla.scala 114:39]
  wire [5:0] _decode_result_orMatrixOutputs_T_48 = {_decode_result_T_51,_decode_result_T_104,_decode_result_T_126,
    _decode_result_T_128,_decode_result_T_168,_decode_result_T_170}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_49 = |_decode_result_orMatrixOutputs_T_48; // @[pla.scala 114:39]
  wire [4:0] _decode_result_orMatrixOutputs_T_50 = {_decode_result_T_88,_decode_result_T_108,_decode_result_T_110,
    _decode_result_T_114,_decode_result_T_126}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_51 = |_decode_result_orMatrixOutputs_T_50; // @[pla.scala 114:39]
  wire [3:0] _decode_result_orMatrixOutputs_T_52 = {_decode_result_T_88,_decode_result_T_114,_decode_result_T_168,
    _decode_result_T_170}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_53 = |_decode_result_orMatrixOutputs_T_52; // @[pla.scala 114:39]
  wire [6:0] decode_result_orMatrixOutputs_lo_12 = {_decode_result_T_67,_decode_result_T_94,_decode_result_T_98,
    _decode_result_T_118,_decode_result_T_150,_decode_result_T_156,_decode_result_T_162}; // @[Cat.scala 33:92]
  wire [13:0] _decode_result_orMatrixOutputs_T_54 = {_decode_result_T_9,_decode_result_T_11,_decode_result_T_13,
    _decode_result_T_27,_decode_result_T_57,_decode_result_T_63,_decode_result_T_65,decode_result_orMatrixOutputs_lo_12}
    ; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_55 = |_decode_result_orMatrixOutputs_T_54; // @[pla.scala 114:39]
  wire [8:0] _decode_result_orMatrixOutputs_T_56 = {_decode_result_T_9,_decode_result_T_11,_decode_result_T_13,
    _decode_result_T_94,_decode_result_T_98,_decode_result_T_134,_decode_result_T_136,_decode_result_T_140,
    _decode_result_T_150}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_57 = |_decode_result_orMatrixOutputs_T_56; // @[pla.scala 114:39]
  wire [5:0] _decode_result_orMatrixOutputs_T_58 = {_decode_result_T_27,_decode_result_T_67,_decode_result_T_84,
    _decode_result_T_102,_decode_result_T_156,_decode_result_T_162}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_59 = |_decode_result_orMatrixOutputs_T_58; // @[pla.scala 114:39]
  wire  _decode_result_orMatrixOutputs_T_60 = |_decode_result_T_67; // @[pla.scala 114:39]
  wire  _decode_result_orMatrixOutputs_T_61 = |_decode_result_T_130; // @[pla.scala 114:39]
  wire [5:0] decode_result_orMatrixOutputs_lo_lo_4 = {_decode_result_T_122,_decode_result_T_142,_decode_result_T_148,
    _decode_result_T_154,_decode_result_T_158,_decode_result_T_160}; // @[Cat.scala 33:92]
  wire [12:0] decode_result_orMatrixOutputs_lo_15 = {_decode_result_T_82,_decode_result_T_90,_decode_result_T_92,
    _decode_result_T_96,_decode_result_T_102,_decode_result_T_112,_decode_result_T_118,
    decode_result_orMatrixOutputs_lo_lo_4}; // @[Cat.scala 33:92]
  wire [6:0] decode_result_orMatrixOutputs_hi_lo_5 = {_decode_result_T_39,_decode_result_T_41,_decode_result_T_43,
    _decode_result_T_59,_decode_result_T_61,_decode_result_T_65,_decode_result_T_76}; // @[Cat.scala 33:92]
  wire [26:0] _decode_result_orMatrixOutputs_T_62 = {_decode_result_T_7,_decode_result_T_11,_decode_result_T_13,
    _decode_result_T_17,_decode_result_T_27,_decode_result_T_33,_decode_result_T_37,
    decode_result_orMatrixOutputs_hi_lo_5,decode_result_orMatrixOutputs_lo_15}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_63 = |_decode_result_orMatrixOutputs_T_62; // @[pla.scala 114:39]
  wire [6:0] decode_result_orMatrixOutputs_lo_lo_5 = {_decode_result_T_122,_decode_result_T_136,_decode_result_T_140,
    _decode_result_T_150,_decode_result_T_156,_decode_result_T_158,_decode_result_T_162}; // @[Cat.scala 33:92]
  wire [13:0] decode_result_orMatrixOutputs_lo_16 = {_decode_result_T_84,_decode_result_T_90,_decode_result_T_94,
    _decode_result_T_98,_decode_result_T_102,_decode_result_T_112,_decode_result_T_118,
    decode_result_orMatrixOutputs_lo_lo_5}; // @[Cat.scala 33:92]
  wire [6:0] decode_result_orMatrixOutputs_hi_lo_6 = {_decode_result_T_37,_decode_result_T_57,_decode_result_T_61,
    _decode_result_T_63,_decode_result_T_65,_decode_result_T_67,_decode_result_T_74}; // @[Cat.scala 33:92]
  wire [27:0] _decode_result_orMatrixOutputs_T_64 = {_decode_result_T_7,_decode_result_T_11,_decode_result_T_13,
    _decode_result_T_27,_decode_result_T_29,_decode_result_T_31,_decode_result_T_33,
    decode_result_orMatrixOutputs_hi_lo_6,decode_result_orMatrixOutputs_lo_16}; // @[Cat.scala 33:92]
  wire  _decode_result_orMatrixOutputs_T_65 = |_decode_result_orMatrixOutputs_T_64; // @[pla.scala 114:39]
  wire [9:0] decode_result_orMatrixOutputs_lo_hi_10 = {_decode_result_orMatrixOutputs_T_34,
    _decode_result_orMatrixOutputs_T_32,_decode_result_orMatrixOutputs_T_30,_decode_result_orMatrixOutputs_T_28,
    _decode_result_orMatrixOutputs_T_26,_decode_result_orMatrixOutputs_T_25,_decode_result_orMatrixOutputs_T_24,
    _decode_result_orMatrixOutputs_T_23,_decode_result_orMatrixOutputs_T_21,_decode_result_orMatrixOutputs_T_19}; // @[Cat.scala 33:92]
  wire [18:0] decode_result_orMatrixOutputs_lo_17 = {decode_result_orMatrixOutputs_lo_hi_10,
    _decode_result_orMatrixOutputs_T_17,_decode_result_orMatrixOutputs_T_15,_decode_result_orMatrixOutputs_T_13,
    _decode_result_orMatrixOutputs_T_11,_decode_result_orMatrixOutputs_T_9,_decode_result_orMatrixOutputs_T_7,
    _decode_result_orMatrixOutputs_T_5,_decode_result_orMatrixOutputs_T_3,_decode_result_orMatrixOutputs_T_1}; // @[Cat.scala 33:92]
  wire [9:0] decode_result_orMatrixOutputs_hi_hi_13 = {_decode_result_orMatrixOutputs_T_65,
    _decode_result_orMatrixOutputs_T_63,_decode_result_orMatrixOutputs_T_61,_decode_result_orMatrixOutputs_T_60,
    _decode_result_orMatrixOutputs_T_59,_decode_result_orMatrixOutputs_T_57,_decode_result_orMatrixOutputs_T_55,
    _decode_result_orMatrixOutputs_T_53,_decode_result_orMatrixOutputs_T_51,_decode_result_orMatrixOutputs_T_49}; // @[Cat.scala 33:92]
  wire [18:0] decode_result_orMatrixOutputs_hi_22 = {decode_result_orMatrixOutputs_hi_hi_13,
    _decode_result_orMatrixOutputs_T_47,_decode_result_orMatrixOutputs_T_45,_decode_result_orMatrixOutputs_T_43,1'h0,
    _decode_result_orMatrixOutputs_T_41,_decode_result_orMatrixOutputs_T_40,_decode_result_orMatrixOutputs_T_39,
    _decode_result_orMatrixOutputs_T_37,_decode_result_orMatrixOutputs_T_36}; // @[Cat.scala 33:92]
  wire [37:0] decode_result_orMatrixOutputs = {decode_result_orMatrixOutputs_hi_22,decode_result_orMatrixOutputs_lo_17}; // @[Cat.scala 33:92]
  wire  _decode_result_invMatrixOutputs_T_1 = ~decode_result_orMatrixOutputs[0]; // @[pla.scala 123:40]
  wire  _decode_result_invMatrixOutputs_T_38 = ~decode_result_orMatrixOutputs[36]; // @[pla.scala 123:40]
  wire [9:0] decode_result_invMatrixOutputs_lo_hi = {decode_result_orMatrixOutputs[18],decode_result_orMatrixOutputs[17]
    ,decode_result_orMatrixOutputs[16],decode_result_orMatrixOutputs[15],decode_result_orMatrixOutputs[14],
    decode_result_orMatrixOutputs[13],decode_result_orMatrixOutputs[12],decode_result_orMatrixOutputs[11],
    decode_result_orMatrixOutputs[10],decode_result_orMatrixOutputs[9]}; // @[Cat.scala 33:92]
  wire [18:0] decode_result_invMatrixOutputs_lo = {decode_result_invMatrixOutputs_lo_hi,decode_result_orMatrixOutputs[8]
    ,decode_result_orMatrixOutputs[7],decode_result_orMatrixOutputs[6],decode_result_orMatrixOutputs[5],
    decode_result_orMatrixOutputs[4],decode_result_orMatrixOutputs[3],decode_result_orMatrixOutputs[2],
    decode_result_orMatrixOutputs[1],_decode_result_invMatrixOutputs_T_1}; // @[Cat.scala 33:92]
  wire [9:0] decode_result_invMatrixOutputs_hi_hi = {decode_result_orMatrixOutputs[37],
    _decode_result_invMatrixOutputs_T_38,decode_result_orMatrixOutputs[35],decode_result_orMatrixOutputs[34],
    decode_result_orMatrixOutputs[33],decode_result_orMatrixOutputs[32],decode_result_orMatrixOutputs[31],
    decode_result_orMatrixOutputs[30],decode_result_orMatrixOutputs[29],decode_result_orMatrixOutputs[28]}; // @[Cat.scala 33:92]
  wire [18:0] decode_result_invMatrixOutputs_hi = {decode_result_invMatrixOutputs_hi_hi,decode_result_orMatrixOutputs[27
    ],decode_result_orMatrixOutputs[26],decode_result_orMatrixOutputs[25],decode_result_orMatrixOutputs[24],
    decode_result_orMatrixOutputs[23],decode_result_orMatrixOutputs[22],decode_result_orMatrixOutputs[21],
    decode_result_orMatrixOutputs[20],decode_result_orMatrixOutputs[19]}; // @[Cat.scala 33:92]
  wire [37:0] decode_result_invMatrixOutputs = {decode_result_invMatrixOutputs_hi,decode_result_invMatrixOutputs_lo}; // @[Cat.scala 33:92]
  wire  uop_dw = decode_result_invMatrixOutputs[0]; // @[MicroOp.scala 56:20]
  wire [2:0] imm_type = decode_result_invMatrixOutputs[3:1]; // @[MicroOp.scala 58:20]
  wire  uop_rd_wen = decode_result_invMatrixOutputs[4]; // @[MicroOp.scala 56:20]
  wire [1:0] uop_rs2_src = decode_result_invMatrixOutputs[6:5]; // @[MicroOp.scala 58:20]
  wire [1:0] uop_rs1_src = decode_result_invMatrixOutputs[8:7]; // @[MicroOp.scala 58:20]
  wire [2:0] uop_sys_op = decode_result_invMatrixOutputs[11:9]; // @[MicroOp.scala 58:20]
  wire [1:0] uop_csr_op = decode_result_invMatrixOutputs[13:12]; // @[MicroOp.scala 58:20]
  wire [1:0] uop_mem_len = decode_result_invMatrixOutputs[15:14]; // @[MicroOp.scala 58:20]
  wire [4:0] uop_lsu_op = decode_result_invMatrixOutputs[20:16]; // @[MicroOp.scala 58:20]
  wire [3:0] uop_mdu_op = decode_result_invMatrixOutputs[24:21]; // @[MicroOp.scala 58:20]
  wire [1:0] uop_jmp_op = decode_result_invMatrixOutputs[26:25]; // @[MicroOp.scala 58:20]
  wire [3:0] uop_alu_op = decode_result_invMatrixOutputs[30:27]; // @[MicroOp.scala 58:20]
  wire [2:0] uop_fu = decode_result_invMatrixOutputs[33:31]; // @[MicroOp.scala 58:20]
  wire [20:0] _imm_i_T_2 = decode_result_andMatrixInput_4_58 ? 21'h1fffff : 21'h0; // @[Bitwise.scala 77:12]
  wire [31:0] imm_i = {_imm_i_T_2,io_in_instr[30:20]}; // @[Cat.scala 33:92]
  wire [31:0] imm_s = {_imm_i_T_2,io_in_instr[30:25],uop_rd_index}; // @[Cat.scala 33:92]
  wire [19:0] _imm_b_T_2 = decode_result_andMatrixInput_4_58 ? 20'hfffff : 20'h0; // @[Bitwise.scala 77:12]
  wire [31:0] imm_b = {_imm_b_T_2,io_in_instr[7],io_in_instr[30:25],io_in_instr[11:8],1'h0}; // @[Cat.scala 33:92]
  wire [31:0] imm_u = {io_in_instr[31:12],12'h0}; // @[Cat.scala 33:92]
  wire [11:0] _imm_j_T_2 = decode_result_andMatrixInput_4_58 ? 12'hfff : 12'h0; // @[Bitwise.scala 77:12]
  wire [31:0] imm_j = {_imm_j_T_2,io_in_instr[19:12],decode_result_andMatrixInput_20_2,io_in_instr[30:21],1'h0}; // @[Cat.scala 33:92]
  wire [31:0] imm_csr = {27'h0,uop_rs1_index}; // @[Cat.scala 33:92]
  wire [31:0] _uop_imm_T_1 = 3'h0 == imm_type ? imm_i : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] _uop_imm_T_3 = 3'h1 == imm_type ? imm_s : _uop_imm_T_1; // @[Mux.scala 81:58]
  wire [31:0] _uop_imm_T_5 = 3'h2 == imm_type ? imm_b : _uop_imm_T_3; // @[Mux.scala 81:58]
  wire [31:0] _uop_imm_T_7 = 3'h3 == imm_type ? imm_u : _uop_imm_T_5; // @[Mux.scala 81:58]
  wire [31:0] _uop_imm_T_9 = 3'h4 == imm_type ? imm_j : _uop_imm_T_7; // @[Mux.scala 81:58]
  wire [31:0] uop_imm = 3'h5 == imm_type ? imm_csr : _uop_imm_T_9; // @[Mux.scala 81:58]
  wire [2:0] _GEN_0 = io_in_access_fault ? 3'h2 : decode_result_invMatrixOutputs[36:34]; // @[Decode.scala 30:36 31:17 MicroOp.scala 58:15]
  wire  _GEN_1 = io_in_access_fault ? 1'h0 : decode_result_invMatrixOutputs[37]; // @[Decode.scala 30:36 32:17 MicroOp.scala 56:15]
  wire [2:0] _GEN_2 = io_in_page_fault ? 3'h3 : _GEN_0; // @[Decode.scala 27:28 28:17]
  wire  _GEN_3 = io_in_page_fault ? 1'h0 : _GEN_1; // @[Decode.scala 27:28 29:17]
  wire [2:0] uop_exc = io_in_valid ? _GEN_2 : decode_result_invMatrixOutputs[36:34]; // @[Decode.scala 26:21 MicroOp.scala 58:15]
  wire  uop_valid = io_in_valid ? _GEN_3 : decode_result_invMatrixOutputs[37]; // @[Decode.scala 26:21 MicroOp.scala 56:15]
  assign io_out_valid = io_in_valid & uop_valid; // @[Decode.scala 36:16]
  assign io_out_exc = io_in_valid ? uop_exc : 3'h0; // @[Decode.scala 36:16]
  assign io_out_pc = io_in_valid ? io_in_pc : 64'h0; // @[Decode.scala 36:16]
  assign io_out_npc = io_in_valid ? uop_npc : 64'h0; // @[Decode.scala 36:16]
  assign io_out_instr = io_in_valid ? io_in_instr : 32'h0; // @[Decode.scala 36:16]
  assign io_out_fu = io_in_valid ? uop_fu : 3'h0; // @[Decode.scala 36:16]
  assign io_out_alu_op = io_in_valid ? uop_alu_op : 4'h0; // @[Decode.scala 36:16]
  assign io_out_jmp_op = io_in_valid ? uop_jmp_op : 2'h0; // @[Decode.scala 36:16]
  assign io_out_mdu_op = io_in_valid ? uop_mdu_op : 4'h0; // @[Decode.scala 36:16]
  assign io_out_lsu_op = io_in_valid ? uop_lsu_op : 5'h0; // @[Decode.scala 36:16]
  assign io_out_mem_len = io_in_valid ? uop_mem_len : 2'h0; // @[Decode.scala 36:16]
  assign io_out_csr_op = io_in_valid ? uop_csr_op : 2'h0; // @[Decode.scala 36:16]
  assign io_out_sys_op = io_in_valid ? uop_sys_op : 3'h0; // @[Decode.scala 36:16]
  assign io_out_rs1_src = io_in_valid ? uop_rs1_src : 2'h0; // @[Decode.scala 36:16]
  assign io_out_rs2_src = io_in_valid ? uop_rs2_src : 2'h0; // @[Decode.scala 36:16]
  assign io_out_rs1_index = io_in_valid ? uop_rs1_index : 5'h0; // @[Decode.scala 36:16]
  assign io_out_rs2_index = io_in_valid ? uop_rs2_index : 5'h0; // @[Decode.scala 36:16]
  assign io_out_rd_index = io_in_valid ? uop_rd_index : 5'h0; // @[Decode.scala 36:16]
  assign io_out_rd_wen = io_in_valid & uop_rd_wen; // @[Decode.scala 36:16]
  assign io_out_imm = io_in_valid ? uop_imm : 32'h0; // @[Decode.scala 36:16]
  assign io_out_dw = io_in_valid & uop_dw; // @[Decode.scala 36:16]
endmodule
module RegFile(
  input         clock,
  input         reset,
  input  [4:0]  io_rs1_index,
  input  [4:0]  io_rs2_index,
  output [63:0] io_rs1_data,
  output [63:0] io_rs2_data,
  input  [4:0]  io_rd_index,
  input  [63:0] io_rd_data,
  input         io_rd_wen
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] rf_0; // @[RegFile.scala 21:19]
  reg [63:0] rf_1; // @[RegFile.scala 21:19]
  reg [63:0] rf_2; // @[RegFile.scala 21:19]
  reg [63:0] rf_3; // @[RegFile.scala 21:19]
  reg [63:0] rf_4; // @[RegFile.scala 21:19]
  reg [63:0] rf_5; // @[RegFile.scala 21:19]
  reg [63:0] rf_6; // @[RegFile.scala 21:19]
  reg [63:0] rf_7; // @[RegFile.scala 21:19]
  reg [63:0] rf_8; // @[RegFile.scala 21:19]
  reg [63:0] rf_9; // @[RegFile.scala 21:19]
  reg [63:0] rf_10; // @[RegFile.scala 21:19]
  reg [63:0] rf_11; // @[RegFile.scala 21:19]
  reg [63:0] rf_12; // @[RegFile.scala 21:19]
  reg [63:0] rf_13; // @[RegFile.scala 21:19]
  reg [63:0] rf_14; // @[RegFile.scala 21:19]
  reg [63:0] rf_15; // @[RegFile.scala 21:19]
  reg [63:0] rf_16; // @[RegFile.scala 21:19]
  reg [63:0] rf_17; // @[RegFile.scala 21:19]
  reg [63:0] rf_18; // @[RegFile.scala 21:19]
  reg [63:0] rf_19; // @[RegFile.scala 21:19]
  reg [63:0] rf_20; // @[RegFile.scala 21:19]
  reg [63:0] rf_21; // @[RegFile.scala 21:19]
  reg [63:0] rf_22; // @[RegFile.scala 21:19]
  reg [63:0] rf_23; // @[RegFile.scala 21:19]
  reg [63:0] rf_24; // @[RegFile.scala 21:19]
  reg [63:0] rf_25; // @[RegFile.scala 21:19]
  reg [63:0] rf_26; // @[RegFile.scala 21:19]
  reg [63:0] rf_27; // @[RegFile.scala 21:19]
  reg [63:0] rf_28; // @[RegFile.scala 21:19]
  reg [63:0] rf_29; // @[RegFile.scala 21:19]
  reg [63:0] rf_30; // @[RegFile.scala 21:19]
  wire  _T_1 = io_rd_wen & io_rd_index != 5'h0; // @[RegFile.scala 23:18]
  wire [4:0] _T_2 = ~io_rd_index; // @[RegFile.scala 18:28]
  wire [4:0] _io_rs1_data_T_1 = ~io_rs1_index; // @[RegFile.scala 18:28]
  wire [63:0] _GEN_63 = 5'h1 == _io_rs1_data_T_1 ? rf_1 : rf_0; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_64 = 5'h2 == _io_rs1_data_T_1 ? rf_2 : _GEN_63; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_65 = 5'h3 == _io_rs1_data_T_1 ? rf_3 : _GEN_64; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_66 = 5'h4 == _io_rs1_data_T_1 ? rf_4 : _GEN_65; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_67 = 5'h5 == _io_rs1_data_T_1 ? rf_5 : _GEN_66; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_68 = 5'h6 == _io_rs1_data_T_1 ? rf_6 : _GEN_67; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_69 = 5'h7 == _io_rs1_data_T_1 ? rf_7 : _GEN_68; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_70 = 5'h8 == _io_rs1_data_T_1 ? rf_8 : _GEN_69; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_71 = 5'h9 == _io_rs1_data_T_1 ? rf_9 : _GEN_70; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_72 = 5'ha == _io_rs1_data_T_1 ? rf_10 : _GEN_71; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_73 = 5'hb == _io_rs1_data_T_1 ? rf_11 : _GEN_72; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_74 = 5'hc == _io_rs1_data_T_1 ? rf_12 : _GEN_73; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_75 = 5'hd == _io_rs1_data_T_1 ? rf_13 : _GEN_74; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_76 = 5'he == _io_rs1_data_T_1 ? rf_14 : _GEN_75; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_77 = 5'hf == _io_rs1_data_T_1 ? rf_15 : _GEN_76; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_78 = 5'h10 == _io_rs1_data_T_1 ? rf_16 : _GEN_77; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_79 = 5'h11 == _io_rs1_data_T_1 ? rf_17 : _GEN_78; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_80 = 5'h12 == _io_rs1_data_T_1 ? rf_18 : _GEN_79; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_81 = 5'h13 == _io_rs1_data_T_1 ? rf_19 : _GEN_80; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_82 = 5'h14 == _io_rs1_data_T_1 ? rf_20 : _GEN_81; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_83 = 5'h15 == _io_rs1_data_T_1 ? rf_21 : _GEN_82; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_84 = 5'h16 == _io_rs1_data_T_1 ? rf_22 : _GEN_83; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_85 = 5'h17 == _io_rs1_data_T_1 ? rf_23 : _GEN_84; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_86 = 5'h18 == _io_rs1_data_T_1 ? rf_24 : _GEN_85; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_87 = 5'h19 == _io_rs1_data_T_1 ? rf_25 : _GEN_86; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_88 = 5'h1a == _io_rs1_data_T_1 ? rf_26 : _GEN_87; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_89 = 5'h1b == _io_rs1_data_T_1 ? rf_27 : _GEN_88; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_90 = 5'h1c == _io_rs1_data_T_1 ? rf_28 : _GEN_89; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_91 = 5'h1d == _io_rs1_data_T_1 ? rf_29 : _GEN_90; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _GEN_92 = 5'h1e == _io_rs1_data_T_1 ? rf_30 : _GEN_91; // @[RegFile.scala 27:{21,21}]
  wire [63:0] _io_rs1_data_T_2 = io_rs1_index != 5'h0 ? _GEN_92 : 64'h0; // @[RegFile.scala 27:21]
  wire [4:0] _io_rs2_data_T_1 = ~io_rs2_index; // @[RegFile.scala 18:28]
  wire [63:0] _GEN_94 = 5'h1 == _io_rs2_data_T_1 ? rf_1 : rf_0; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_95 = 5'h2 == _io_rs2_data_T_1 ? rf_2 : _GEN_94; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_96 = 5'h3 == _io_rs2_data_T_1 ? rf_3 : _GEN_95; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_97 = 5'h4 == _io_rs2_data_T_1 ? rf_4 : _GEN_96; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_98 = 5'h5 == _io_rs2_data_T_1 ? rf_5 : _GEN_97; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_99 = 5'h6 == _io_rs2_data_T_1 ? rf_6 : _GEN_98; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_100 = 5'h7 == _io_rs2_data_T_1 ? rf_7 : _GEN_99; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_101 = 5'h8 == _io_rs2_data_T_1 ? rf_8 : _GEN_100; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_102 = 5'h9 == _io_rs2_data_T_1 ? rf_9 : _GEN_101; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_103 = 5'ha == _io_rs2_data_T_1 ? rf_10 : _GEN_102; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_104 = 5'hb == _io_rs2_data_T_1 ? rf_11 : _GEN_103; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_105 = 5'hc == _io_rs2_data_T_1 ? rf_12 : _GEN_104; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_106 = 5'hd == _io_rs2_data_T_1 ? rf_13 : _GEN_105; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_107 = 5'he == _io_rs2_data_T_1 ? rf_14 : _GEN_106; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_108 = 5'hf == _io_rs2_data_T_1 ? rf_15 : _GEN_107; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_109 = 5'h10 == _io_rs2_data_T_1 ? rf_16 : _GEN_108; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_110 = 5'h11 == _io_rs2_data_T_1 ? rf_17 : _GEN_109; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_111 = 5'h12 == _io_rs2_data_T_1 ? rf_18 : _GEN_110; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_112 = 5'h13 == _io_rs2_data_T_1 ? rf_19 : _GEN_111; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_113 = 5'h14 == _io_rs2_data_T_1 ? rf_20 : _GEN_112; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_114 = 5'h15 == _io_rs2_data_T_1 ? rf_21 : _GEN_113; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_115 = 5'h16 == _io_rs2_data_T_1 ? rf_22 : _GEN_114; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_116 = 5'h17 == _io_rs2_data_T_1 ? rf_23 : _GEN_115; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_117 = 5'h18 == _io_rs2_data_T_1 ? rf_24 : _GEN_116; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_118 = 5'h19 == _io_rs2_data_T_1 ? rf_25 : _GEN_117; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_119 = 5'h1a == _io_rs2_data_T_1 ? rf_26 : _GEN_118; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_120 = 5'h1b == _io_rs2_data_T_1 ? rf_27 : _GEN_119; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_121 = 5'h1c == _io_rs2_data_T_1 ? rf_28 : _GEN_120; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_122 = 5'h1d == _io_rs2_data_T_1 ? rf_29 : _GEN_121; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _GEN_123 = 5'h1e == _io_rs2_data_T_1 ? rf_30 : _GEN_122; // @[RegFile.scala 28:{21,21}]
  wire [63:0] _io_rs2_data_T_2 = io_rs2_index != 5'h0 ? _GEN_123 : 64'h0; // @[RegFile.scala 28:21]
  wire [63:0] _GEN_124 = io_rd_index == io_rs1_index ? io_rd_data : _io_rs1_data_T_2; // @[RegFile.scala 27:15 32:40 33:19]
  wire [63:0] _GEN_125 = io_rd_index == io_rs2_index ? io_rd_data : _io_rs2_data_T_2; // @[RegFile.scala 28:15 35:40 36:19]
  assign io_rs1_data = _T_1 ? _GEN_124 : _io_rs1_data_T_2; // @[RegFile.scala 27:15 31:44]
  assign io_rs2_data = _T_1 ? _GEN_125 : _io_rs2_data_T_2; // @[RegFile.scala 28:15 31:44]
  always @(posedge clock) begin
    if (reset) begin // @[RegFile.scala 21:19]
      rf_0 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h0 == _T_2) begin // @[RegFile.scala 24:25]
        rf_0 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_1 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h1 == _T_2) begin // @[RegFile.scala 24:25]
        rf_1 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_2 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h2 == _T_2) begin // @[RegFile.scala 24:25]
        rf_2 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_3 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h3 == _T_2) begin // @[RegFile.scala 24:25]
        rf_3 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_4 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h4 == _T_2) begin // @[RegFile.scala 24:25]
        rf_4 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_5 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h5 == _T_2) begin // @[RegFile.scala 24:25]
        rf_5 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_6 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h6 == _T_2) begin // @[RegFile.scala 24:25]
        rf_6 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_7 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h7 == _T_2) begin // @[RegFile.scala 24:25]
        rf_7 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_8 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h8 == _T_2) begin // @[RegFile.scala 24:25]
        rf_8 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_9 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h9 == _T_2) begin // @[RegFile.scala 24:25]
        rf_9 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_10 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'ha == _T_2) begin // @[RegFile.scala 24:25]
        rf_10 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_11 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'hb == _T_2) begin // @[RegFile.scala 24:25]
        rf_11 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_12 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'hc == _T_2) begin // @[RegFile.scala 24:25]
        rf_12 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_13 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'hd == _T_2) begin // @[RegFile.scala 24:25]
        rf_13 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_14 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'he == _T_2) begin // @[RegFile.scala 24:25]
        rf_14 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_15 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'hf == _T_2) begin // @[RegFile.scala 24:25]
        rf_15 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_16 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h10 == _T_2) begin // @[RegFile.scala 24:25]
        rf_16 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_17 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h11 == _T_2) begin // @[RegFile.scala 24:25]
        rf_17 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_18 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h12 == _T_2) begin // @[RegFile.scala 24:25]
        rf_18 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_19 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h13 == _T_2) begin // @[RegFile.scala 24:25]
        rf_19 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_20 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h14 == _T_2) begin // @[RegFile.scala 24:25]
        rf_20 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_21 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h15 == _T_2) begin // @[RegFile.scala 24:25]
        rf_21 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_22 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h16 == _T_2) begin // @[RegFile.scala 24:25]
        rf_22 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_23 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h17 == _T_2) begin // @[RegFile.scala 24:25]
        rf_23 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_24 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h18 == _T_2) begin // @[RegFile.scala 24:25]
        rf_24 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_25 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h19 == _T_2) begin // @[RegFile.scala 24:25]
        rf_25 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_26 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h1a == _T_2) begin // @[RegFile.scala 24:25]
        rf_26 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_27 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h1b == _T_2) begin // @[RegFile.scala 24:25]
        rf_27 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_28 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h1c == _T_2) begin // @[RegFile.scala 24:25]
        rf_28 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_29 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h1d == _T_2) begin // @[RegFile.scala 24:25]
        rf_29 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
    if (reset) begin // @[RegFile.scala 21:19]
      rf_30 <= 64'h0; // @[RegFile.scala 21:19]
    end else if (io_rd_wen & io_rd_index != 5'h0) begin // @[RegFile.scala 23:44]
      if (5'h1e == _T_2) begin // @[RegFile.scala 24:25]
        rf_30 <= io_rd_data; // @[RegFile.scala 24:25]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  rf_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  rf_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  rf_2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  rf_3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  rf_4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  rf_5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  rf_6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  rf_7 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  rf_8 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  rf_9 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  rf_10 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  rf_11 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  rf_12 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  rf_13 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  rf_14 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  rf_15 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  rf_16 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  rf_17 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  rf_18 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  rf_19 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  rf_20 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  rf_21 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  rf_22 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  rf_23 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  rf_24 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  rf_25 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  rf_26 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  rf_27 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  rf_28 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  rf_29 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  rf_30 = _RAND_30[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PipelineReg(
  input         clock,
  input         reset,
  input         io_in_uop_valid,
  input  [2:0]  io_in_uop_exc,
  input  [63:0] io_in_uop_pc,
  input  [63:0] io_in_uop_npc,
  input  [31:0] io_in_uop_instr,
  input  [2:0]  io_in_uop_fu,
  input  [3:0]  io_in_uop_alu_op,
  input  [1:0]  io_in_uop_jmp_op,
  input  [3:0]  io_in_uop_mdu_op,
  input  [4:0]  io_in_uop_lsu_op,
  input  [1:0]  io_in_uop_mem_len,
  input  [1:0]  io_in_uop_csr_op,
  input  [2:0]  io_in_uop_sys_op,
  input  [4:0]  io_in_uop_rd_index,
  input         io_in_uop_rd_wen,
  input  [31:0] io_in_uop_imm,
  input         io_in_uop_dw,
  input  [63:0] io_in_rs1_data,
  input  [63:0] io_in_rs2_data,
  input  [63:0] io_in_rs2_data_from_rf,
  input  [63:0] io_in_bp_npc,
  output        io_out_uop_valid,
  output [2:0]  io_out_uop_exc,
  output [63:0] io_out_uop_pc,
  output [63:0] io_out_uop_npc,
  output [31:0] io_out_uop_instr,
  output [2:0]  io_out_uop_fu,
  output [3:0]  io_out_uop_alu_op,
  output [1:0]  io_out_uop_jmp_op,
  output [3:0]  io_out_uop_mdu_op,
  output [4:0]  io_out_uop_lsu_op,
  output [1:0]  io_out_uop_mem_len,
  output [1:0]  io_out_uop_csr_op,
  output [2:0]  io_out_uop_sys_op,
  output [4:0]  io_out_uop_rd_index,
  output        io_out_uop_rd_wen,
  output [31:0] io_out_uop_imm,
  output        io_out_uop_dw,
  output [63:0] io_out_rs1_data,
  output [63:0] io_out_rs2_data,
  output [63:0] io_out_rs2_data_from_rf,
  output [63:0] io_out_bp_npc,
  input         io_en,
  input         io_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
`endif // RANDOMIZE_REG_INIT
  reg  reg_uop_valid; // @[Reg.scala 35:20]
  reg [2:0] reg_uop_exc; // @[Reg.scala 35:20]
  reg [63:0] reg_uop_pc; // @[Reg.scala 35:20]
  reg [63:0] reg_uop_npc; // @[Reg.scala 35:20]
  reg [31:0] reg_uop_instr; // @[Reg.scala 35:20]
  reg [2:0] reg_uop_fu; // @[Reg.scala 35:20]
  reg [3:0] reg_uop_alu_op; // @[Reg.scala 35:20]
  reg [1:0] reg_uop_jmp_op; // @[Reg.scala 35:20]
  reg [3:0] reg_uop_mdu_op; // @[Reg.scala 35:20]
  reg [4:0] reg_uop_lsu_op; // @[Reg.scala 35:20]
  reg [1:0] reg_uop_mem_len; // @[Reg.scala 35:20]
  reg [1:0] reg_uop_csr_op; // @[Reg.scala 35:20]
  reg [2:0] reg_uop_sys_op; // @[Reg.scala 35:20]
  reg [4:0] reg_uop_rd_index; // @[Reg.scala 35:20]
  reg  reg_uop_rd_wen; // @[Reg.scala 35:20]
  reg [31:0] reg_uop_imm; // @[Reg.scala 35:20]
  reg  reg_uop_dw; // @[Reg.scala 35:20]
  reg [63:0] reg_rs1_data; // @[Reg.scala 35:20]
  reg [63:0] reg_rs2_data; // @[Reg.scala 35:20]
  reg [63:0] reg_rs2_data_from_rf; // @[Reg.scala 35:20]
  reg [63:0] reg_bp_npc; // @[Reg.scala 35:20]
  assign io_out_uop_valid = reg_uop_valid; // @[DataType.scala 41:10]
  assign io_out_uop_exc = reg_uop_exc; // @[DataType.scala 41:10]
  assign io_out_uop_pc = reg_uop_pc; // @[DataType.scala 41:10]
  assign io_out_uop_npc = reg_uop_npc; // @[DataType.scala 41:10]
  assign io_out_uop_instr = reg_uop_instr; // @[DataType.scala 41:10]
  assign io_out_uop_fu = reg_uop_fu; // @[DataType.scala 41:10]
  assign io_out_uop_alu_op = reg_uop_alu_op; // @[DataType.scala 41:10]
  assign io_out_uop_jmp_op = reg_uop_jmp_op; // @[DataType.scala 41:10]
  assign io_out_uop_mdu_op = reg_uop_mdu_op; // @[DataType.scala 41:10]
  assign io_out_uop_lsu_op = reg_uop_lsu_op; // @[DataType.scala 41:10]
  assign io_out_uop_mem_len = reg_uop_mem_len; // @[DataType.scala 41:10]
  assign io_out_uop_csr_op = reg_uop_csr_op; // @[DataType.scala 41:10]
  assign io_out_uop_sys_op = reg_uop_sys_op; // @[DataType.scala 41:10]
  assign io_out_uop_rd_index = reg_uop_rd_index; // @[DataType.scala 41:10]
  assign io_out_uop_rd_wen = reg_uop_rd_wen; // @[DataType.scala 41:10]
  assign io_out_uop_imm = reg_uop_imm; // @[DataType.scala 41:10]
  assign io_out_uop_dw = reg_uop_dw; // @[DataType.scala 41:10]
  assign io_out_rs1_data = reg_rs1_data; // @[DataType.scala 41:10]
  assign io_out_rs2_data = reg_rs2_data; // @[DataType.scala 41:10]
  assign io_out_rs2_data_from_rf = reg_rs2_data_from_rf; // @[DataType.scala 41:10]
  assign io_out_bp_npc = reg_bp_npc; // @[DataType.scala 41:10]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 35:20]
      reg_uop_valid <= 1'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_flush) begin // @[DataType.scala 40:26]
        reg_uop_valid <= 1'h0;
      end else begin
        reg_uop_valid <= io_in_uop_valid;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      reg_uop_exc <= 3'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_flush) begin // @[DataType.scala 40:26]
        reg_uop_exc <= 3'h0;
      end else begin
        reg_uop_exc <= io_in_uop_exc;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      reg_uop_pc <= 64'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_flush) begin // @[DataType.scala 40:26]
        reg_uop_pc <= 64'h0;
      end else begin
        reg_uop_pc <= io_in_uop_pc;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      reg_uop_npc <= 64'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_flush) begin // @[DataType.scala 40:26]
        reg_uop_npc <= 64'h0;
      end else begin
        reg_uop_npc <= io_in_uop_npc;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      reg_uop_instr <= 32'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_flush) begin // @[DataType.scala 40:26]
        reg_uop_instr <= 32'h0;
      end else begin
        reg_uop_instr <= io_in_uop_instr;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      reg_uop_fu <= 3'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_flush) begin // @[DataType.scala 40:26]
        reg_uop_fu <= 3'h0;
      end else begin
        reg_uop_fu <= io_in_uop_fu;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      reg_uop_alu_op <= 4'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_flush) begin // @[DataType.scala 40:26]
        reg_uop_alu_op <= 4'h0;
      end else begin
        reg_uop_alu_op <= io_in_uop_alu_op;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      reg_uop_jmp_op <= 2'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_flush) begin // @[DataType.scala 40:26]
        reg_uop_jmp_op <= 2'h0;
      end else begin
        reg_uop_jmp_op <= io_in_uop_jmp_op;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      reg_uop_mdu_op <= 4'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_flush) begin // @[DataType.scala 40:26]
        reg_uop_mdu_op <= 4'h0;
      end else begin
        reg_uop_mdu_op <= io_in_uop_mdu_op;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      reg_uop_lsu_op <= 5'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_flush) begin // @[DataType.scala 40:26]
        reg_uop_lsu_op <= 5'h0;
      end else begin
        reg_uop_lsu_op <= io_in_uop_lsu_op;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      reg_uop_mem_len <= 2'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_flush) begin // @[DataType.scala 40:26]
        reg_uop_mem_len <= 2'h0;
      end else begin
        reg_uop_mem_len <= io_in_uop_mem_len;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      reg_uop_csr_op <= 2'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_flush) begin // @[DataType.scala 40:26]
        reg_uop_csr_op <= 2'h0;
      end else begin
        reg_uop_csr_op <= io_in_uop_csr_op;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      reg_uop_sys_op <= 3'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_flush) begin // @[DataType.scala 40:26]
        reg_uop_sys_op <= 3'h0;
      end else begin
        reg_uop_sys_op <= io_in_uop_sys_op;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      reg_uop_rd_index <= 5'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_flush) begin // @[DataType.scala 40:26]
        reg_uop_rd_index <= 5'h0;
      end else begin
        reg_uop_rd_index <= io_in_uop_rd_index;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      reg_uop_rd_wen <= 1'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_flush) begin // @[DataType.scala 40:26]
        reg_uop_rd_wen <= 1'h0;
      end else begin
        reg_uop_rd_wen <= io_in_uop_rd_wen;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      reg_uop_imm <= 32'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_flush) begin // @[DataType.scala 40:26]
        reg_uop_imm <= 32'h0;
      end else begin
        reg_uop_imm <= io_in_uop_imm;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      reg_uop_dw <= 1'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_flush) begin // @[DataType.scala 40:26]
        reg_uop_dw <= 1'h0;
      end else begin
        reg_uop_dw <= io_in_uop_dw;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      reg_rs1_data <= 64'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_flush) begin // @[DataType.scala 40:26]
        reg_rs1_data <= 64'h0;
      end else begin
        reg_rs1_data <= io_in_rs1_data;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      reg_rs2_data <= 64'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_flush) begin // @[DataType.scala 40:26]
        reg_rs2_data <= 64'h0;
      end else begin
        reg_rs2_data <= io_in_rs2_data;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      reg_rs2_data_from_rf <= 64'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_flush) begin // @[DataType.scala 40:26]
        reg_rs2_data_from_rf <= 64'h0;
      end else begin
        reg_rs2_data_from_rf <= io_in_rs2_data_from_rf;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      reg_bp_npc <= 64'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_flush) begin // @[DataType.scala 40:26]
        reg_bp_npc <= 64'h0;
      end else begin
        reg_bp_npc <= io_in_bp_npc;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_uop_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  reg_uop_exc = _RAND_1[2:0];
  _RAND_2 = {2{`RANDOM}};
  reg_uop_pc = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  reg_uop_npc = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  reg_uop_instr = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  reg_uop_fu = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  reg_uop_alu_op = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  reg_uop_jmp_op = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  reg_uop_mdu_op = _RAND_8[3:0];
  _RAND_9 = {1{`RANDOM}};
  reg_uop_lsu_op = _RAND_9[4:0];
  _RAND_10 = {1{`RANDOM}};
  reg_uop_mem_len = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  reg_uop_csr_op = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  reg_uop_sys_op = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  reg_uop_rd_index = _RAND_13[4:0];
  _RAND_14 = {1{`RANDOM}};
  reg_uop_rd_wen = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  reg_uop_imm = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  reg_uop_dw = _RAND_16[0:0];
  _RAND_17 = {2{`RANDOM}};
  reg_rs1_data = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  reg_rs2_data = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  reg_rs2_data_from_rf = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  reg_bp_npc = _RAND_20[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ALU(
  input  [3:0]  io_uop_alu_op,
  input  [1:0]  io_uop_jmp_op,
  input         io_uop_dw,
  input  [63:0] io_in1,
  input  [63:0] io_in2,
  output [63:0] io_out,
  output [63:0] io_adder_out,
  output        io_cmp_out
);
  wire  is_sub = io_uop_alu_op[3]; // @[ALU.scala 19:24]
  wire  is_cmp = io_uop_alu_op >= 4'hc; // @[ALU.scala 20:25]
  wire  cmp_unsigned = io_uop_alu_op[1]; // @[ALU.scala 21:24]
  wire  cmp_inverted = io_uop_alu_op[0]; // @[ALU.scala 22:24]
  wire  cmp_eq = ~is_sub; // @[ALU.scala 23:22]
  wire [63:0] _in2_inv_T = ~io_in2; // @[ALU.scala 26:34]
  wire [63:0] in2_inv = is_sub ? _in2_inv_T : io_in2; // @[ALU.scala 26:24]
  wire [63:0] in1_xor_in2 = io_in1 ^ in2_inv; // @[ALU.scala 27:28]
  wire [63:0] _io_adder_out_T_1 = io_in1 + in2_inv; // @[ALU.scala 28:26]
  wire [63:0] _GEN_1 = {{63'd0}, is_sub}; // @[ALU.scala 28:36]
  wire  _slt_T_2 = io_in1[63] == io_in2[63]; // @[ALU.scala 32:22]
  wire  _slt_T_6 = cmp_unsigned ? io_in2[63] : io_in1[63]; // @[ALU.scala 34:8]
  wire  slt = _slt_T_2 ? io_adder_out[63] : _slt_T_6; // @[ALU.scala 31:16]
  wire  _io_cmp_out_T_1 = cmp_eq ? in1_xor_in2 == 64'h0 : slt; // @[ALU.scala 36:35]
  wire  _T_1 = is_sub & io_in1[31]; // @[ALU.scala 43:40]
  wire [31:0] _T_3 = _T_1 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [31:0] _T_5 = io_uop_dw ? io_in1[63:32] : _T_3; // @[ALU.scala 44:27]
  wire  _T_7 = io_in2[5] & io_uop_dw; // @[ALU.scala 45:38]
  wire [5:0] shamt = {_T_7,io_in2[4:0]}; // @[Cat.scala 33:92]
  wire [63:0] shin_r = {_T_5,io_in1[31:0]}; // @[Cat.scala 33:92]
  wire  _shin_T_2 = io_uop_alu_op == 4'h5 | io_uop_alu_op == 4'hb; // @[ALU.scala 48:43]
  wire [63:0] _GEN_2 = {{32'd0}, shin_r[63:32]}; // @[Bitwise.scala 108:31]
  wire [63:0] _shin_T_6 = _GEN_2 & 64'hffffffff; // @[Bitwise.scala 108:31]
  wire [63:0] _shin_T_8 = {shin_r[31:0], 32'h0}; // @[Bitwise.scala 108:70]
  wire [63:0] _shin_T_10 = _shin_T_8 & 64'hffffffff00000000; // @[Bitwise.scala 108:80]
  wire [63:0] _shin_T_11 = _shin_T_6 | _shin_T_10; // @[Bitwise.scala 108:39]
  wire [63:0] _GEN_3 = {{16'd0}, _shin_T_11[63:16]}; // @[Bitwise.scala 108:31]
  wire [63:0] _shin_T_16 = _GEN_3 & 64'hffff0000ffff; // @[Bitwise.scala 108:31]
  wire [63:0] _shin_T_18 = {_shin_T_11[47:0], 16'h0}; // @[Bitwise.scala 108:70]
  wire [63:0] _shin_T_20 = _shin_T_18 & 64'hffff0000ffff0000; // @[Bitwise.scala 108:80]
  wire [63:0] _shin_T_21 = _shin_T_16 | _shin_T_20; // @[Bitwise.scala 108:39]
  wire [63:0] _GEN_4 = {{8'd0}, _shin_T_21[63:8]}; // @[Bitwise.scala 108:31]
  wire [63:0] _shin_T_26 = _GEN_4 & 64'hff00ff00ff00ff; // @[Bitwise.scala 108:31]
  wire [63:0] _shin_T_28 = {_shin_T_21[55:0], 8'h0}; // @[Bitwise.scala 108:70]
  wire [63:0] _shin_T_30 = _shin_T_28 & 64'hff00ff00ff00ff00; // @[Bitwise.scala 108:80]
  wire [63:0] _shin_T_31 = _shin_T_26 | _shin_T_30; // @[Bitwise.scala 108:39]
  wire [63:0] _GEN_5 = {{4'd0}, _shin_T_31[63:4]}; // @[Bitwise.scala 108:31]
  wire [63:0] _shin_T_36 = _GEN_5 & 64'hf0f0f0f0f0f0f0f; // @[Bitwise.scala 108:31]
  wire [63:0] _shin_T_38 = {_shin_T_31[59:0], 4'h0}; // @[Bitwise.scala 108:70]
  wire [63:0] _shin_T_40 = _shin_T_38 & 64'hf0f0f0f0f0f0f0f0; // @[Bitwise.scala 108:80]
  wire [63:0] _shin_T_41 = _shin_T_36 | _shin_T_40; // @[Bitwise.scala 108:39]
  wire [63:0] _GEN_6 = {{2'd0}, _shin_T_41[63:2]}; // @[Bitwise.scala 108:31]
  wire [63:0] _shin_T_46 = _GEN_6 & 64'h3333333333333333; // @[Bitwise.scala 108:31]
  wire [63:0] _shin_T_48 = {_shin_T_41[61:0], 2'h0}; // @[Bitwise.scala 108:70]
  wire [63:0] _shin_T_50 = _shin_T_48 & 64'hcccccccccccccccc; // @[Bitwise.scala 108:80]
  wire [63:0] _shin_T_51 = _shin_T_46 | _shin_T_50; // @[Bitwise.scala 108:39]
  wire [63:0] _GEN_7 = {{1'd0}, _shin_T_51[63:1]}; // @[Bitwise.scala 108:31]
  wire [63:0] _shin_T_56 = _GEN_7 & 64'h5555555555555555; // @[Bitwise.scala 108:31]
  wire [63:0] _shin_T_58 = {_shin_T_51[62:0], 1'h0}; // @[Bitwise.scala 108:70]
  wire [63:0] _shin_T_60 = _shin_T_58 & 64'haaaaaaaaaaaaaaaa; // @[Bitwise.scala 108:80]
  wire [63:0] _shin_T_61 = _shin_T_56 | _shin_T_60; // @[Bitwise.scala 108:39]
  wire [63:0] shin = io_uop_alu_op == 4'h5 | io_uop_alu_op == 4'hb ? shin_r : _shin_T_61; // @[ALU.scala 48:20]
  wire  _shout_r_T_1 = is_sub & shin[63]; // @[ALU.scala 49:29]
  wire [64:0] _shout_r_T_3 = {_shout_r_T_1,shin}; // @[ALU.scala 49:53]
  wire [64:0] _shout_r_T_4 = $signed(_shout_r_T_3) >>> shamt; // @[ALU.scala 49:60]
  wire [63:0] shout_r = _shout_r_T_4[63:0]; // @[ALU.scala 49:69]
  wire [63:0] _GEN_8 = {{32'd0}, shout_r[63:32]}; // @[Bitwise.scala 108:31]
  wire [63:0] _shout_l_T_3 = _GEN_8 & 64'hffffffff; // @[Bitwise.scala 108:31]
  wire [63:0] _shout_l_T_5 = {shout_r[31:0], 32'h0}; // @[Bitwise.scala 108:70]
  wire [63:0] _shout_l_T_7 = _shout_l_T_5 & 64'hffffffff00000000; // @[Bitwise.scala 108:80]
  wire [63:0] _shout_l_T_8 = _shout_l_T_3 | _shout_l_T_7; // @[Bitwise.scala 108:39]
  wire [63:0] _GEN_9 = {{16'd0}, _shout_l_T_8[63:16]}; // @[Bitwise.scala 108:31]
  wire [63:0] _shout_l_T_13 = _GEN_9 & 64'hffff0000ffff; // @[Bitwise.scala 108:31]
  wire [63:0] _shout_l_T_15 = {_shout_l_T_8[47:0], 16'h0}; // @[Bitwise.scala 108:70]
  wire [63:0] _shout_l_T_17 = _shout_l_T_15 & 64'hffff0000ffff0000; // @[Bitwise.scala 108:80]
  wire [63:0] _shout_l_T_18 = _shout_l_T_13 | _shout_l_T_17; // @[Bitwise.scala 108:39]
  wire [63:0] _GEN_10 = {{8'd0}, _shout_l_T_18[63:8]}; // @[Bitwise.scala 108:31]
  wire [63:0] _shout_l_T_23 = _GEN_10 & 64'hff00ff00ff00ff; // @[Bitwise.scala 108:31]
  wire [63:0] _shout_l_T_25 = {_shout_l_T_18[55:0], 8'h0}; // @[Bitwise.scala 108:70]
  wire [63:0] _shout_l_T_27 = _shout_l_T_25 & 64'hff00ff00ff00ff00; // @[Bitwise.scala 108:80]
  wire [63:0] _shout_l_T_28 = _shout_l_T_23 | _shout_l_T_27; // @[Bitwise.scala 108:39]
  wire [63:0] _GEN_11 = {{4'd0}, _shout_l_T_28[63:4]}; // @[Bitwise.scala 108:31]
  wire [63:0] _shout_l_T_33 = _GEN_11 & 64'hf0f0f0f0f0f0f0f; // @[Bitwise.scala 108:31]
  wire [63:0] _shout_l_T_35 = {_shout_l_T_28[59:0], 4'h0}; // @[Bitwise.scala 108:70]
  wire [63:0] _shout_l_T_37 = _shout_l_T_35 & 64'hf0f0f0f0f0f0f0f0; // @[Bitwise.scala 108:80]
  wire [63:0] _shout_l_T_38 = _shout_l_T_33 | _shout_l_T_37; // @[Bitwise.scala 108:39]
  wire [63:0] _GEN_12 = {{2'd0}, _shout_l_T_38[63:2]}; // @[Bitwise.scala 108:31]
  wire [63:0] _shout_l_T_43 = _GEN_12 & 64'h3333333333333333; // @[Bitwise.scala 108:31]
  wire [63:0] _shout_l_T_45 = {_shout_l_T_38[61:0], 2'h0}; // @[Bitwise.scala 108:70]
  wire [63:0] _shout_l_T_47 = _shout_l_T_45 & 64'hcccccccccccccccc; // @[Bitwise.scala 108:80]
  wire [63:0] _shout_l_T_48 = _shout_l_T_43 | _shout_l_T_47; // @[Bitwise.scala 108:39]
  wire [63:0] _GEN_13 = {{1'd0}, _shout_l_T_48[63:1]}; // @[Bitwise.scala 108:31]
  wire [63:0] _shout_l_T_53 = _GEN_13 & 64'h5555555555555555; // @[Bitwise.scala 108:31]
  wire [63:0] _shout_l_T_55 = {_shout_l_T_48[62:0], 1'h0}; // @[Bitwise.scala 108:70]
  wire [63:0] _shout_l_T_57 = _shout_l_T_55 & 64'haaaaaaaaaaaaaaaa; // @[Bitwise.scala 108:80]
  wire [63:0] shout_l = _shout_l_T_53 | _shout_l_T_57; // @[Bitwise.scala 108:39]
  wire [63:0] _shout_T_3 = _shin_T_2 ? shout_r : 64'h0; // @[ALU.scala 51:18]
  wire [63:0] _shout_T_5 = io_uop_alu_op == 4'h1 ? shout_l : 64'h0; // @[ALU.scala 52:8]
  wire [63:0] shout = _shout_T_3 | _shout_T_5; // @[ALU.scala 51:81]
  wire  _logic_T_1 = io_uop_alu_op == 4'h6; // @[ALU.scala 55:47]
  wire [63:0] _logic_T_3 = io_uop_alu_op == 4'h4 | io_uop_alu_op == 4'h6 ? in1_xor_in2 : 64'h0; // @[ALU.scala 55:18]
  wire [63:0] _logic_T_7 = io_in1 & io_in2; // @[ALU.scala 56:63]
  wire [63:0] _logic_T_8 = _logic_T_1 | io_uop_alu_op == 4'h7 ? _logic_T_7 : 64'h0; // @[ALU.scala 56:8]
  wire [63:0] logic_ = _logic_T_3 | _logic_T_8; // @[ALU.scala 55:84]
  wire  _shift_logic_T = is_cmp & slt; // @[ALU.scala 57:29]
  wire [63:0] _GEN_14 = {{63'd0}, _shift_logic_T}; // @[ALU.scala 57:37]
  wire [63:0] _shift_logic_T_1 = _GEN_14 | logic_; // @[ALU.scala 57:37]
  wire [63:0] shift_logic = _shift_logic_T_1 | shout; // @[ALU.scala 57:45]
  wire [63:0] out = io_uop_alu_op == 4'h0 | io_uop_alu_op == 4'ha ? io_adder_out : shift_logic; // @[ALU.scala 58:24]
  wire [31:0] _io_out_T_2 = out[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _io_out_T_4 = {_io_out_T_2,out[31:0]}; // @[Cat.scala 33:92]
  assign io_out = ~io_uop_dw ? _io_out_T_4 : out; // @[ALU.scala 60:10 63:{22,31}]
  assign io_adder_out = _io_adder_out_T_1 + _GEN_1; // @[ALU.scala 28:36]
  assign io_cmp_out = cmp_inverted ^ _io_cmp_out_T_1; // @[ALU.scala 36:30]
endmodule
module LSU(
  input         clock,
  input         reset,
  input  [4:0]  io_uop_lsu_op,
  input  [1:0]  io_uop_mem_len,
  input         io_is_mem,
  input         io_is_store,
  input         io_is_amo,
  input  [63:0] io_addr,
  input  [63:0] io_wdata,
  output [63:0] io_rdata,
  output        io_valid,
  output [3:0]  io_exc_code,
  input         io_dmem_req_ready,
  output        io_dmem_req_valid,
  output [38:0] io_dmem_req_bits_addr,
  output [63:0] io_dmem_req_bits_wdata,
  output [7:0]  io_dmem_req_bits_wmask,
  output        io_dmem_req_bits_wen,
  output [1:0]  io_dmem_req_bits_len,
  output        io_dmem_req_bits_lrsc,
  output [4:0]  io_dmem_req_bits_amo,
  output        io_dmem_resp_ready,
  input         io_dmem_resp_valid,
  input  [63:0] io_dmem_resp_bits_rdata,
  input         io_dmem_resp_bits_page_fault,
  input         io_dmem_resp_bits_access_fault,
  output        io_ready
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[LSU.scala 31:58]
  wire [2:0] addr_offset = io_addr[2:0]; // @[LSU.scala 33:28]
  wire [5:0] _wdata_T = {addr_offset, 3'h0}; // @[LSU.scala 35:41]
  wire [126:0] _GEN_7 = {{63'd0}, io_wdata}; // @[LSU.scala 35:25]
  wire [126:0] _wdata_T_1 = _GEN_7 << _wdata_T; // @[LSU.scala 35:25]
  wire [7:0] _wmask_T_1 = 2'h1 == io_uop_mem_len ? 8'h3 : 8'h1; // @[Mux.scala 81:58]
  wire [7:0] _wmask_T_3 = 2'h2 == io_uop_mem_len ? 8'hf : _wmask_T_1; // @[Mux.scala 81:58]
  wire [7:0] _wmask_T_5 = 2'h3 == io_uop_mem_len ? 8'hff : _wmask_T_3; // @[Mux.scala 81:58]
  wire [14:0] _GEN_8 = {{7'd0}, _wmask_T_5}; // @[LSU.scala 45:5]
  wire [14:0] _wmask_T_6 = _GEN_8 << addr_offset; // @[LSU.scala 45:5]
  wire  _io_dmem_req_bits_wen_T = io_is_store | io_is_amo; // @[LSU.scala 51:33]
  wire  _io_dmem_req_bits_lrsc_T_2 = ~io_uop_lsu_op[4]; // @[Constant.scala 85:32]
  wire  _io_dmem_resp_ready_T = state == 2'h2; // @[LSU.scala 55:28]
  wire  _misaligned_T_3 = io_addr[1:0] != 2'h0; // @[LSU.scala 63:42]
  wire  _misaligned_T_5 = addr_offset != 3'h0; // @[LSU.scala 64:42]
  wire  _misaligned_T_9 = 2'h2 == io_uop_mem_len ? _misaligned_T_3 : 2'h1 == io_uop_mem_len & io_addr[0]; // @[Mux.scala 81:58]
  wire  misaligned = 2'h3 == io_uop_mem_len ? _misaligned_T_5 : _misaligned_T_9; // @[Mux.scala 81:58]
  wire  _T_2 = io_dmem_req_ready & io_dmem_req_valid; // @[Decoupled.scala 51:35]
  wire  _T_4 = io_dmem_resp_ready & io_dmem_resp_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _state_T_2 = io_dmem_resp_bits_page_fault | io_dmem_resp_bits_access_fault ? 2'h3 : 2'h0; // @[LSU.scala 81:21]
  wire [1:0] _GEN_2 = _T_4 ? _state_T_2 : state; // @[LSU.scala 80:23 81:15 31:58]
  wire [1:0] _GEN_3 = 2'h3 == state ? 2'h0 : state; // @[LSU.scala 68:17 85:13 31:58]
  wire [63:0] resp_data = io_dmem_resp_bits_rdata >> _wdata_T; // @[LSU.scala 89:35]
  wire  _sign_T_5 = _io_dmem_req_bits_lrsc_T_2 & io_uop_lsu_op[1]; // @[Constant.scala 83:45]
  wire  _sign_T_8 = _sign_T_5 & io_uop_lsu_op[2]; // @[Constant.scala 84:42]
  wire  _sign_T_16 = 2'h1 == io_uop_mem_len ? resp_data[15] : 2'h0 == io_uop_mem_len & resp_data[7]; // @[Mux.scala 81:58]
  wire  _sign_T_18 = 2'h2 == io_uop_mem_len ? resp_data[31] : _sign_T_16; // @[Mux.scala 81:58]
  wire  sign = ~_sign_T_8 & _sign_T_18; // @[LSU.scala 90:37]
  wire [55:0] _rdata_T_1 = sign ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _rdata_T_3 = {_rdata_T_1,resp_data[7:0]}; // @[Cat.scala 33:92]
  wire [47:0] _rdata_T_5 = sign ? 48'hffffffffffff : 48'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _rdata_T_7 = {_rdata_T_5,resp_data[15:0]}; // @[Cat.scala 33:92]
  wire [31:0] _rdata_T_9 = sign ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _rdata_T_11 = {_rdata_T_9,resp_data[31:0]}; // @[Cat.scala 33:92]
  wire [63:0] _rdata_T_13 = 2'h1 == io_uop_mem_len ? _rdata_T_7 : _rdata_T_3; // @[Mux.scala 81:58]
  wire [63:0] _rdata_T_15 = 2'h2 == io_uop_mem_len ? _rdata_T_11 : _rdata_T_13; // @[Mux.scala 81:58]
  wire  _io_valid_T_7 = state == 2'h3; // @[LSU.scala 111:115]
  reg  exc_code_REG; // @[LSU.scala 131:20]
  wire [3:0] _exc_code_T_1 = exc_code_REG ? 4'h7 : 4'hf; // @[LSU.scala 131:12]
  wire [3:0] _exc_code_T_2 = misaligned ? 4'h6 : _exc_code_T_1; // @[LSU.scala 128:10]
  reg  exc_code_REG_1; // @[LSU.scala 136:20]
  wire [3:0] _exc_code_T_3 = exc_code_REG_1 ? 4'h5 : 4'hd; // @[LSU.scala 136:12]
  wire [3:0] _exc_code_T_4 = misaligned ? 4'h4 : _exc_code_T_3; // @[LSU.scala 133:10]
  wire [3:0] exc_code = _io_dmem_req_bits_wen_T ? _exc_code_T_2 : _exc_code_T_4; // @[LSU.scala 126:8]
  assign io_rdata = 2'h3 == io_uop_mem_len ? resp_data : _rdata_T_15; // @[Mux.scala 81:58]
  assign io_valid = _io_dmem_resp_ready_T & (_T_4 & ~io_dmem_resp_bits_page_fault & ~io_dmem_resp_bits_access_fault) |
    state == 2'h3; // @[LSU.scala 111:105]
  assign io_exc_code = _io_valid_T_7 ? exc_code : 4'h0; // @[LSU.scala 139:21]
  assign io_dmem_req_valid = state == 2'h1; // @[LSU.scala 54:28]
  assign io_dmem_req_bits_addr = io_addr[38:0]; // @[LSU.scala 47:18]
  assign io_dmem_req_bits_wdata = _wdata_T_1[63:0]; // @[LSU.scala 35:47]
  assign io_dmem_req_bits_wmask = _wmask_T_6[7:0]; // @[LSU.scala 45:20]
  assign io_dmem_req_bits_wen = io_is_store | io_is_amo; // @[LSU.scala 51:33]
  assign io_dmem_req_bits_len = io_uop_mem_len; // @[LSU.scala 50:18]
  assign io_dmem_req_bits_lrsc = ~io_uop_lsu_op[4] & io_uop_lsu_op[3]; // @[Constant.scala 85:45]
  assign io_dmem_req_bits_amo = io_uop_lsu_op; // @[LSU.scala 53:18]
  assign io_dmem_resp_ready = state == 2'h2; // @[LSU.scala 55:28]
  assign io_ready = state == 2'h0 & ~io_is_mem | io_valid; // @[LSU.scala 113:52]
  always @(posedge clock) begin
    if (reset) begin // @[LSU.scala 31:58]
      state <= 2'h0; // @[LSU.scala 31:58]
    end else if (2'h0 == state) begin // @[LSU.scala 68:17]
      if (io_is_mem) begin // @[LSU.scala 70:23]
        if (misaligned) begin // @[LSU.scala 71:21]
          state <= 2'h3;
        end else begin
          state <= 2'h1;
        end
      end
    end else if (2'h1 == state) begin // @[LSU.scala 68:17]
      if (_T_2) begin // @[LSU.scala 75:22]
        state <= 2'h2; // @[LSU.scala 76:15]
      end
    end else if (2'h2 == state) begin // @[LSU.scala 68:17]
      state <= _GEN_2;
    end else begin
      state <= _GEN_3;
    end
    exc_code_REG <= io_dmem_resp_bits_access_fault; // @[LSU.scala 131:20]
    exc_code_REG_1 <= io_dmem_resp_bits_access_fault; // @[LSU.scala 136:20]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  exc_code_REG = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  exc_code_REG_1 = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MulDiv(
  input         clock,
  input         reset,
  output        io_req_ready,
  input         io_req_valid,
  input  [3:0]  io_req_bits_fn,
  input         io_req_bits_dw,
  input  [63:0] io_req_bits_in1,
  input  [63:0] io_req_bits_in2,
  input         io_resp_ready,
  output        io_resp_valid,
  output [63:0] io_resp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [95:0] _RAND_6;
  reg [159:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] state; // @[Multiplier.scala 48:22]
  reg  req_dw; // @[Multiplier.scala 50:16]
  reg [6:0] count; // @[Multiplier.scala 51:18]
  reg  neg_out; // @[Multiplier.scala 54:20]
  reg  isHi; // @[Multiplier.scala 55:17]
  reg  resHi; // @[Multiplier.scala 56:18]
  reg [64:0] divisor; // @[Multiplier.scala 57:20]
  reg [129:0] remainder; // @[Multiplier.scala 58:22]
  wire [2:0] decoded_plaInput = io_req_bits_fn[2:0]; // @[decoder.scala 40:16 pla.scala 77:22]
  wire [2:0] decoded_invInputs = ~decoded_plaInput; // @[pla.scala 78:21]
  wire  decoded_andMatrixInput_0 = decoded_invInputs[0]; // @[pla.scala 91:29]
  wire  _decoded_T = &decoded_andMatrixInput_0; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_0_1 = decoded_invInputs[2]; // @[pla.scala 91:29]
  wire  _decoded_T_1 = &decoded_andMatrixInput_0_1; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_0_2 = decoded_invInputs[1]; // @[pla.scala 91:29]
  wire [1:0] _decoded_T_2 = {decoded_andMatrixInput_0_2,decoded_andMatrixInput_0_1}; // @[Cat.scala 33:92]
  wire  _decoded_T_3 = &_decoded_T_2; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_0_3 = decoded_plaInput[0]; // @[pla.scala 90:45]
  wire [1:0] _decoded_T_4 = {decoded_andMatrixInput_0_3,decoded_andMatrixInput_0_1}; // @[Cat.scala 33:92]
  wire  _decoded_T_5 = &_decoded_T_4; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_0_4 = decoded_plaInput[1]; // @[pla.scala 90:45]
  wire  _decoded_T_6 = &decoded_andMatrixInput_0_4; // @[pla.scala 98:74]
  wire  decoded_andMatrixInput_1_2 = decoded_plaInput[2]; // @[pla.scala 90:45]
  wire [1:0] _decoded_T_7 = {decoded_andMatrixInput_0,decoded_andMatrixInput_1_2}; // @[Cat.scala 33:92]
  wire  _decoded_T_8 = &_decoded_T_7; // @[pla.scala 98:74]
  wire [1:0] _decoded_orMatrixOutputs_T = {_decoded_T_3,_decoded_T_8}; // @[Cat.scala 33:92]
  wire  _decoded_orMatrixOutputs_T_1 = |_decoded_orMatrixOutputs_T; // @[pla.scala 114:39]
  wire [1:0] _decoded_orMatrixOutputs_T_2 = {_decoded_T,_decoded_T_3}; // @[Cat.scala 33:92]
  wire  _decoded_orMatrixOutputs_T_3 = |_decoded_orMatrixOutputs_T_2; // @[pla.scala 114:39]
  wire [1:0] _decoded_orMatrixOutputs_T_4 = {_decoded_T_5,_decoded_T_6}; // @[Cat.scala 33:92]
  wire  _decoded_orMatrixOutputs_T_5 = |_decoded_orMatrixOutputs_T_4; // @[pla.scala 114:39]
  wire  _decoded_orMatrixOutputs_T_6 = |_decoded_T_1; // @[pla.scala 114:39]
  wire [3:0] decoded_orMatrixOutputs = {_decoded_orMatrixOutputs_T_6,_decoded_orMatrixOutputs_T_5,
    _decoded_orMatrixOutputs_T_3,_decoded_orMatrixOutputs_T_1}; // @[Cat.scala 33:92]
  wire [3:0] decoded_invMatrixOutputs = {decoded_orMatrixOutputs[3],decoded_orMatrixOutputs[2],decoded_orMatrixOutputs[1
    ],decoded_orMatrixOutputs[0]}; // @[Cat.scala 33:92]
  wire  cmdMul = decoded_invMatrixOutputs[3]; // @[Decode.scala 50:77]
  wire  cmdHi = decoded_invMatrixOutputs[2]; // @[Decode.scala 50:77]
  wire  lhsSigned = decoded_invMatrixOutputs[1]; // @[Decode.scala 50:77]
  wire  rhsSigned = decoded_invMatrixOutputs[0]; // @[Decode.scala 50:77]
  wire  _T_4 = ~io_req_bits_dw; // @[Multiplier.scala 75:60]
  wire  _sign_T_2 = _T_4 ? io_req_bits_in1[31] : io_req_bits_in1[63]; // @[Multiplier.scala 78:29]
  wire  lhs_sign = lhsSigned & _sign_T_2; // @[Multiplier.scala 78:23]
  wire [31:0] _hi_T_1 = lhs_sign ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [31:0] hi = _T_4 ? _hi_T_1 : io_req_bits_in1[63:32]; // @[Multiplier.scala 79:17]
  wire [63:0] lhs_in = {hi,io_req_bits_in1[31:0]}; // @[Cat.scala 33:92]
  wire  _sign_T_5 = _T_4 ? io_req_bits_in2[31] : io_req_bits_in2[63]; // @[Multiplier.scala 78:29]
  wire  rhs_sign = rhsSigned & _sign_T_5; // @[Multiplier.scala 78:23]
  wire [31:0] _hi_T_4 = rhs_sign ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [31:0] hi_1 = _T_4 ? _hi_T_4 : io_req_bits_in2[63:32]; // @[Multiplier.scala 79:17]
  wire [64:0] subtractor = remainder[128:64] - divisor; // @[Multiplier.scala 85:37]
  wire [63:0] result = resHi ? remainder[128:65] : remainder[63:0]; // @[Multiplier.scala 86:19]
  wire [63:0] negated_remainder = 64'h0 - result; // @[Multiplier.scala 87:27]
  wire [129:0] _GEN_0 = remainder[63] ? {{66'd0}, negated_remainder} : remainder; // @[Multiplier.scala 90:27 91:17 58:22]
  wire [129:0] _GEN_2 = state == 3'h1 ? _GEN_0 : remainder; // @[Multiplier.scala 58:22 89:57]
  wire [2:0] _GEN_4 = state == 3'h1 ? 3'h3 : state; // @[Multiplier.scala 89:57 96:11 48:22]
  wire [2:0] _GEN_6 = state == 3'h5 ? 3'h7 : _GEN_4; // @[Multiplier.scala 100:11 98:57]
  wire  _GEN_7 = state == 3'h5 ? 1'h0 : resHi; // @[Multiplier.scala 101:11 56:18 98:57]
  wire [128:0] mulReg = {remainder[129:65],remainder[63:0]}; // @[Cat.scala 33:92]
  wire  mplierSign = remainder[64]; // @[Multiplier.scala 105:31]
  wire [63:0] mplier = mulReg[63:0]; // @[Multiplier.scala 106:24]
  wire [64:0] accum = mulReg[128:64]; // @[Multiplier.scala 107:37]
  wire [1:0] _prod_T_2 = {mplierSign,mplier[0]}; // @[Multiplier.scala 109:60]
  wire [66:0] _prod_T_3 = $signed(_prod_T_2) * $signed(divisor); // @[Multiplier.scala 109:67]
  wire [66:0] _GEN_35 = {{2{accum[64]}},accum}; // @[Multiplier.scala 109:76]
  wire [66:0] nextMulReg_hi = $signed(_prod_T_3) + $signed(_GEN_35); // @[Cat.scala 33:92]
  wire [129:0] nextMulReg = {nextMulReg_hi,mplier[63:1]}; // @[Cat.scala 33:92]
  wire  nextMplierSign = count == 7'h3e & neg_out; // @[Multiplier.scala 111:61]
  wire  _eOut_T_4 = ~isHi; // @[Multiplier.scala 115:7]
  wire [128:0] nextMulReg1 = {nextMulReg[128:64],nextMulReg[63:0]}; // @[Cat.scala 33:92]
  wire [129:0] _remainder_T_2 = {nextMulReg1[128:64],nextMplierSign,nextMulReg1[63:0]}; // @[Cat.scala 33:92]
  wire [6:0] _count_T_1 = count + 7'h1; // @[Multiplier.scala 120:20]
  wire [2:0] _GEN_8 = count == 7'h3f ? 3'h6 : _GEN_6; // @[Multiplier.scala 121:55 122:13]
  wire  _GEN_9 = count == 7'h3f ? isHi : _GEN_7; // @[Multiplier.scala 121:55 123:13]
  wire [2:0] _GEN_12 = state == 3'h2 ? _GEN_8 : _GEN_6; // @[Multiplier.scala 103:50]
  wire  _GEN_13 = state == 3'h2 ? _GEN_9 : _GEN_7; // @[Multiplier.scala 103:50]
  wire  unrolls_less = subtractor[64]; // @[Multiplier.scala 130:28]
  wire [63:0] _unrolls_T_2 = unrolls_less ? remainder[127:64] : subtractor[63:0]; // @[Multiplier.scala 131:14]
  wire  _unrolls_T_4 = ~unrolls_less; // @[Multiplier.scala 131:67]
  wire [128:0] unrolls_0 = {_unrolls_T_2,remainder[63:0],_unrolls_T_4}; // @[Cat.scala 33:92]
  wire [2:0] _state_T = neg_out ? 3'h5 : 3'h7; // @[Multiplier.scala 136:19]
  wire [2:0] _GEN_14 = count == 7'h40 ? _state_T : _GEN_12; // @[Multiplier.scala 135:42 136:13]
  wire  divby0 = count == 7'h0 & _unrolls_T_4; // @[Multiplier.scala 143:32]
  wire  _T_23 = io_req_ready & io_req_valid; // @[Decoupled.scala 51:35]
  wire [5:0] _count_T_7 = cmdMul & _T_4 ? 6'h20 : 6'h0; // @[Multiplier.scala 165:38]
  wire [64:0] _divisor_T = {rhs_sign,hi_1,io_req_bits_in2[31:0]}; // @[Cat.scala 33:92]
  wire [2:0] _outMul_T_1 = state & 3'h1; // @[Multiplier.scala 172:23]
  wire  outMul = _outMul_T_1 == 3'h0; // @[Multiplier.scala 172:52]
  wire  _loOut_T = ~req_dw; // @[Multiplier.scala 75:60]
  wire [31:0] loOut = _loOut_T & outMul ? result[63:32] : result[31:0]; // @[Multiplier.scala 173:18]
  wire [31:0] _hiOut_T_4 = loOut[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [31:0] hiOut = _loOut_T ? _hiOut_T_4 : result[63:32]; // @[Multiplier.scala 174:18]
  assign io_req_ready = state == 3'h0; // @[Multiplier.scala 179:25]
  assign io_resp_valid = state == 3'h6 | state == 3'h7; // @[Multiplier.scala 178:42]
  assign io_resp_bits_data = {hiOut,loOut}; // @[Cat.scala 33:92]
  always @(posedge clock) begin
    if (reset) begin // @[Multiplier.scala 48:22]
      state <= 3'h0; // @[Multiplier.scala 48:22]
    end else if (_T_23) begin // @[Multiplier.scala 161:24]
      if (cmdMul) begin // @[Multiplier.scala 162:17]
        state <= 3'h2;
      end else if (lhs_sign | rhs_sign) begin // @[Multiplier.scala 162:36]
        state <= 3'h1;
      end else begin
        state <= 3'h3;
      end
    end else if (io_resp_valid) begin // @[Multiplier.scala 158:36]
      state <= 3'h0; // @[Multiplier.scala 159:11]
    end else if (state == 3'h3) begin // @[Multiplier.scala 126:50]
      state <= _GEN_14;
    end else begin
      state <= _GEN_12;
    end
    if (_T_23) begin // @[Multiplier.scala 161:24]
      req_dw <= io_req_bits_dw; // @[Multiplier.scala 169:9]
    end
    if (_T_23) begin // @[Multiplier.scala 161:24]
      count <= {{1'd0}, _count_T_7}; // @[Multiplier.scala 165:11]
    end else if (state == 3'h3) begin // @[Multiplier.scala 126:50]
      count <= _count_T_1; // @[Multiplier.scala 141:11]
    end else if (state == 3'h2) begin // @[Multiplier.scala 103:50]
      count <= _count_T_1; // @[Multiplier.scala 120:11]
    end
    if (_T_23) begin // @[Multiplier.scala 161:24]
      if (cmdHi) begin // @[Multiplier.scala 166:19]
        neg_out <= lhs_sign;
      end else begin
        neg_out <= lhs_sign != rhs_sign;
      end
    end else if (state == 3'h3) begin // @[Multiplier.scala 126:50]
      if (divby0 & _eOut_T_4) begin // @[Multiplier.scala 156:28]
        neg_out <= 1'h0; // @[Multiplier.scala 156:38]
      end
    end
    if (_T_23) begin // @[Multiplier.scala 161:24]
      isHi <= cmdHi; // @[Multiplier.scala 163:10]
    end
    if (_T_23) begin // @[Multiplier.scala 161:24]
      resHi <= 1'h0; // @[Multiplier.scala 164:11]
    end else if (state == 3'h3) begin // @[Multiplier.scala 126:50]
      if (count == 7'h40) begin // @[Multiplier.scala 135:42]
        resHi <= isHi; // @[Multiplier.scala 137:13]
      end else begin
        resHi <= _GEN_13;
      end
    end else begin
      resHi <= _GEN_13;
    end
    if (_T_23) begin // @[Multiplier.scala 161:24]
      divisor <= _divisor_T; // @[Multiplier.scala 167:13]
    end else if (state == 3'h1) begin // @[Multiplier.scala 89:57]
      if (divisor[63]) begin // @[Multiplier.scala 93:25]
        divisor <= subtractor; // @[Multiplier.scala 94:15]
      end
    end
    if (_T_23) begin // @[Multiplier.scala 161:24]
      remainder <= {{66'd0}, lhs_in}; // @[Multiplier.scala 168:15]
    end else if (state == 3'h3) begin // @[Multiplier.scala 126:50]
      remainder <= {{1'd0}, unrolls_0}; // @[Multiplier.scala 134:15]
    end else if (state == 3'h2) begin // @[Multiplier.scala 103:50]
      remainder <= _remainder_T_2; // @[Multiplier.scala 118:15]
    end else if (state == 3'h5) begin // @[Multiplier.scala 98:57]
      remainder <= {{66'd0}, negated_remainder}; // @[Multiplier.scala 99:15]
    end else begin
      remainder <= _GEN_2;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  req_dw = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  count = _RAND_2[6:0];
  _RAND_3 = {1{`RANDOM}};
  neg_out = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  isHi = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  resHi = _RAND_5[0:0];
  _RAND_6 = {3{`RANDOM}};
  divisor = _RAND_6[64:0];
  _RAND_7 = {5{`RANDOM}};
  remainder = _RAND_7[129:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MDU(
  input         clock,
  input         reset,
  input         io_uop_valid,
  input  [3:0]  io_uop_mdu_op,
  input         io_uop_dw,
  input         io_is_mdu,
  input  [63:0] io_in1,
  input  [63:0] io_in2,
  output [63:0] io_out,
  output        io_valid,
  output        io_ready
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  rocket_mdu_clock; // @[MDU.scala 26:26]
  wire  rocket_mdu_reset; // @[MDU.scala 26:26]
  wire  rocket_mdu_io_req_ready; // @[MDU.scala 26:26]
  wire  rocket_mdu_io_req_valid; // @[MDU.scala 26:26]
  wire [3:0] rocket_mdu_io_req_bits_fn; // @[MDU.scala 26:26]
  wire  rocket_mdu_io_req_bits_dw; // @[MDU.scala 26:26]
  wire [63:0] rocket_mdu_io_req_bits_in1; // @[MDU.scala 26:26]
  wire [63:0] rocket_mdu_io_req_bits_in2; // @[MDU.scala 26:26]
  wire  rocket_mdu_io_resp_ready; // @[MDU.scala 26:26]
  wire  rocket_mdu_io_resp_valid; // @[MDU.scala 26:26]
  wire [63:0] rocket_mdu_io_resp_bits_data; // @[MDU.scala 26:26]
  reg [1:0] state; // @[MDU.scala 24:49]
  wire  _T_2 = rocket_mdu_io_req_ready & rocket_mdu_io_req_valid; // @[Decoupled.scala 51:35]
  wire  _T_4 = rocket_mdu_io_resp_ready & rocket_mdu_io_resp_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _GEN_2 = _T_4 ? 2'h0 : state; // @[MDU.scala 48:37 49:15 24:49]
  MulDiv rocket_mdu ( // @[MDU.scala 26:26]
    .clock(rocket_mdu_clock),
    .reset(rocket_mdu_reset),
    .io_req_ready(rocket_mdu_io_req_ready),
    .io_req_valid(rocket_mdu_io_req_valid),
    .io_req_bits_fn(rocket_mdu_io_req_bits_fn),
    .io_req_bits_dw(rocket_mdu_io_req_bits_dw),
    .io_req_bits_in1(rocket_mdu_io_req_bits_in1),
    .io_req_bits_in2(rocket_mdu_io_req_bits_in2),
    .io_resp_ready(rocket_mdu_io_resp_ready),
    .io_resp_valid(rocket_mdu_io_resp_valid),
    .io_resp_bits_data(rocket_mdu_io_resp_bits_data)
  );
  assign io_out = rocket_mdu_io_resp_bits_data; // @[MDU.scala 54:12]
  assign io_valid = state == 2'h2 & _T_4; // @[MDU.scala 55:34]
  assign io_ready = state == 2'h0 & ~io_is_mdu | io_valid; // @[MDU.scala 56:47]
  assign rocket_mdu_clock = clock;
  assign rocket_mdu_reset = reset;
  assign rocket_mdu_io_req_valid = state == 2'h1 & io_uop_valid & io_is_mdu; // @[MDU.scala 27:64]
  assign rocket_mdu_io_req_bits_fn = io_uop_mdu_op; // @[MDU.scala 28:30]
  assign rocket_mdu_io_req_bits_dw = io_uop_dw; // @[MDU.scala 29:30]
  assign rocket_mdu_io_req_bits_in1 = io_in1; // @[MDU.scala 30:30]
  assign rocket_mdu_io_req_bits_in2 = io_in2; // @[MDU.scala 31:30]
  assign rocket_mdu_io_resp_ready = 1'h1; // @[MDU.scala 34:30]
  always @(posedge clock) begin
    if (reset) begin // @[MDU.scala 24:49]
      state <= 2'h0; // @[MDU.scala 24:49]
    end else if (2'h0 == state) begin // @[MDU.scala 36:17]
      if (io_is_mdu) begin // @[MDU.scala 38:20]
        state <= 2'h1; // @[MDU.scala 39:15]
      end
    end else if (2'h1 == state) begin // @[MDU.scala 36:17]
      if (_T_2) begin // @[MDU.scala 43:36]
        state <= 2'h2; // @[MDU.scala 44:15]
      end
    end else if (2'h2 == state) begin // @[MDU.scala 36:17]
      state <= _GEN_2;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CSR(
  input         clock,
  input         reset,
  input         io_uop_valid,
  input  [2:0]  io_uop_exc,
  input  [63:0] io_uop_pc,
  input  [63:0] io_uop_npc,
  input  [2:0]  io_uop_fu,
  input  [2:0]  io_uop_sys_op,
  input  [11:0] io_rw_addr,
  input  [1:0]  io_rw_cmd,
  input  [63:0] io_rw_wdata,
  output [63:0] io_rw_rdata,
  output        io_rw_valid,
  output [1:0]  io_prv,
  output        io_mprv,
  output [1:0]  io_mpp,
  output        io_sv39_en,
  output [15:0] io_satp_asid,
  output [43:0] io_satp_ppn,
  output        io_sfence_vma,
  output        io_fence_i,
  output        io_jmp_packet_valid,
  output [63:0] io_jmp_packet_target,
  input  [63:0] io_lsu_addr,
  input  [3:0]  io_lsu_exc_code,
  input         io_interrupt_mtip,
  input         io_interrupt_msip,
  input         io_interrupt_meip,
  input         io_interrupt_seip,
  output        io_is_int,
  input         io_commit
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] prv; // @[CSR.scala 49:26]
  wire  mret_legal = prv == 2'h3; // @[CSR.scala 50:24]
  wire  prv_is_s = prv == 2'h1; // @[CSR.scala 51:24]
  wire  prv_is_ms = mret_legal | prv_is_s; // @[CSR.scala 52:28]
  wire  prv_is_u = prv == 2'h0; // @[CSR.scala 53:24]
  wire  _wen_T = io_rw_cmd != 2'h0; // @[CSR.scala 58:30]
  reg [63:0] mcounteren; // @[CSR.scala 477:27]
  reg [63:0] scounteren; // @[CSR.scala 208:27]
  reg  mstatus_tvm; // @[CSR.scala 117:29]
  wire  tvm_en = prv_is_s & mstatus_tvm; // @[CSR.scala 285:31]
  wire  _csr_legal_T_1 = prv_is_ms & ~tvm_en; // @[CSR.scala 300:28]
  wire  _GEN_13 = io_rw_addr == 12'h100 & prv_is_ms; // @[CSR.scala 151:39 162:15 55:30]
  wire  _GEN_41 = io_rw_addr == 12'h300 ? mret_legal : _GEN_13; // @[CSR.scala 164:39 182:15]
  wire  _GEN_45 = io_rw_addr == 12'h105 ? prv_is_ms : _GEN_41; // @[CSR.scala 194:37 199:15]
  wire  _GEN_49 = io_rw_addr == 12'h106 ? prv_is_ms : _GEN_45; // @[CSR.scala 209:42 214:15]
  wire  _GEN_53 = io_rw_addr == 12'h140 ? prv_is_ms : _GEN_49; // @[CSR.scala 224:40 229:15]
  wire  _GEN_57 = io_rw_addr == 12'h141 ? prv_is_ms : _GEN_53; // @[CSR.scala 239:36 244:15]
  wire  _GEN_61 = io_rw_addr == 12'h142 ? prv_is_ms : _GEN_57; // @[CSR.scala 254:38 259:15]
  wire  _GEN_65 = io_rw_addr == 12'h143 ? prv_is_ms : _GEN_61; // @[CSR.scala 269:37 274:15]
  wire  _GEN_77 = io_rw_addr == 12'h180 ? prv_is_ms & ~tvm_en : _GEN_65; // @[CSR.scala 291:36 300:15]
  wire  _GEN_79 = io_rw_addr == 12'hf11 ? mret_legal : _GEN_77; // @[CSR.scala 309:41 311:15]
  wire  _GEN_81 = io_rw_addr == 12'hf12 ? mret_legal : _GEN_79; // @[CSR.scala 320:39 322:15]
  wire  _GEN_83 = io_rw_addr == 12'hf13 ? mret_legal : _GEN_81; // @[CSR.scala 331:38 333:15]
  wire  _GEN_89 = io_rw_addr == 12'hf14 ? mret_legal : _GEN_83; // @[CSR.scala 344:39 350:15]
  wire  _GEN_91 = io_rw_addr == 12'h301 ? mret_legal : _GEN_89; // @[CSR.scala 361:36 363:15]
  wire  _GEN_95 = io_rw_addr == 12'h302 ? mret_legal : _GEN_91; // @[CSR.scala 373:39 378:15]
  wire  _GEN_99 = io_rw_addr == 12'h303 ? mret_legal : _GEN_95; // @[CSR.scala 388:39 393:15]
  wire  _GEN_113 = io_rw_addr == 12'h304 ? mret_legal : _GEN_99; // @[CSR.scala 434:35 444:15]
  wire  _GEN_121 = io_rw_addr == 12'h104 ? prv_is_ms : _GEN_113; // @[CSR.scala 446:35 453:15]
  wire  _GEN_125 = io_rw_addr == 12'h305 ? mret_legal : _GEN_121; // @[CSR.scala 463:37 468:15]
  wire  _GEN_129 = io_rw_addr == 12'h306 ? mret_legal : _GEN_125; // @[CSR.scala 478:42 483:15]
  wire  _GEN_133 = io_rw_addr == 12'h340 ? mret_legal : _GEN_129; // @[CSR.scala 493:40 498:15]
  wire  _GEN_137 = io_rw_addr == 12'h341 ? mret_legal : _GEN_133; // @[CSR.scala 508:36 513:15]
  wire  _GEN_141 = io_rw_addr == 12'h342 ? mret_legal : _GEN_137; // @[CSR.scala 523:38 528:15]
  wire  _GEN_145 = io_rw_addr == 12'h343 ? mret_legal : _GEN_141; // @[CSR.scala 538:37 543:15]
  wire  _GEN_153 = io_rw_addr == 12'h344 ? mret_legal : _GEN_145; // @[CSR.scala 585:35 592:15]
  wire  _GEN_157 = io_rw_addr == 12'h144 ? prv_is_ms : _GEN_153; // @[CSR.scala 594:35 599:15]
  wire  _GEN_161 = io_rw_addr == 12'hb00 ? mret_legal : _GEN_157; // @[CSR.scala 610:38 615:15]
  wire  _GEN_163 = io_rw_addr == 12'hc00 ? mret_legal | prv_is_s & mcounteren[0] | prv_is_u & mcounteren[0] & scounteren
    [0] : _GEN_161; // @[CSR.scala 617:37 619:15]
  wire  _GEN_167 = io_rw_addr == 12'hb02 ? mret_legal : _GEN_163; // @[CSR.scala 632:40 637:15]
  wire  csr_legal = io_rw_addr == 12'hc02 ? mret_legal | prv_is_s & mcounteren[2] | prv_is_u & mcounteren[2] &
    scounteren[2] : _GEN_167; // @[CSR.scala 639:39 641:15]
  wire  wen = io_rw_cmd != 2'h0 & io_uop_exc == 3'h0 & csr_legal; // @[CSR.scala 58:81]
  reg [63:0] instret; // @[CSR.scala 630:24]
  reg [63:0] cycle; // @[CSR.scala 608:22]
  reg  ip_seip_r; // @[CSR.scala 558:26]
  wire  ip_seip = io_interrupt_seip | ip_seip_r; // @[CSR.scala 559:38]
  reg  ip_stip; // @[CSR.scala 556:26]
  reg  ip_ssip; // @[CSR.scala 554:26]
  wire [63:0] sip = {54'h0,ip_seip,3'h0,ip_stip,3'h0,ip_ssip,1'h0}; // @[Cat.scala 33:92]
  wire [5:0] mip_lo = {ip_stip,1'h0,io_interrupt_msip,1'h0,ip_ssip,1'h0}; // @[Cat.scala 33:92]
  wire [63:0] mip = {52'h0,io_interrupt_meip,1'h0,ip_seip,1'h0,io_interrupt_mtip,1'h0,mip_lo}; // @[Cat.scala 33:92]
  reg [63:0] mtval; // @[CSR.scala 537:22]
  reg [63:0] mcause; // @[CSR.scala 522:23]
  reg [63:0] mepc; // @[CSR.scala 507:21]
  reg [63:0] mscratch; // @[CSR.scala 492:25]
  reg [63:0] mtvec; // @[CSR.scala 462:22]
  reg  ie_seie; // @[CSR.scala 408:24]
  reg  ie_stie; // @[CSR.scala 406:24]
  reg  ie_ssie; // @[CSR.scala 404:24]
  wire [63:0] sie = {54'h0,ie_seie,3'h0,ie_stie,3'h0,ie_ssie,1'h0}; // @[Cat.scala 33:92]
  reg  ie_meie; // @[CSR.scala 409:24]
  reg  ie_mtie; // @[CSR.scala 407:24]
  reg  ie_msie; // @[CSR.scala 405:24]
  wire [5:0] mie_lo = {ie_stie,1'h0,ie_msie,1'h0,ie_ssie,1'h0}; // @[Cat.scala 33:92]
  wire [63:0] mie = {52'h0,ie_meie,1'h0,ie_seie,1'h0,ie_mtie,1'h0,mie_lo}; // @[Cat.scala 33:92]
  reg [63:0] mideleg; // @[CSR.scala 387:24]
  reg [63:0] medeleg; // @[CSR.scala 372:24]
  reg [63:0] mhartid; // @[CSR.scala 342:33]
  reg [63:0] satp; // @[CSR.scala 283:29]
  reg [63:0] stval; // @[CSR.scala 268:22]
  reg [63:0] scause; // @[CSR.scala 253:23]
  reg [63:0] sepc; // @[CSR.scala 238:21]
  reg [63:0] sscratch; // @[CSR.scala 223:25]
  reg [63:0] stvec; // @[CSR.scala 193:22]
  reg [1:0] status_fs; // @[CSR.scala 86:28]
  wire  status_sd = |status_fs; // @[CSR.scala 91:31]
  reg  mstatus_tsr; // @[CSR.scala 119:29]
  reg  mstatus_tw; // @[CSR.scala 118:29]
  reg  status_mxr; // @[CSR.scala 89:28]
  reg  status_sum; // @[CSR.scala 88:28]
  reg  mstatus_mprv; // @[CSR.scala 116:29]
  wire [46:0] mstatus_hi = {status_sd,25'h0,2'h0,13'h1400,mstatus_tsr,mstatus_tw,mstatus_tvm,status_mxr,status_sum,
    mstatus_mprv}; // @[Cat.scala 33:92]
  reg [1:0] mstatus_mpp; // @[CSR.scala 115:29]
  reg  status_spp; // @[CSR.scala 84:28]
  reg  mstatus_mpie; // @[CSR.scala 114:29]
  reg  status_spie; // @[CSR.scala 82:28]
  reg  mstatus_mie; // @[CSR.scala 113:29]
  reg  status_sie; // @[CSR.scala 81:28]
  wire [5:0] mstatus_lo_lo = {status_spie,1'h0,mstatus_mie,1'h0,status_sie,1'h0}; // @[Cat.scala 33:92]
  wire [63:0] mstatus = {mstatus_hi,2'h0,status_fs,mstatus_mpp,2'h0,status_spp,mstatus_mpie,1'h0,mstatus_lo_lo}; // @[Cat.scala 33:92]
  wire [12:0] sstatus_lo = {4'h0,status_spp,2'h0,status_spie,3'h0,status_sie,1'h0}; // @[Cat.scala 33:92]
  wire [63:0] sstatus = {status_sd,29'h0,2'h2,12'h0,status_mxr,status_sum,1'h0,2'h0,status_fs,sstatus_lo}; // @[Cat.scala 33:92]
  wire [63:0] _GEN_6 = io_rw_addr == 12'h100 ? sstatus : 64'h0; // @[CSR.scala 151:39 152:11 56:30]
  wire [63:0] _GEN_27 = io_rw_addr == 12'h300 ? mstatus : _GEN_6; // @[CSR.scala 164:39 165:11]
  wire [63:0] _GEN_43 = io_rw_addr == 12'h105 ? stvec : _GEN_27; // @[CSR.scala 194:37 195:11]
  wire [63:0] _GEN_47 = io_rw_addr == 12'h106 ? scounteren : _GEN_43; // @[CSR.scala 209:42 210:11]
  wire [63:0] _GEN_51 = io_rw_addr == 12'h140 ? sscratch : _GEN_47; // @[CSR.scala 224:40 225:11]
  wire [63:0] _GEN_55 = io_rw_addr == 12'h141 ? sepc : _GEN_51; // @[CSR.scala 239:36 240:11]
  wire [63:0] _GEN_59 = io_rw_addr == 12'h142 ? scause : _GEN_55; // @[CSR.scala 254:38 255:11]
  wire [63:0] _GEN_63 = io_rw_addr == 12'h143 ? stval : _GEN_59; // @[CSR.scala 269:37 270:11]
  wire [63:0] _GEN_71 = io_rw_addr == 12'h180 ? satp : _GEN_63; // @[CSR.scala 291:36 292:11]
  wire [63:0] _GEN_78 = io_rw_addr == 12'hf11 ? 64'h0 : _GEN_71; // @[CSR.scala 309:41 310:15]
  wire [63:0] _GEN_80 = io_rw_addr == 12'hf12 ? 64'h0 : _GEN_78; // @[CSR.scala 320:39 321:15]
  wire [63:0] _GEN_82 = io_rw_addr == 12'hf13 ? 64'h0 : _GEN_80; // @[CSR.scala 331:38 332:15]
  wire [63:0] _GEN_86 = io_rw_addr == 12'hf14 ? mhartid : _GEN_82; // @[CSR.scala 344:39 345:11]
  wire [63:0] _GEN_90 = io_rw_addr == 12'h301 ? 64'h8000000000141101 : _GEN_86; // @[CSR.scala 361:36 362:15]
  wire [63:0] _GEN_93 = io_rw_addr == 12'h302 ? medeleg : _GEN_90; // @[CSR.scala 373:39 374:11]
  wire [63:0] _GEN_97 = io_rw_addr == 12'h303 ? mideleg : _GEN_93; // @[CSR.scala 388:39 389:11]
  wire [63:0] _GEN_106 = io_rw_addr == 12'h304 ? mie : _GEN_97; // @[CSR.scala 434:35 435:11]
  wire [63:0] _GEN_117 = io_rw_addr == 12'h104 ? sie : _GEN_106; // @[CSR.scala 446:35 447:11]
  wire [63:0] _GEN_123 = io_rw_addr == 12'h305 ? mtvec : _GEN_117; // @[CSR.scala 463:37 464:11]
  wire [63:0] _GEN_127 = io_rw_addr == 12'h306 ? mcounteren : _GEN_123; // @[CSR.scala 478:42 479:11]
  wire [63:0] _GEN_131 = io_rw_addr == 12'h340 ? mscratch : _GEN_127; // @[CSR.scala 493:40 494:11]
  wire [63:0] _GEN_135 = io_rw_addr == 12'h341 ? mepc : _GEN_131; // @[CSR.scala 508:36 509:11]
  wire [63:0] _GEN_139 = io_rw_addr == 12'h342 ? mcause : _GEN_135; // @[CSR.scala 523:38 524:11]
  wire [63:0] _GEN_143 = io_rw_addr == 12'h343 ? mtval : _GEN_139; // @[CSR.scala 538:37 539:11]
  wire [63:0] _GEN_149 = io_rw_addr == 12'h344 ? mip : _GEN_143; // @[CSR.scala 585:35 586:11]
  wire [63:0] _GEN_155 = io_rw_addr == 12'h144 ? sip : _GEN_149; // @[CSR.scala 594:35 595:11]
  wire [63:0] _GEN_159 = io_rw_addr == 12'hb00 ? cycle : _GEN_155; // @[CSR.scala 610:38 611:11]
  wire [63:0] _GEN_162 = io_rw_addr == 12'hc00 ? cycle : _GEN_159; // @[CSR.scala 617:37 618:15]
  wire [63:0] _GEN_165 = io_rw_addr == 12'hb02 ? instret : _GEN_162; // @[CSR.scala 632:40 633:11]
  wire [63:0] rdata = io_rw_addr == 12'hc02 ? instret : _GEN_165; // @[CSR.scala 639:39 640:15]
  wire [63:0] _wdata_T = rdata | io_rw_wdata; // @[CSR.scala 64:31]
  wire [63:0] _wdata_T_1 = ~io_rw_wdata; // @[CSR.scala 65:33]
  wire [63:0] _wdata_T_2 = rdata & _wdata_T_1; // @[CSR.scala 65:31]
  wire [63:0] _wdata_T_4 = 2'h1 == io_rw_cmd ? io_rw_wdata : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _wdata_T_6 = 2'h2 == io_rw_cmd ? _wdata_T : _wdata_T_4; // @[Mux.scala 81:58]
  wire [63:0] wdata = 2'h3 == io_rw_cmd ? _wdata_T_2 : _wdata_T_6; // @[Mux.scala 81:58]
  wire  _GEN_0 = wen ? wdata[1] : status_sie; // @[CSR.scala 153:15 154:19 81:28]
  wire  _GEN_1 = wen ? wdata[5] : status_spie; // @[CSR.scala 153:15 155:19 82:28]
  wire  _GEN_2 = wen ? wdata[8] : status_spp; // @[CSR.scala 153:15 156:19 84:28]
  wire [1:0] _GEN_3 = wen ? wdata[14:13] : status_fs; // @[CSR.scala 153:15 157:19 86:28]
  wire  _GEN_4 = wen ? wdata[18] : status_sum; // @[CSR.scala 153:15 159:18 88:28]
  wire  _GEN_5 = wen ? wdata[19] : status_mxr; // @[CSR.scala 153:15 160:18 89:28]
  wire  _GEN_7 = io_rw_addr == 12'h100 ? _GEN_0 : status_sie; // @[CSR.scala 151:39 81:28]
  wire  _GEN_8 = io_rw_addr == 12'h100 ? _GEN_1 : status_spie; // @[CSR.scala 151:39 82:28]
  wire  _GEN_9 = io_rw_addr == 12'h100 ? _GEN_2 : status_spp; // @[CSR.scala 151:39 84:28]
  wire [1:0] _GEN_10 = io_rw_addr == 12'h100 ? _GEN_3 : status_fs; // @[CSR.scala 151:39 86:28]
  wire  _GEN_11 = io_rw_addr == 12'h100 ? _GEN_4 : status_sum; // @[CSR.scala 151:39 88:28]
  wire  _GEN_12 = io_rw_addr == 12'h100 ? _GEN_5 : status_mxr; // @[CSR.scala 151:39 89:28]
  wire  _GEN_14 = wen ? wdata[1] : _GEN_7; // @[CSR.scala 166:15 167:19]
  wire  _GEN_15 = wen ? wdata[5] : _GEN_8; // @[CSR.scala 166:15 168:19]
  wire  _GEN_16 = wen ? wdata[8] : _GEN_9; // @[CSR.scala 166:15 169:19]
  wire  _GEN_20 = wen ? wdata[3] : mstatus_mie; // @[CSR.scala 166:15 174:20 113:29]
  wire  _GEN_21 = wen ? wdata[7] : mstatus_mpie; // @[CSR.scala 166:15 175:20 114:29]
  wire [1:0] _GEN_22 = wen ? wdata[12:11] : mstatus_mpp; // @[CSR.scala 166:15 176:20 115:29]
  wire  _GEN_23 = wen ? wdata[17] : mstatus_mprv; // @[CSR.scala 166:15 177:20 116:29]
  wire  _GEN_29 = io_rw_addr == 12'h300 ? _GEN_15 : _GEN_8; // @[CSR.scala 164:39]
  wire  _GEN_30 = io_rw_addr == 12'h300 ? _GEN_16 : _GEN_9; // @[CSR.scala 164:39]
  wire  _GEN_35 = io_rw_addr == 12'h300 ? _GEN_21 : mstatus_mpie; // @[CSR.scala 114:29 164:39]
  wire  _GEN_37 = io_rw_addr == 12'h300 ? _GEN_23 : mstatus_mprv; // @[CSR.scala 116:29 164:39]
  wire  satp_wen = wdata[62:60] == 3'h0; // @[CSR.scala 287:33]
  wire  _GEN_67 = wen & satp_wen ? wdata[63] : satp[63]; // @[CSR.scala 288:16 293:27 295:20]
  wire [15:0] _GEN_68 = wen & satp_wen ? wdata[59:44] : satp[59:44]; // @[CSR.scala 289:16 293:27 296:20]
  wire [43:0] _GEN_69 = wen & satp_wen ? wdata[43:0] : satp[43:0]; // @[CSR.scala 290:16 293:27 297:20]
  wire  _GEN_70 = wen & satp_wen & prv_is_s; // @[CSR.scala 293:27 298:20 284:33]
  wire  satp_updated = io_rw_addr == 12'h180 & _GEN_70; // @[CSR.scala 284:33 291:36]
  reg  mhartid_writable; // @[CSR.scala 343:33]
  wire  _GEN_85 = wen & mhartid_writable ? 1'h0 : mhartid_writable; // @[CSR.scala 346:35 348:24 343:33]
  wire  _GEN_88 = io_rw_addr == 12'hf14 ? _GEN_85 : mhartid_writable; // @[CSR.scala 343:33 344:39]
  wire [63:0] _medeleg_T = wdata & 64'hf7ff; // @[CSR.scala 376:24]
  wire [63:0] _mideleg_T = wdata & 64'h222; // @[CSR.scala 391:24]
  wire  _GEN_100 = wen ? wdata[1] : ie_ssie; // @[CSR.scala 436:15 437:15 404:24]
  wire  _GEN_102 = wen ? wdata[5] : ie_stie; // @[CSR.scala 436:15 439:15 406:24]
  wire  _GEN_104 = wen ? wdata[9] : ie_seie; // @[CSR.scala 436:15 441:15 408:24]
  wire  _GEN_107 = io_rw_addr == 12'h304 ? _GEN_100 : ie_ssie; // @[CSR.scala 404:24 434:35]
  wire  _GEN_109 = io_rw_addr == 12'h304 ? _GEN_102 : ie_stie; // @[CSR.scala 406:24 434:35]
  wire  _GEN_111 = io_rw_addr == 12'h304 ? _GEN_104 : ie_seie; // @[CSR.scala 408:24 434:35]
  wire  _GEN_146 = wen ? wdata[1] : ip_ssip; // @[CSR.scala 587:15 588:17 554:26]
  wire  _GEN_150 = io_rw_addr == 12'h344 ? _GEN_146 : ip_ssip; // @[CSR.scala 554:26 585:35]
  wire [63:0] _cycle_T_1 = cycle + 64'h1; // @[CSR.scala 609:18]
  wire [63:0] _GEN_218 = {{63'd0}, io_commit}; // @[CSR.scala 631:22]
  wire [63:0] _instret_T_1 = instret + _GEN_218; // @[CSR.scala 631:22]
  wire  is_mret = io_uop_sys_op == 3'h1; // @[CSR.scala 656:34]
  wire  _T_32 = is_mret & mret_legal; // @[CSR.scala 658:16]
  wire  _GEN_170 = mstatus_mpp != 2'h3 ? 1'h0 : _GEN_37; // @[CSR.scala 664:35 665:20]
  wire [1:0] _GEN_171 = is_mret & mret_legal ? mstatus_mpp : prv; // @[CSR.scala 658:31 659:18 49:26]
  wire  _GEN_173 = is_mret & mret_legal | _GEN_35; // @[CSR.scala 658:31 662:18]
  wire  _GEN_175 = is_mret & mret_legal ? _GEN_170 : _GEN_37; // @[CSR.scala 658:31]
  wire  is_sret = io_uop_sys_op == 3'h2; // @[CSR.scala 669:34]
  wire  sret_legal = prv_is_ms & ~mstatus_tsr; // @[CSR.scala 670:30]
  wire  _T_34 = is_sret & sret_legal; // @[CSR.scala 671:16]
  wire [1:0] _GEN_219 = {{1'd0}, status_spp}; // @[CSR.scala 677:21]
  wire [1:0] _GEN_177 = is_sret & sret_legal ? {{1'd0}, status_spp} : _GEN_171; // @[CSR.scala 671:31 672:17]
  wire  _GEN_179 = is_sret & sret_legal | _GEN_29; // @[CSR.scala 671:31 675:17]
  wire  _GEN_180 = is_sret & sret_legal ? 1'h0 : _GEN_30; // @[CSR.scala 671:31 676:17]
  wire  is_sfv = io_uop_sys_op == 3'h6 & io_uop_valid; // @[CSR.scala 685:55]
  wire  is_fence_i = io_uop_sys_op == 3'h5 & io_uop_valid; // @[CSR.scala 687:58]
  wire  is_sys = io_sfence_vma | is_fence_i; // @[CSR.scala 688:34]
  wire  is_exc_from_prev = io_uop_exc != 3'h0; // @[CSR.scala 695:38]
  wire  is_exc_from_lsu = io_lsu_exc_code != 4'h0; // @[CSR.scala 696:43]
  wire  is_exc_from_csr = ~csr_legal & _wen_T; // @[CSR.scala 697:37]
  wire  _is_exc_from_sys_T = ~mret_legal; // @[CSR.scala 698:38]
  wire  is_exc_from_sys = is_mret & ~mret_legal | is_sret & ~sret_legal | is_sfv & ~_csr_legal_T_1; // @[CSR.scala 698:79]
  wire  is_exc = is_exc_from_prev | is_exc_from_lsu | is_exc_from_csr; // @[CSR.scala 699:62]
  wire  int_attach = io_uop_valid & (io_uop_fu == 3'h0 | io_uop_fu == 3'h1); // @[CSR.scala 719:37]
  wire [63:0] int_bits = mip & mie; // @[CSR.scala 720:28]
  wire [63:0] _int_bits_mmode_T = ~mideleg; // @[CSR.scala 721:36]
  wire [63:0] int_bits_mmode = int_bits & _int_bits_mmode_T; // @[CSR.scala 721:33]
  wire [3:0] _GEN_182 = int_bits[5] ? 4'h5 : 4'h0; // @[CSR.scala 713:22 702:24 714:9]
  wire [3:0] _GEN_183 = int_bits[1] ? 4'h1 : _GEN_182; // @[CSR.scala 711:22 712:9]
  wire [3:0] _GEN_184 = int_bits[9] ? 4'h9 : _GEN_183; // @[CSR.scala 709:22 710:9]
  wire [3:0] _GEN_185 = int_bits[7] ? 4'h7 : _GEN_184; // @[CSR.scala 707:22 708:9]
  wire [3:0] _GEN_186 = int_bits[3] ? 4'h3 : _GEN_185; // @[CSR.scala 705:22 706:9]
  wire [3:0] int_index_tmp = int_bits[11] ? 4'hb : _GEN_186; // @[CSR.scala 703:17 704:9]
  wire [3:0] _GEN_188 = int_bits_mmode[5] ? 4'h5 : 4'h0; // @[CSR.scala 713:22 702:24 714:9]
  wire [3:0] _GEN_189 = int_bits_mmode[1] ? 4'h1 : _GEN_188; // @[CSR.scala 711:22 712:9]
  wire [3:0] _GEN_190 = int_bits_mmode[9] ? 4'h9 : _GEN_189; // @[CSR.scala 709:22 710:9]
  wire [3:0] _GEN_191 = int_bits_mmode[7] ? 4'h7 : _GEN_190; // @[CSR.scala 707:22 708:9]
  wire [3:0] _GEN_192 = int_bits_mmode[3] ? 4'h3 : _GEN_191; // @[CSR.scala 705:22 706:9]
  wire [3:0] int_index_y = int_bits_mmode[11] ? 4'hb : _GEN_192; // @[CSR.scala 703:17 704:9]
  wire [3:0] _GEN_194 = mstatus_mie ? int_index_y : 4'h0; // @[CSR.scala 726:30 727:17 723:34]
  wire [15:0] _T_38 = 16'h1 << int_index_tmp; // @[CSR.scala 730:16]
  wire [63:0] _GEN_220 = {{48'd0}, _T_38}; // @[CSR.scala 730:34]
  wire [63:0] _T_39 = _GEN_220 & mideleg; // @[CSR.scala 730:34]
  wire [3:0] _GEN_195 = status_sie | prv_is_u ? int_index_tmp : 4'h0; // @[CSR.scala 731:50 732:19 723:34]
  wire [3:0] _GEN_196 = mstatus_mie | prv_is_u | prv_is_s ? int_index_tmp : 4'h0; // @[CSR.scala 735:70 736:19 723:34]
  wire [3:0] _GEN_197 = _T_39 != 64'h0 ? _GEN_195 : _GEN_196; // @[CSR.scala 730:54]
  wire [3:0] int_index = mret_legal ? _GEN_194 : _GEN_197; // @[CSR.scala 725:25]
  wire  is_int = int_attach & int_index != 4'h0; // @[CSR.scala 740:27]
  wire [1:0] _cause_exc_T_2 = is_exc_from_csr | is_exc_from_sys ? 2'h2 : 2'h0; // @[CSR.scala 751:10]
  wire [3:0] _cause_exc_T_3 = is_exc_from_lsu ? io_lsu_exc_code : {{2'd0}, _cause_exc_T_2}; // @[CSR.scala 748:8]
  wire [3:0] _cause_exc_T_4 = {2'h2,prv}; // @[Cat.scala 33:92]
  wire [3:0] _cause_exc_T_6 = 3'h1 == io_uop_exc ? 4'h0 : _cause_exc_T_3; // @[Mux.scala 81:58]
  wire [3:0] _cause_exc_T_8 = 3'h2 == io_uop_exc ? 4'h1 : _cause_exc_T_6; // @[Mux.scala 81:58]
  wire [3:0] _cause_exc_T_10 = 3'h4 == io_uop_exc ? 4'h2 : _cause_exc_T_8; // @[Mux.scala 81:58]
  wire [3:0] _cause_exc_T_12 = 3'h7 == io_uop_exc ? 4'h3 : _cause_exc_T_10; // @[Mux.scala 81:58]
  wire [3:0] _cause_exc_T_14 = 3'h5 == io_uop_exc ? _cause_exc_T_4 : _cause_exc_T_12; // @[Mux.scala 81:58]
  wire [3:0] cause_exc = 3'h3 == io_uop_exc ? 4'hc : _cause_exc_T_14; // @[Mux.scala 81:58]
  wire [15:0] cause_exc_onehot = 16'h1 << cause_exc; // @[OneHot.scala 57:35]
  wire [15:0] cause_int_onehot = 16'h1 << int_index; // @[OneHot.scala 57:35]
  wire  trap = is_exc | is_int; // @[CSR.scala 796:26]
  wire [63:0] _GEN_221 = {{48'd0}, cause_exc_onehot}; // @[CSR.scala 801:37]
  wire [63:0] _trap_to_s_T = _GEN_221 & medeleg; // @[CSR.scala 801:37]
  wire [63:0] _GEN_222 = {{48'd0}, cause_int_onehot}; // @[CSR.scala 802:37]
  wire [63:0] _trap_to_s_T_3 = _GEN_222 & mideleg; // @[CSR.scala 802:37]
  wire  _trap_to_s_T_5 = is_int & _trap_to_s_T_3 != 64'h0; // @[CSR.scala 802:15]
  wire  _trap_to_s_T_6 = is_exc & _trap_to_s_T != 64'h0 | _trap_to_s_T_5; // @[CSR.scala 801:58]
  wire  trap_to_s = _is_exc_from_sys_T & _trap_to_s_T_6; // @[CSR.scala 799:19 800:15 797:30]
  wire [63:0] _scause_T = {60'h800000000000000,int_index}; // @[Cat.scala 33:92]
  wire [3:0] _trap_pc_T_4 = is_int & stvec[1:0] == 2'h1 ? int_index : 4'h0; // @[CSR.scala 813:48]
  wire [61:0] _GEN_223 = {{58'd0}, _trap_pc_T_4}; // @[CSR.scala 813:43]
  wire [61:0] _trap_pc_T_6 = stvec[63:2] + _GEN_223; // @[CSR.scala 813:43]
  wire [63:0] _trap_pc_T_7 = {_trap_pc_T_6,2'h0}; // @[Cat.scala 33:92]
  wire [1:0] _GEN_207 = trap_to_s & trap ? prv : {{1'd0}, _GEN_180}; // @[CSR.scala 804:27 810:17]
  wire [1:0] _GEN_208 = trap_to_s & trap ? 2'h1 : _GEN_177; // @[CSR.scala 804:27 811:17]
  wire [63:0] _GEN_209 = trap_to_s & trap ? _trap_pc_T_7 : 64'h0; // @[CSR.scala 804:27 813:17 798:30]
  wire [3:0] _trap_pc_T_12 = is_int & mtvec[1:0] == 2'h1 ? int_index : 4'h0; // @[CSR.scala 824:49]
  wire [61:0] _GEN_224 = {{58'd0}, _trap_pc_T_12}; // @[CSR.scala 824:44]
  wire [61:0] _trap_pc_T_14 = mtvec[63:2] + _GEN_224; // @[CSR.scala 824:44]
  wire [63:0] _trap_pc_T_15 = {_trap_pc_T_14,2'h0}; // @[Cat.scala 33:92]
  wire [63:0] trap_pc = ~trap_to_s & trap ? _trap_pc_T_15 : _GEN_209; // @[CSR.scala 815:28 824:18]
  wire [63:0] _io_jmp_packet_target_T_1 = is_mret ? mepc : sepc; // @[CSR.scala 830:89]
  wire [63:0] _io_jmp_packet_target_T_2 = is_sys | satp_updated ? io_uop_npc : _io_jmp_packet_target_T_1; // @[CSR.scala 830:49]
  wire [1:0] _GEN_225 = reset ? 2'h0 : _GEN_207; // @[CSR.scala 84:{28,28}]
  assign io_rw_rdata = io_rw_addr == 12'hc02 ? instret : _GEN_165; // @[CSR.scala 639:39 640:15]
  assign io_rw_valid = io_rw_addr == 12'hc02 ? mret_legal | prv_is_s & mcounteren[2] | prv_is_u & mcounteren[2] &
    scounteren[2] : _GEN_167; // @[CSR.scala 639:39 641:15]
  assign io_prv = ~trap_to_s & trap ? 2'h3 : _GEN_208; // @[CSR.scala 815:28 822:18]
  assign io_mprv = mstatus_mprv; // @[CSR.scala 184:11]
  assign io_mpp = mstatus_mpp; // @[CSR.scala 185:11]
  assign io_sv39_en = io_rw_addr == 12'h180 ? _GEN_67 : satp[63]; // @[CSR.scala 288:16 291:36]
  assign io_satp_asid = io_rw_addr == 12'h180 ? _GEN_68 : satp[59:44]; // @[CSR.scala 289:16 291:36]
  assign io_satp_ppn = io_rw_addr == 12'h180 ? _GEN_69 : satp[43:0]; // @[CSR.scala 290:16 291:36]
  assign io_sfence_vma = is_sfv & _csr_legal_T_1; // @[CSR.scala 689:27]
  assign io_fence_i = io_uop_sys_op == 3'h5 & io_uop_valid; // @[CSR.scala 687:58]
  assign io_jmp_packet_valid = trap | is_sys | satp_updated | _T_32 | _T_34; // @[CSR.scala 829:85]
  assign io_jmp_packet_target = trap ? trap_pc : _io_jmp_packet_target_T_2; // @[CSR.scala 830:30]
  assign io_is_int = int_attach & int_index != 4'h0; // @[CSR.scala 740:27]
  always @(posedge clock) begin
    if (reset) begin // @[CSR.scala 49:26]
      prv <= 2'h3; // @[CSR.scala 49:26]
    end else if (~trap_to_s & trap) begin // @[CSR.scala 815:28]
      prv <= 2'h3; // @[CSR.scala 822:18]
    end else if (trap_to_s & trap) begin // @[CSR.scala 804:27]
      prv <= 2'h1; // @[CSR.scala 811:17]
    end else if (is_sret & sret_legal) begin // @[CSR.scala 671:31]
      prv <= {{1'd0}, status_spp}; // @[CSR.scala 672:17]
    end else begin
      prv <= _GEN_171;
    end
    if (reset) begin // @[CSR.scala 477:27]
      mcounteren <= 64'h0; // @[CSR.scala 477:27]
    end else if (io_rw_addr == 12'h306) begin // @[CSR.scala 478:42]
      if (wen) begin // @[CSR.scala 480:15]
        if (2'h3 == io_rw_cmd) begin // @[Mux.scala 81:58]
          mcounteren <= _wdata_T_2;
        end else begin
          mcounteren <= _wdata_T_6;
        end
      end
    end
    if (reset) begin // @[CSR.scala 208:27]
      scounteren <= 64'h0; // @[CSR.scala 208:27]
    end else if (io_rw_addr == 12'h106) begin // @[CSR.scala 209:42]
      if (wen) begin // @[CSR.scala 211:15]
        if (2'h3 == io_rw_cmd) begin // @[Mux.scala 81:58]
          scounteren <= _wdata_T_2;
        end else begin
          scounteren <= _wdata_T_6;
        end
      end
    end
    if (reset) begin // @[CSR.scala 117:29]
      mstatus_tvm <= 1'h0; // @[CSR.scala 117:29]
    end else if (io_rw_addr == 12'h300) begin // @[CSR.scala 164:39]
      if (wen) begin // @[CSR.scala 166:15]
        mstatus_tvm <= wdata[20]; // @[CSR.scala 178:20]
      end
    end
    if (reset) begin // @[CSR.scala 630:24]
      instret <= 64'h0; // @[CSR.scala 630:24]
    end else if (io_rw_addr == 12'hb02) begin // @[CSR.scala 632:40]
      if (wen) begin // @[CSR.scala 634:15]
        if (2'h3 == io_rw_cmd) begin // @[Mux.scala 81:58]
          instret <= _wdata_T_2;
        end else begin
          instret <= _wdata_T_6;
        end
      end else begin
        instret <= _instret_T_1; // @[CSR.scala 631:11]
      end
    end else begin
      instret <= _instret_T_1; // @[CSR.scala 631:11]
    end
    if (reset) begin // @[CSR.scala 608:22]
      cycle <= 64'h0; // @[CSR.scala 608:22]
    end else if (io_rw_addr == 12'hb00) begin // @[CSR.scala 610:38]
      if (wen) begin // @[CSR.scala 612:15]
        if (2'h3 == io_rw_cmd) begin // @[Mux.scala 81:58]
          cycle <= _wdata_T_2;
        end else begin
          cycle <= _wdata_T_6;
        end
      end else begin
        cycle <= _cycle_T_1; // @[CSR.scala 609:9]
      end
    end else begin
      cycle <= _cycle_T_1; // @[CSR.scala 609:9]
    end
    if (reset) begin // @[CSR.scala 558:26]
      ip_seip_r <= 1'h0; // @[CSR.scala 558:26]
    end else if (io_rw_addr == 12'h344) begin // @[CSR.scala 585:35]
      if (wen) begin // @[CSR.scala 587:15]
        ip_seip_r <= wdata[9]; // @[CSR.scala 590:17]
      end
    end
    if (reset) begin // @[CSR.scala 556:26]
      ip_stip <= 1'h0; // @[CSR.scala 556:26]
    end else if (io_rw_addr == 12'h344) begin // @[CSR.scala 585:35]
      if (wen) begin // @[CSR.scala 587:15]
        ip_stip <= wdata[5]; // @[CSR.scala 589:17]
      end
    end
    if (reset) begin // @[CSR.scala 554:26]
      ip_ssip <= 1'h0; // @[CSR.scala 554:26]
    end else if (io_rw_addr == 12'h144) begin // @[CSR.scala 594:35]
      if (wen) begin // @[CSR.scala 596:15]
        ip_ssip <= wdata[1]; // @[CSR.scala 597:15]
      end else begin
        ip_ssip <= _GEN_150;
      end
    end else begin
      ip_ssip <= _GEN_150;
    end
    if (reset) begin // @[CSR.scala 537:22]
      mtval <= 64'h0; // @[CSR.scala 537:22]
    end else if (~trap_to_s & trap) begin // @[CSR.scala 815:28]
      if (io_uop_exc == 3'h3) begin // @[CSR.scala 792:39]
        mtval <= io_uop_pc; // @[CSR.scala 793:10]
      end else if (is_exc_from_lsu) begin // @[CSR.scala 789:25]
        mtval <= io_lsu_addr; // @[CSR.scala 790:10]
      end else begin
        mtval <= 64'h0; // @[CSR.scala 788:25]
      end
    end else if (io_rw_addr == 12'h343) begin // @[CSR.scala 538:37]
      if (wen) begin // @[CSR.scala 540:15]
        mtval <= wdata; // @[CSR.scala 541:13]
      end
    end
    if (reset) begin // @[CSR.scala 522:23]
      mcause <= 64'h0; // @[CSR.scala 522:23]
    end else if (~trap_to_s & trap) begin // @[CSR.scala 815:28]
      if (is_exc) begin // @[CSR.scala 806:23]
        mcause <= {{60'd0}, cause_exc};
      end else begin
        mcause <= _scause_T;
      end
    end else if (io_rw_addr == 12'h342) begin // @[CSR.scala 523:38]
      if (wen) begin // @[CSR.scala 525:15]
        mcause <= wdata; // @[CSR.scala 526:14]
      end
    end
    if (reset) begin // @[CSR.scala 507:21]
      mepc <= 64'h0; // @[CSR.scala 507:21]
    end else if (~trap_to_s & trap) begin // @[CSR.scala 815:28]
      mepc <= io_uop_pc; // @[CSR.scala 818:18]
    end else if (io_rw_addr == 12'h341) begin // @[CSR.scala 508:36]
      if (wen) begin // @[CSR.scala 510:15]
        mepc <= wdata; // @[CSR.scala 511:12]
      end
    end
    if (reset) begin // @[CSR.scala 492:25]
      mscratch <= 64'h0; // @[CSR.scala 492:25]
    end else if (io_rw_addr == 12'h340) begin // @[CSR.scala 493:40]
      if (wen) begin // @[CSR.scala 495:15]
        if (2'h3 == io_rw_cmd) begin // @[Mux.scala 81:58]
          mscratch <= _wdata_T_2;
        end else begin
          mscratch <= _wdata_T_6;
        end
      end
    end
    if (reset) begin // @[CSR.scala 462:22]
      mtvec <= 64'h0; // @[CSR.scala 462:22]
    end else if (io_rw_addr == 12'h305) begin // @[CSR.scala 463:37]
      if (wen) begin // @[CSR.scala 465:15]
        if (2'h3 == io_rw_cmd) begin // @[Mux.scala 81:58]
          mtvec <= _wdata_T_2;
        end else begin
          mtvec <= _wdata_T_6;
        end
      end
    end
    if (reset) begin // @[CSR.scala 408:24]
      ie_seie <= 1'h0; // @[CSR.scala 408:24]
    end else if (io_rw_addr == 12'h104) begin // @[CSR.scala 446:35]
      if (wen) begin // @[CSR.scala 448:15]
        ie_seie <= wdata[9]; // @[CSR.scala 451:15]
      end else begin
        ie_seie <= _GEN_111;
      end
    end else begin
      ie_seie <= _GEN_111;
    end
    if (reset) begin // @[CSR.scala 406:24]
      ie_stie <= 1'h0; // @[CSR.scala 406:24]
    end else if (io_rw_addr == 12'h104) begin // @[CSR.scala 446:35]
      if (wen) begin // @[CSR.scala 448:15]
        ie_stie <= wdata[5]; // @[CSR.scala 450:15]
      end else begin
        ie_stie <= _GEN_109;
      end
    end else begin
      ie_stie <= _GEN_109;
    end
    if (reset) begin // @[CSR.scala 404:24]
      ie_ssie <= 1'h0; // @[CSR.scala 404:24]
    end else if (io_rw_addr == 12'h104) begin // @[CSR.scala 446:35]
      if (wen) begin // @[CSR.scala 448:15]
        ie_ssie <= wdata[1]; // @[CSR.scala 449:15]
      end else begin
        ie_ssie <= _GEN_107;
      end
    end else begin
      ie_ssie <= _GEN_107;
    end
    if (reset) begin // @[CSR.scala 409:24]
      ie_meie <= 1'h0; // @[CSR.scala 409:24]
    end else if (io_rw_addr == 12'h304) begin // @[CSR.scala 434:35]
      if (wen) begin // @[CSR.scala 436:15]
        ie_meie <= wdata[11]; // @[CSR.scala 442:15]
      end
    end
    if (reset) begin // @[CSR.scala 407:24]
      ie_mtie <= 1'h0; // @[CSR.scala 407:24]
    end else if (io_rw_addr == 12'h304) begin // @[CSR.scala 434:35]
      if (wen) begin // @[CSR.scala 436:15]
        ie_mtie <= wdata[7]; // @[CSR.scala 440:15]
      end
    end
    if (reset) begin // @[CSR.scala 405:24]
      ie_msie <= 1'h0; // @[CSR.scala 405:24]
    end else if (io_rw_addr == 12'h304) begin // @[CSR.scala 434:35]
      if (wen) begin // @[CSR.scala 436:15]
        ie_msie <= wdata[3]; // @[CSR.scala 438:15]
      end
    end
    if (reset) begin // @[CSR.scala 387:24]
      mideleg <= 64'h0; // @[CSR.scala 387:24]
    end else if (io_rw_addr == 12'h303) begin // @[CSR.scala 388:39]
      if (wen) begin // @[CSR.scala 390:15]
        mideleg <= _mideleg_T; // @[CSR.scala 391:15]
      end
    end
    if (reset) begin // @[CSR.scala 372:24]
      medeleg <= 64'h0; // @[CSR.scala 372:24]
    end else if (io_rw_addr == 12'h302) begin // @[CSR.scala 373:39]
      if (wen) begin // @[CSR.scala 375:15]
        medeleg <= _medeleg_T; // @[CSR.scala 376:15]
      end
    end
    if (reset) begin // @[CSR.scala 342:33]
      mhartid <= 64'h0; // @[CSR.scala 342:33]
    end else if (io_rw_addr == 12'hf14) begin // @[CSR.scala 344:39]
      if (wen & mhartid_writable) begin // @[CSR.scala 346:35]
        if (2'h3 == io_rw_cmd) begin // @[Mux.scala 81:58]
          mhartid <= _wdata_T_2;
        end else begin
          mhartid <= _wdata_T_6;
        end
      end
    end
    if (reset) begin // @[CSR.scala 283:29]
      satp <= 64'h0; // @[CSR.scala 283:29]
    end else if (io_rw_addr == 12'h180) begin // @[CSR.scala 291:36]
      if (wen & satp_wen) begin // @[CSR.scala 293:27]
        if (2'h3 == io_rw_cmd) begin // @[Mux.scala 81:58]
          satp <= _wdata_T_2;
        end else begin
          satp <= _wdata_T_6;
        end
      end
    end
    if (reset) begin // @[CSR.scala 268:22]
      stval <= 64'h0; // @[CSR.scala 268:22]
    end else if (trap_to_s & trap) begin // @[CSR.scala 804:27]
      if (io_uop_exc == 3'h3) begin // @[CSR.scala 792:39]
        stval <= io_uop_pc; // @[CSR.scala 793:10]
      end else if (is_exc_from_lsu) begin // @[CSR.scala 789:25]
        stval <= io_lsu_addr; // @[CSR.scala 790:10]
      end else begin
        stval <= 64'h0; // @[CSR.scala 788:25]
      end
    end else if (io_rw_addr == 12'h143) begin // @[CSR.scala 269:37]
      if (wen) begin // @[CSR.scala 271:15]
        stval <= wdata; // @[CSR.scala 272:13]
      end
    end
    if (reset) begin // @[CSR.scala 253:23]
      scause <= 64'h0; // @[CSR.scala 253:23]
    end else if (trap_to_s & trap) begin // @[CSR.scala 804:27]
      if (is_exc) begin // @[CSR.scala 806:23]
        scause <= {{60'd0}, cause_exc};
      end else begin
        scause <= _scause_T;
      end
    end else if (io_rw_addr == 12'h142) begin // @[CSR.scala 254:38]
      if (wen) begin // @[CSR.scala 256:15]
        scause <= wdata; // @[CSR.scala 257:14]
      end
    end
    if (reset) begin // @[CSR.scala 238:21]
      sepc <= 64'h0; // @[CSR.scala 238:21]
    end else if (trap_to_s & trap) begin // @[CSR.scala 804:27]
      sepc <= io_uop_pc; // @[CSR.scala 807:17]
    end else if (io_rw_addr == 12'h141) begin // @[CSR.scala 239:36]
      if (wen) begin // @[CSR.scala 241:15]
        sepc <= wdata; // @[CSR.scala 242:12]
      end
    end
    if (reset) begin // @[CSR.scala 223:25]
      sscratch <= 64'h0; // @[CSR.scala 223:25]
    end else if (io_rw_addr == 12'h140) begin // @[CSR.scala 224:40]
      if (wen) begin // @[CSR.scala 226:15]
        if (2'h3 == io_rw_cmd) begin // @[Mux.scala 81:58]
          sscratch <= _wdata_T_2;
        end else begin
          sscratch <= _wdata_T_6;
        end
      end
    end
    if (reset) begin // @[CSR.scala 193:22]
      stvec <= 64'h0; // @[CSR.scala 193:22]
    end else if (io_rw_addr == 12'h105) begin // @[CSR.scala 194:37]
      if (wen) begin // @[CSR.scala 196:15]
        if (2'h3 == io_rw_cmd) begin // @[Mux.scala 81:58]
          stvec <= _wdata_T_2;
        end else begin
          stvec <= _wdata_T_6;
        end
      end
    end
    if (reset) begin // @[CSR.scala 86:28]
      status_fs <= 2'h0; // @[CSR.scala 86:28]
    end else if (io_rw_addr == 12'h300) begin // @[CSR.scala 164:39]
      if (wen) begin // @[CSR.scala 166:15]
        status_fs <= wdata[14:13]; // @[CSR.scala 170:19]
      end else begin
        status_fs <= _GEN_10;
      end
    end else begin
      status_fs <= _GEN_10;
    end
    if (reset) begin // @[CSR.scala 119:29]
      mstatus_tsr <= 1'h0; // @[CSR.scala 119:29]
    end else if (io_rw_addr == 12'h300) begin // @[CSR.scala 164:39]
      if (wen) begin // @[CSR.scala 166:15]
        mstatus_tsr <= wdata[22]; // @[CSR.scala 180:20]
      end
    end
    if (reset) begin // @[CSR.scala 118:29]
      mstatus_tw <= 1'h0; // @[CSR.scala 118:29]
    end else if (io_rw_addr == 12'h300) begin // @[CSR.scala 164:39]
      if (wen) begin // @[CSR.scala 166:15]
        mstatus_tw <= wdata[21]; // @[CSR.scala 179:20]
      end
    end
    if (reset) begin // @[CSR.scala 89:28]
      status_mxr <= 1'h0; // @[CSR.scala 89:28]
    end else if (io_rw_addr == 12'h300) begin // @[CSR.scala 164:39]
      if (wen) begin // @[CSR.scala 166:15]
        status_mxr <= wdata[19]; // @[CSR.scala 173:20]
      end else begin
        status_mxr <= _GEN_12;
      end
    end else begin
      status_mxr <= _GEN_12;
    end
    if (reset) begin // @[CSR.scala 88:28]
      status_sum <= 1'h0; // @[CSR.scala 88:28]
    end else if (io_rw_addr == 12'h300) begin // @[CSR.scala 164:39]
      if (wen) begin // @[CSR.scala 166:15]
        status_sum <= wdata[18]; // @[CSR.scala 172:20]
      end else begin
        status_sum <= _GEN_11;
      end
    end else begin
      status_sum <= _GEN_11;
    end
    if (reset) begin // @[CSR.scala 116:29]
      mstatus_mprv <= 1'h0; // @[CSR.scala 116:29]
    end else if (is_sret & sret_legal) begin // @[CSR.scala 671:31]
      if (_GEN_219 != 2'h3) begin // @[CSR.scala 677:34]
        mstatus_mprv <= 1'h0; // @[CSR.scala 678:20]
      end else begin
        mstatus_mprv <= _GEN_175;
      end
    end else begin
      mstatus_mprv <= _GEN_175;
    end
    if (reset) begin // @[CSR.scala 115:29]
      mstatus_mpp <= 2'h0; // @[CSR.scala 115:29]
    end else if (~trap_to_s & trap) begin // @[CSR.scala 815:28]
      mstatus_mpp <= prv; // @[CSR.scala 821:18]
    end else if (is_mret & mret_legal) begin // @[CSR.scala 658:31]
      mstatus_mpp <= 2'h0; // @[CSR.scala 663:18]
    end else if (io_rw_addr == 12'h300) begin // @[CSR.scala 164:39]
      mstatus_mpp <= _GEN_22;
    end
    status_spp <= _GEN_225[0]; // @[CSR.scala 84:{28,28}]
    if (reset) begin // @[CSR.scala 114:29]
      mstatus_mpie <= 1'h0; // @[CSR.scala 114:29]
    end else if (~trap_to_s & trap) begin // @[CSR.scala 815:28]
      mstatus_mpie <= mstatus_mie; // @[CSR.scala 819:18]
    end else begin
      mstatus_mpie <= _GEN_173;
    end
    if (reset) begin // @[CSR.scala 82:28]
      status_spie <= 1'h0; // @[CSR.scala 82:28]
    end else if (trap_to_s & trap) begin // @[CSR.scala 804:27]
      status_spie <= status_sie; // @[CSR.scala 808:17]
    end else begin
      status_spie <= _GEN_179;
    end
    if (reset) begin // @[CSR.scala 113:29]
      mstatus_mie <= 1'h0; // @[CSR.scala 113:29]
    end else if (~trap_to_s & trap) begin // @[CSR.scala 815:28]
      mstatus_mie <= 1'h0; // @[CSR.scala 820:18]
    end else if (is_mret & mret_legal) begin // @[CSR.scala 658:31]
      mstatus_mie <= mstatus_mpie; // @[CSR.scala 661:18]
    end else if (io_rw_addr == 12'h300) begin // @[CSR.scala 164:39]
      mstatus_mie <= _GEN_20;
    end
    if (reset) begin // @[CSR.scala 81:28]
      status_sie <= 1'h0; // @[CSR.scala 81:28]
    end else if (trap_to_s & trap) begin // @[CSR.scala 804:27]
      status_sie <= 1'h0; // @[CSR.scala 809:17]
    end else if (is_sret & sret_legal) begin // @[CSR.scala 671:31]
      status_sie <= status_spie; // @[CSR.scala 674:17]
    end else if (io_rw_addr == 12'h300) begin // @[CSR.scala 164:39]
      status_sie <= _GEN_14;
    end else begin
      status_sie <= _GEN_7;
    end
    mhartid_writable <= reset | _GEN_88; // @[CSR.scala 343:{33,33}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  prv = _RAND_0[1:0];
  _RAND_1 = {2{`RANDOM}};
  mcounteren = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  scounteren = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  mstatus_tvm = _RAND_3[0:0];
  _RAND_4 = {2{`RANDOM}};
  instret = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  cycle = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  ip_seip_r = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  ip_stip = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  ip_ssip = _RAND_8[0:0];
  _RAND_9 = {2{`RANDOM}};
  mtval = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  mcause = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  mepc = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  mscratch = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  mtvec = _RAND_13[63:0];
  _RAND_14 = {1{`RANDOM}};
  ie_seie = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  ie_stie = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  ie_ssie = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  ie_meie = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  ie_mtie = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  ie_msie = _RAND_19[0:0];
  _RAND_20 = {2{`RANDOM}};
  mideleg = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  medeleg = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  mhartid = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  satp = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  stval = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  scause = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  sepc = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  sscratch = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  stvec = _RAND_28[63:0];
  _RAND_29 = {1{`RANDOM}};
  status_fs = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  mstatus_tsr = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  mstatus_tw = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  status_mxr = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  status_sum = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  mstatus_mprv = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  mstatus_mpp = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  status_spp = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  mstatus_mpie = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  status_spie = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  mstatus_mie = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  status_sie = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  mhartid_writable = _RAND_41[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CachePortProxy_1(
  input         clock,
  input         reset,
  input  [1:0]  io_prv,
  input         io_sv39_en,
  input  [15:0] io_satp_asid,
  input  [43:0] io_satp_ppn,
  input         io_sfence_vma,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [38:0] io_in_req_bits_addr,
  input  [63:0] io_in_req_bits_wdata,
  input  [7:0]  io_in_req_bits_wmask,
  input         io_in_req_bits_wen,
  input  [1:0]  io_in_req_bits_len,
  input         io_in_req_bits_lrsc,
  input  [4:0]  io_in_req_bits_amo,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [63:0] io_in_resp_bits_rdata,
  output        io_in_resp_bits_page_fault,
  output        io_in_resp_bits_access_fault,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [38:0] io_out_req_bits_addr,
  output [63:0] io_out_req_bits_wdata,
  output [7:0]  io_out_req_bits_wmask,
  output        io_out_req_bits_wen,
  output [1:0]  io_out_req_bits_len,
  output        io_out_req_bits_lrsc,
  output [4:0]  io_out_req_bits_amo,
  output        io_out_resp_ready,
  input         io_out_resp_valid,
  input  [63:0] io_out_resp_bits_rdata,
  input         io_ptw_req_ready,
  output        io_ptw_req_valid,
  output [38:0] io_ptw_req_bits_addr,
  output        io_ptw_resp_ready,
  input         io_ptw_resp_valid,
  input  [63:0] io_ptw_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
`endif // RANDOMIZE_REG_INIT
  wire  tlb_clock; // @[CachePortProxy.scala 28:19]
  wire  tlb_reset; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_sfence_vma; // @[CachePortProxy.scala 28:19]
  wire [8:0] tlb_io_vaddr_vpn2; // @[CachePortProxy.scala 28:19]
  wire [8:0] tlb_io_vaddr_vpn1; // @[CachePortProxy.scala 28:19]
  wire [8:0] tlb_io_vaddr_vpn0; // @[CachePortProxy.scala 28:19]
  wire [1:0] tlb_io_rpte_ppn2; // @[CachePortProxy.scala 28:19]
  wire [8:0] tlb_io_rpte_ppn1; // @[CachePortProxy.scala 28:19]
  wire [8:0] tlb_io_rpte_ppn0; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_rpte_flag_d; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_rpte_flag_a; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_rpte_flag_u; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_rpte_flag_x; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_rpte_flag_w; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_rpte_flag_r; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_rpte_flag_v; // @[CachePortProxy.scala 28:19]
  wire [1:0] tlb_io_rlevel; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_hit; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_wen; // @[CachePortProxy.scala 28:19]
  wire [8:0] tlb_io_wvaddr_vpn2; // @[CachePortProxy.scala 28:19]
  wire [8:0] tlb_io_wvaddr_vpn1; // @[CachePortProxy.scala 28:19]
  wire [8:0] tlb_io_wvaddr_vpn0; // @[CachePortProxy.scala 28:19]
  wire [1:0] tlb_io_wpte_ppn2; // @[CachePortProxy.scala 28:19]
  wire [8:0] tlb_io_wpte_ppn1; // @[CachePortProxy.scala 28:19]
  wire [8:0] tlb_io_wpte_ppn0; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_wpte_flag_d; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_wpte_flag_a; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_wpte_flag_g; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_wpte_flag_u; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_wpte_flag_x; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_wpte_flag_w; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_wpte_flag_r; // @[CachePortProxy.scala 28:19]
  wire  tlb_io_wpte_flag_v; // @[CachePortProxy.scala 28:19]
  wire [1:0] tlb_io_wlevel; // @[CachePortProxy.scala 28:19]
  wire [15:0] tlb_io_satp_asid; // @[CachePortProxy.scala 28:19]
  reg [2:0] state; // @[CachePortProxy.scala 21:93]
  wire  _in_req_bits_T = state == 3'h0; // @[CachePortProxy.scala 24:54]
  reg [38:0] in_req_bits_r_addr; // @[Reg.scala 35:20]
  reg [63:0] in_req_bits_r_wdata; // @[Reg.scala 35:20]
  reg [7:0] in_req_bits_r_wmask; // @[Reg.scala 35:20]
  reg  in_req_bits_r_wen; // @[Reg.scala 35:20]
  reg [1:0] in_req_bits_r_len; // @[Reg.scala 35:20]
  reg  in_req_bits_r_lrsc; // @[Reg.scala 35:20]
  reg [4:0] in_req_bits_r_amo; // @[Reg.scala 35:20]
  wire [38:0] _GEN_0 = _in_req_bits_T ? io_in_req_bits_addr : in_req_bits_r_addr; // @[Reg.scala 36:18 35:20 36:22]
  wire  _GEN_3 = _in_req_bits_T ? io_in_req_bits_wen : in_req_bits_r_wen; // @[Reg.scala 36:18 35:20 36:22]
  wire [11:0] in_vaddr_offset = _GEN_0[11:0]; // @[CachePortProxy.scala 25:46]
  wire [8:0] in_vaddr_vpn0 = _GEN_0[20:12]; // @[CachePortProxy.scala 25:46]
  wire [8:0] in_vaddr_vpn1 = _GEN_0[29:21]; // @[CachePortProxy.scala 25:46]
  wire [8:0] in_vaddr_vpn2 = _GEN_0[38:30]; // @[CachePortProxy.scala 25:46]
  wire  _atp_en_T_1 = io_prv != 2'h3 & io_sv39_en; // @[CachePortProxy.scala 38:48]
  reg  atp_en_r; // @[Reg.scala 35:20]
  wire  _GEN_7 = _in_req_bits_T ? _atp_en_T_1 : atp_en_r; // @[Reg.scala 36:18 35:20 36:22]
  wire  in_addr_invalid = io_in_req_bits_addr < 39'h10000; // @[CachePortProxy.scala 42:34]
  wire  _access_fault_T_3 = ~_GEN_7; // @[CachePortProxy.scala 43:73]
  wire  access_fault = ~io_in_req_bits_addr[31] & (io_prv == 2'h3 | ~_GEN_7) & in_addr_invalid; // @[CachePortProxy.scala 43:82]
  reg [1:0] ptw_level; // @[CachePortProxy.scala 46:29]
  wire  ptw_pte_flag_v = io_ptw_resp_bits_rdata[0]; // @[CachePortProxy.scala 47:53]
  wire  ptw_pte_flag_r = io_ptw_resp_bits_rdata[1]; // @[CachePortProxy.scala 47:53]
  wire  ptw_pte_flag_w = io_ptw_resp_bits_rdata[2]; // @[CachePortProxy.scala 47:53]
  wire  ptw_pte_flag_x = io_ptw_resp_bits_rdata[3]; // @[CachePortProxy.scala 47:53]
  wire  ptw_pte_flag_u = io_ptw_resp_bits_rdata[4]; // @[CachePortProxy.scala 47:53]
  wire  ptw_pte_flag_g = io_ptw_resp_bits_rdata[5]; // @[CachePortProxy.scala 47:53]
  wire  ptw_pte_flag_a = io_ptw_resp_bits_rdata[6]; // @[CachePortProxy.scala 47:53]
  wire  ptw_pte_flag_d = io_ptw_resp_bits_rdata[7]; // @[CachePortProxy.scala 47:53]
  wire [8:0] ptw_pte_ppn0 = io_ptw_resp_bits_rdata[18:10]; // @[CachePortProxy.scala 47:53]
  wire [8:0] ptw_pte_ppn1 = io_ptw_resp_bits_rdata[27:19]; // @[CachePortProxy.scala 47:53]
  wire [1:0] ptw_pte_ppn2 = io_ptw_resp_bits_rdata[29:28]; // @[CachePortProxy.scala 47:53]
  wire  _ptw_pte_reg_T = io_ptw_resp_ready & io_ptw_resp_valid; // @[Decoupled.scala 51:35]
  reg [1:0] ptw_pte_reg_ppn2; // @[Reg.scala 35:20]
  reg [8:0] ptw_pte_reg_ppn1; // @[Reg.scala 35:20]
  reg [8:0] ptw_pte_reg_ppn0; // @[Reg.scala 35:20]
  reg  ptw_pte_reg_flag_d; // @[Reg.scala 35:20]
  reg  ptw_pte_reg_flag_a; // @[Reg.scala 35:20]
  reg  ptw_pte_reg_flag_g; // @[Reg.scala 35:20]
  reg  ptw_pte_reg_flag_u; // @[Reg.scala 35:20]
  reg  ptw_pte_reg_flag_x; // @[Reg.scala 35:20]
  reg  ptw_pte_reg_flag_w; // @[Reg.scala 35:20]
  reg  ptw_pte_reg_flag_r; // @[Reg.scala 35:20]
  reg  ptw_pte_reg_flag_v; // @[Reg.scala 35:20]
  wire  _ptw_complete_T_4 = ptw_pte_flag_r | ptw_pte_flag_x; // @[CachePortProxy.scala 7:37]
  wire  ptw_complete = ~ptw_pte_flag_v | ~ptw_pte_flag_r & ptw_pte_flag_w | _ptw_complete_T_4 | ptw_level == 2'h0; // @[CachePortProxy.scala 49:96]
  wire  _T_1 = io_in_req_ready & io_in_req_valid; // @[Decoupled.scala 51:35]
  wire  _T_2 = ~tlb_io_hit; // @[CachePortProxy.scala 55:24]
  wire [2:0] _GEN_20 = _GEN_7 & ~tlb_io_hit ? 3'h1 : state; // @[CachePortProxy.scala 55:37 56:17 21:93]
  wire [2:0] _GEN_21 = _T_1 ? _GEN_20 : state; // @[CachePortProxy.scala 54:28 21:93]
  wire  _T_7 = io_ptw_req_ready & io_ptw_req_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _ptw_level_T_1 = ptw_level - 2'h1; // @[CachePortProxy.scala 77:34]
  wire [2:0] _GEN_25 = ptw_complete ? 3'h3 : 3'h1; // @[CachePortProxy.scala 73:28 74:17 76:21]
  wire [1:0] _GEN_26 = ptw_complete ? ptw_level : _ptw_level_T_1; // @[CachePortProxy.scala 73:28 46:29 77:21]
  wire [2:0] _GEN_27 = _ptw_pte_reg_T ? _GEN_25 : state; // @[CachePortProxy.scala 72:30 21:93]
  wire [1:0] _GEN_28 = _ptw_pte_reg_T ? _GEN_26 : ptw_level; // @[CachePortProxy.scala 46:29 72:30]
  wire  _T_11 = io_out_req_ready & io_out_req_valid; // @[Decoupled.scala 51:35]
  wire  pte_flag_v = _in_req_bits_T ? tlb_io_rpte_flag_v : ptw_pte_reg_flag_v; // @[CachePortProxy.scala 117:18]
  wire  pte_flag_r = _in_req_bits_T ? tlb_io_rpte_flag_r : ptw_pte_reg_flag_r; // @[CachePortProxy.scala 117:18]
  wire  _T_16 = ~pte_flag_r; // @[CachePortProxy.scala 132:24]
  wire  pte_flag_w = _in_req_bits_T ? tlb_io_rpte_flag_w : ptw_pte_reg_flag_w; // @[CachePortProxy.scala 117:18]
  wire  pf1 = ~pte_flag_v | ~pte_flag_r & pte_flag_w; // @[CachePortProxy.scala 132:20]
  wire  pte_flag_x = _in_req_bits_T ? tlb_io_rpte_flag_x : ptw_pte_reg_flag_x; // @[CachePortProxy.scala 117:18]
  wire  _T_19 = pte_flag_r | pte_flag_x; // @[CachePortProxy.scala 7:37]
  wire  pte_flag_a = _in_req_bits_T ? tlb_io_rpte_flag_a : ptw_pte_reg_flag_a; // @[CachePortProxy.scala 117:18]
  wire  _T_20 = ~pte_flag_a; // @[CachePortProxy.scala 136:10]
  wire  pf2 = _T_19 & _T_20; // @[CachePortProxy.scala 135:21 128:24]
  reg [1:0] prv_r; // @[Reg.scala 35:20]
  wire [1:0] prv = _in_req_bits_T ? io_prv : prv_r; // @[Utils.scala 50:8]
  wire  pte_flag_u = _in_req_bits_T ? tlb_io_rpte_flag_u : ptw_pte_reg_flag_u; // @[CachePortProxy.scala 117:18]
  wire  _T_23 = prv == 2'h0 & ~pte_flag_u; // @[CachePortProxy.scala 139:26]
  wire  pf3 = _T_19 & _T_23; // @[CachePortProxy.scala 135:21 129:24]
  wire  pte_flag_d = _in_req_bits_T ? tlb_io_rpte_flag_d : ptw_pte_reg_flag_d; // @[CachePortProxy.scala 117:18]
  wire  _T_29 = _GEN_3 & (~pte_flag_w | _T_16 | ~pte_flag_d); // @[CachePortProxy.scala 148:28]
  wire  pf4 = _T_19 & _T_29; // @[CachePortProxy.scala 135:21 130:24]
  wire  _T_30 = state == 3'h3; // @[CachePortProxy.scala 152:16]
  wire [8:0] pte_ppn1 = _in_req_bits_T ? tlb_io_rpte_ppn1 : ptw_pte_reg_ppn1; // @[CachePortProxy.scala 117:18]
  wire [8:0] pte_ppn0 = _in_req_bits_T ? tlb_io_rpte_ppn0 : ptw_pte_reg_ppn0; // @[CachePortProxy.scala 117:18]
  wire [17:0] _T_32 = {pte_ppn1,pte_ppn0}; // @[Cat.scala 33:92]
  wire  _T_38 = ptw_level == 2'h2 & _T_32 != 18'h0 | ptw_level == 2'h1 & pte_ppn0 != 9'h0; // @[CachePortProxy.scala 153:67]
  wire  _GEN_45 = state == 3'h3 & _T_38; // @[CachePortProxy.scala 131:24 152:36]
  wire  pf5 = _T_19 & _GEN_45; // @[CachePortProxy.scala 135:21 131:24]
  wire  page_fault = pf1 | pf2 | pf3 | pf4 | pf5; // @[CachePortProxy.scala 158:42]
  wire [2:0] _GEN_29 = _T_11 | page_fault ? 3'h0 : state; // @[CachePortProxy.scala 82:43 83:15 21:93]
  wire  _T_14 = io_in_resp_ready & io_in_resp_valid; // @[Decoupled.scala 51:35]
  wire [2:0] _GEN_30 = _T_14 ? 3'h0 : state; // @[CachePortProxy.scala 87:29 88:15 21:93]
  wire [2:0] _GEN_31 = 3'h4 == state ? _GEN_30 : state; // @[CachePortProxy.scala 52:17 21:93]
  wire [2:0] _GEN_32 = 3'h3 == state ? _GEN_29 : _GEN_31; // @[CachePortProxy.scala 52:17]
  wire [55:0] _l2_addr_T = {io_satp_ppn,in_vaddr_vpn2,3'h0}; // @[Cat.scala 33:92]
  wire [31:0] l1_addr = {ptw_pte_reg_ppn2,ptw_pte_reg_ppn1,ptw_pte_reg_ppn0,in_vaddr_vpn1,3'h0}; // @[Cat.scala 33:92]
  wire [31:0] l0_addr = {ptw_pte_reg_ppn2,ptw_pte_reg_ppn1,ptw_pte_reg_ppn0,in_vaddr_vpn0,3'h0}; // @[Cat.scala 33:92]
  wire [31:0] l2_addr = _l2_addr_T[31:0]; // @[CachePortProxy.scala 94:21 98:11]
  wire [31:0] _io_ptw_req_bits_addr_T_1 = 2'h2 == ptw_level ? l2_addr : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] _io_ptw_req_bits_addr_T_3 = 2'h1 == ptw_level ? l1_addr : _io_ptw_req_bits_addr_T_1; // @[Mux.scala 81:58]
  wire [31:0] _io_ptw_req_bits_addr_T_5 = 2'h0 == ptw_level ? l0_addr : _io_ptw_req_bits_addr_T_3; // @[Mux.scala 81:58]
  wire [1:0] pte_ppn2 = _in_req_bits_T ? tlb_io_rpte_ppn2 : ptw_pte_reg_ppn2; // @[CachePortProxy.scala 117:18]
  wire [1:0] level = _in_req_bits_T ? tlb_io_rlevel : ptw_level; // @[CachePortProxy.scala 118:18]
  wire  _tlb_io_wen_T_1 = ~page_fault; // @[CachePortProxy.scala 121:50]
  wire  _tlb_io_wen_T_2 = _T_30 & ~page_fault; // @[CachePortProxy.scala 121:47]
  wire [8:0] paddr_ppn0 = level > 2'h0 ? in_vaddr_vpn0 : pte_ppn0; // @[CachePortProxy.scala 163:22]
  wire [8:0] paddr_ppn1 = level > 2'h1 ? in_vaddr_vpn1 : pte_ppn1; // @[CachePortProxy.scala 164:22]
  wire [31:0] _io_out_req_bits_addr_T = {pte_ppn2,paddr_ppn1,paddr_ppn0,in_vaddr_offset}; // @[CachePortProxy.scala 173:43]
  wire [38:0] _io_out_req_bits_addr_WIRE = {{7'd0}, _io_out_req_bits_addr_T}; // @[CachePortProxy.scala 173:{43,43}]
  wire  _page_fault_reg_T_7 = page_fault & _GEN_7 & (_in_req_bits_T & tlb_io_hit & _T_1 | _T_30); // @[CachePortProxy.scala 178:26]
  reg  page_fault_reg; // @[Utils.scala 36:20]
  wire  _GEN_51 = _page_fault_reg_T_7 | page_fault_reg; // @[Utils.scala 41:19 36:20 41:23]
  TLB tlb ( // @[CachePortProxy.scala 28:19]
    .clock(tlb_clock),
    .reset(tlb_reset),
    .io_sfence_vma(tlb_io_sfence_vma),
    .io_vaddr_vpn2(tlb_io_vaddr_vpn2),
    .io_vaddr_vpn1(tlb_io_vaddr_vpn1),
    .io_vaddr_vpn0(tlb_io_vaddr_vpn0),
    .io_rpte_ppn2(tlb_io_rpte_ppn2),
    .io_rpte_ppn1(tlb_io_rpte_ppn1),
    .io_rpte_ppn0(tlb_io_rpte_ppn0),
    .io_rpte_flag_d(tlb_io_rpte_flag_d),
    .io_rpte_flag_a(tlb_io_rpte_flag_a),
    .io_rpte_flag_u(tlb_io_rpte_flag_u),
    .io_rpte_flag_x(tlb_io_rpte_flag_x),
    .io_rpte_flag_w(tlb_io_rpte_flag_w),
    .io_rpte_flag_r(tlb_io_rpte_flag_r),
    .io_rpte_flag_v(tlb_io_rpte_flag_v),
    .io_rlevel(tlb_io_rlevel),
    .io_hit(tlb_io_hit),
    .io_wen(tlb_io_wen),
    .io_wvaddr_vpn2(tlb_io_wvaddr_vpn2),
    .io_wvaddr_vpn1(tlb_io_wvaddr_vpn1),
    .io_wvaddr_vpn0(tlb_io_wvaddr_vpn0),
    .io_wpte_ppn2(tlb_io_wpte_ppn2),
    .io_wpte_ppn1(tlb_io_wpte_ppn1),
    .io_wpte_ppn0(tlb_io_wpte_ppn0),
    .io_wpte_flag_d(tlb_io_wpte_flag_d),
    .io_wpte_flag_a(tlb_io_wpte_flag_a),
    .io_wpte_flag_g(tlb_io_wpte_flag_g),
    .io_wpte_flag_u(tlb_io_wpte_flag_u),
    .io_wpte_flag_x(tlb_io_wpte_flag_x),
    .io_wpte_flag_w(tlb_io_wpte_flag_w),
    .io_wpte_flag_r(tlb_io_wpte_flag_r),
    .io_wpte_flag_v(tlb_io_wpte_flag_v),
    .io_wlevel(tlb_io_wlevel),
    .io_satp_asid(tlb_io_satp_asid)
  );
  assign io_in_req_ready = _in_req_bits_T & (io_out_req_ready | access_fault | _GEN_7 & (_T_2 | page_fault)); // @[CachePortProxy.scala 168:41]
  assign io_in_resp_valid = io_out_resp_valid | io_in_resp_bits_page_fault | io_in_resp_bits_access_fault; // @[CachePortProxy.scala 185:83]
  assign io_in_resp_bits_rdata = io_out_resp_bits_rdata; // @[CachePortProxy.scala 181:32]
  assign io_in_resp_bits_page_fault = page_fault_reg; // @[CachePortProxy.scala 182:32]
  assign io_in_resp_bits_access_fault = state == 3'h4; // @[CachePortProxy.scala 183:42]
  assign io_out_req_valid = _in_req_bits_T & (tlb_io_hit & _tlb_io_wen_T_1 | _access_fault_T_3 & ~access_fault) &
    io_in_req_valid | _tlb_io_wen_T_2; // @[CachePortProxy.scala 169:126]
  assign io_out_req_bits_addr = _GEN_7 ? _io_out_req_bits_addr_WIRE : _GEN_0; // @[CachePortProxy.scala 172:16 171:19 173:26]
  assign io_out_req_bits_wdata = _in_req_bits_T ? io_in_req_bits_wdata : in_req_bits_r_wdata; // @[Utils.scala 50:8]
  assign io_out_req_bits_wmask = _in_req_bits_T ? io_in_req_bits_wmask : in_req_bits_r_wmask; // @[Utils.scala 50:8]
  assign io_out_req_bits_wen = _in_req_bits_T ? io_in_req_bits_wen : in_req_bits_r_wen; // @[Utils.scala 50:8]
  assign io_out_req_bits_len = _in_req_bits_T ? io_in_req_bits_len : in_req_bits_r_len; // @[Utils.scala 50:8]
  assign io_out_req_bits_lrsc = _in_req_bits_T ? io_in_req_bits_lrsc : in_req_bits_r_lrsc; // @[Utils.scala 50:8]
  assign io_out_req_bits_amo = _in_req_bits_T ? io_in_req_bits_amo : in_req_bits_r_amo; // @[Utils.scala 50:8]
  assign io_out_resp_ready = io_in_resp_ready; // @[CachePortProxy.scala 186:32]
  assign io_ptw_req_valid = state == 3'h1; // @[CachePortProxy.scala 113:31]
  assign io_ptw_req_bits_addr = {{7'd0}, _io_ptw_req_bits_addr_T_5}; // @[CachePortProxy.scala 104:24]
  assign io_ptw_resp_ready = state == 3'h2; // @[CachePortProxy.scala 114:31]
  assign tlb_clock = clock;
  assign tlb_reset = reset;
  assign tlb_io_sfence_vma = io_sfence_vma; // @[CachePortProxy.scala 31:21]
  assign tlb_io_vaddr_vpn2 = io_in_req_bits_addr[38:30]; // @[CachePortProxy.scala 32:52]
  assign tlb_io_vaddr_vpn1 = io_in_req_bits_addr[29:21]; // @[CachePortProxy.scala 32:52]
  assign tlb_io_vaddr_vpn0 = io_in_req_bits_addr[20:12]; // @[CachePortProxy.scala 32:52]
  assign tlb_io_wen = _T_30 & ~page_fault; // @[CachePortProxy.scala 121:47]
  assign tlb_io_wvaddr_vpn2 = _GEN_0[38:30]; // @[CachePortProxy.scala 25:46]
  assign tlb_io_wvaddr_vpn1 = _GEN_0[29:21]; // @[CachePortProxy.scala 25:46]
  assign tlb_io_wvaddr_vpn0 = _GEN_0[20:12]; // @[CachePortProxy.scala 25:46]
  assign tlb_io_wpte_ppn2 = ptw_pte_reg_ppn2; // @[CachePortProxy.scala 123:17]
  assign tlb_io_wpte_ppn1 = ptw_pte_reg_ppn1; // @[CachePortProxy.scala 123:17]
  assign tlb_io_wpte_ppn0 = ptw_pte_reg_ppn0; // @[CachePortProxy.scala 123:17]
  assign tlb_io_wpte_flag_d = ptw_pte_reg_flag_d; // @[CachePortProxy.scala 123:17]
  assign tlb_io_wpte_flag_a = ptw_pte_reg_flag_a; // @[CachePortProxy.scala 123:17]
  assign tlb_io_wpte_flag_g = ptw_pte_reg_flag_g; // @[CachePortProxy.scala 123:17]
  assign tlb_io_wpte_flag_u = ptw_pte_reg_flag_u; // @[CachePortProxy.scala 123:17]
  assign tlb_io_wpte_flag_x = ptw_pte_reg_flag_x; // @[CachePortProxy.scala 123:17]
  assign tlb_io_wpte_flag_w = ptw_pte_reg_flag_w; // @[CachePortProxy.scala 123:17]
  assign tlb_io_wpte_flag_r = ptw_pte_reg_flag_r; // @[CachePortProxy.scala 123:17]
  assign tlb_io_wpte_flag_v = ptw_pte_reg_flag_v; // @[CachePortProxy.scala 123:17]
  assign tlb_io_wlevel = ptw_level; // @[CachePortProxy.scala 124:17]
  assign tlb_io_satp_asid = io_satp_asid; // @[CachePortProxy.scala 30:21]
  always @(posedge clock) begin
    if (reset) begin // @[CachePortProxy.scala 21:93]
      state <= 3'h0; // @[CachePortProxy.scala 21:93]
    end else if (3'h0 == state) begin // @[CachePortProxy.scala 52:17]
      if (io_in_req_valid) begin // @[CachePortProxy.scala 59:29]
        if (_access_fault_T_3 & access_fault) begin // @[CachePortProxy.scala 60:39]
          state <= 3'h4; // @[CachePortProxy.scala 61:17]
        end else begin
          state <= _GEN_21;
        end
      end else begin
        state <= _GEN_21;
      end
    end else if (3'h1 == state) begin // @[CachePortProxy.scala 52:17]
      if (_T_7) begin // @[CachePortProxy.scala 67:29]
        state <= 3'h2; // @[CachePortProxy.scala 68:15]
      end
    end else if (3'h2 == state) begin // @[CachePortProxy.scala 52:17]
      state <= _GEN_27;
    end else begin
      state <= _GEN_32;
    end
    if (reset) begin // @[Reg.scala 35:20]
      in_req_bits_r_addr <= 39'h0; // @[Reg.scala 35:20]
    end else if (_in_req_bits_T) begin // @[Reg.scala 36:18]
      in_req_bits_r_addr <= io_in_req_bits_addr; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      in_req_bits_r_wdata <= 64'h0; // @[Reg.scala 35:20]
    end else if (_in_req_bits_T) begin // @[Reg.scala 36:18]
      in_req_bits_r_wdata <= io_in_req_bits_wdata; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      in_req_bits_r_wmask <= 8'h0; // @[Reg.scala 35:20]
    end else if (_in_req_bits_T) begin // @[Reg.scala 36:18]
      in_req_bits_r_wmask <= io_in_req_bits_wmask; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      in_req_bits_r_wen <= 1'h0; // @[Reg.scala 35:20]
    end else if (_in_req_bits_T) begin // @[Reg.scala 36:18]
      in_req_bits_r_wen <= io_in_req_bits_wen; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      in_req_bits_r_len <= 2'h0; // @[Reg.scala 35:20]
    end else if (_in_req_bits_T) begin // @[Reg.scala 36:18]
      in_req_bits_r_len <= io_in_req_bits_len; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      in_req_bits_r_lrsc <= 1'h0; // @[Reg.scala 35:20]
    end else if (_in_req_bits_T) begin // @[Reg.scala 36:18]
      in_req_bits_r_lrsc <= io_in_req_bits_lrsc; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      in_req_bits_r_amo <= 5'h0; // @[Reg.scala 35:20]
    end else if (_in_req_bits_T) begin // @[Reg.scala 36:18]
      in_req_bits_r_amo <= io_in_req_bits_amo; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      atp_en_r <= 1'h0; // @[Reg.scala 35:20]
    end else if (_in_req_bits_T) begin // @[Reg.scala 36:18]
      atp_en_r <= _atp_en_T_1; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[CachePortProxy.scala 46:29]
      ptw_level <= 2'h0; // @[CachePortProxy.scala 46:29]
    end else if (3'h0 == state) begin // @[CachePortProxy.scala 52:17]
      ptw_level <= 2'h2; // @[CachePortProxy.scala 64:17]
    end else if (!(3'h1 == state)) begin // @[CachePortProxy.scala 52:17]
      if (3'h2 == state) begin // @[CachePortProxy.scala 52:17]
        ptw_level <= _GEN_28;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      ptw_pte_reg_ppn2 <= 2'h0; // @[Reg.scala 35:20]
    end else if (_ptw_pte_reg_T) begin // @[Reg.scala 36:18]
      ptw_pte_reg_ppn2 <= ptw_pte_ppn2; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ptw_pte_reg_ppn1 <= 9'h0; // @[Reg.scala 35:20]
    end else if (_ptw_pte_reg_T) begin // @[Reg.scala 36:18]
      ptw_pte_reg_ppn1 <= ptw_pte_ppn1; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ptw_pte_reg_ppn0 <= 9'h0; // @[Reg.scala 35:20]
    end else if (_ptw_pte_reg_T) begin // @[Reg.scala 36:18]
      ptw_pte_reg_ppn0 <= ptw_pte_ppn0; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ptw_pte_reg_flag_d <= 1'h0; // @[Reg.scala 35:20]
    end else if (_ptw_pte_reg_T) begin // @[Reg.scala 36:18]
      ptw_pte_reg_flag_d <= ptw_pte_flag_d; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ptw_pte_reg_flag_a <= 1'h0; // @[Reg.scala 35:20]
    end else if (_ptw_pte_reg_T) begin // @[Reg.scala 36:18]
      ptw_pte_reg_flag_a <= ptw_pte_flag_a; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ptw_pte_reg_flag_g <= 1'h0; // @[Reg.scala 35:20]
    end else if (_ptw_pte_reg_T) begin // @[Reg.scala 36:18]
      ptw_pte_reg_flag_g <= ptw_pte_flag_g; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ptw_pte_reg_flag_u <= 1'h0; // @[Reg.scala 35:20]
    end else if (_ptw_pte_reg_T) begin // @[Reg.scala 36:18]
      ptw_pte_reg_flag_u <= ptw_pte_flag_u; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ptw_pte_reg_flag_x <= 1'h0; // @[Reg.scala 35:20]
    end else if (_ptw_pte_reg_T) begin // @[Reg.scala 36:18]
      ptw_pte_reg_flag_x <= ptw_pte_flag_x; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ptw_pte_reg_flag_w <= 1'h0; // @[Reg.scala 35:20]
    end else if (_ptw_pte_reg_T) begin // @[Reg.scala 36:18]
      ptw_pte_reg_flag_w <= ptw_pte_flag_w; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ptw_pte_reg_flag_r <= 1'h0; // @[Reg.scala 35:20]
    end else if (_ptw_pte_reg_T) begin // @[Reg.scala 36:18]
      ptw_pte_reg_flag_r <= ptw_pte_flag_r; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ptw_pte_reg_flag_v <= 1'h0; // @[Reg.scala 35:20]
    end else if (_ptw_pte_reg_T) begin // @[Reg.scala 36:18]
      ptw_pte_reg_flag_v <= ptw_pte_flag_v; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      prv_r <= 2'h0; // @[Reg.scala 35:20]
    end else if (_in_req_bits_T) begin // @[Utils.scala 50:8]
      prv_r <= io_prv;
    end
    if (reset) begin // @[Utils.scala 36:20]
      page_fault_reg <= 1'h0; // @[Utils.scala 36:20]
    end else if (_T_14) begin // @[Utils.scala 42:18]
      page_fault_reg <= 1'h0; // @[Utils.scala 42:22]
    end else begin
      page_fault_reg <= _GEN_51;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {2{`RANDOM}};
  in_req_bits_r_addr = _RAND_1[38:0];
  _RAND_2 = {2{`RANDOM}};
  in_req_bits_r_wdata = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  in_req_bits_r_wmask = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  in_req_bits_r_wen = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  in_req_bits_r_len = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  in_req_bits_r_lrsc = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  in_req_bits_r_amo = _RAND_7[4:0];
  _RAND_8 = {1{`RANDOM}};
  atp_en_r = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  ptw_level = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  ptw_pte_reg_ppn2 = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  ptw_pte_reg_ppn1 = _RAND_11[8:0];
  _RAND_12 = {1{`RANDOM}};
  ptw_pte_reg_ppn0 = _RAND_12[8:0];
  _RAND_13 = {1{`RANDOM}};
  ptw_pte_reg_flag_d = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  ptw_pte_reg_flag_a = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  ptw_pte_reg_flag_g = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  ptw_pte_reg_flag_u = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  ptw_pte_reg_flag_x = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  ptw_pte_reg_flag_w = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  ptw_pte_reg_flag_r = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  ptw_pte_reg_flag_v = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  prv_r = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  page_fault_reg = _RAND_22[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CachePortXBar1to2(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [38:0] io_in_req_bits_addr,
  input  [63:0] io_in_req_bits_wdata,
  input  [7:0]  io_in_req_bits_wmask,
  input         io_in_req_bits_wen,
  input  [1:0]  io_in_req_bits_len,
  input         io_in_req_bits_lrsc,
  input  [4:0]  io_in_req_bits_amo,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_0_req_ready,
  output        io_out_0_req_valid,
  output [38:0] io_out_0_req_bits_addr,
  output [63:0] io_out_0_req_bits_wdata,
  output [7:0]  io_out_0_req_bits_wmask,
  output        io_out_0_req_bits_wen,
  output [1:0]  io_out_0_req_bits_len,
  output        io_out_0_req_bits_lrsc,
  output [4:0]  io_out_0_req_bits_amo,
  output        io_out_0_resp_ready,
  input         io_out_0_resp_valid,
  input  [63:0] io_out_0_resp_bits_rdata,
  input         io_out_1_req_ready,
  output        io_out_1_req_valid,
  output [38:0] io_out_1_req_bits_addr,
  output [63:0] io_out_1_req_bits_wdata,
  output [7:0]  io_out_1_req_bits_wmask,
  output        io_out_1_req_bits_wen,
  output [1:0]  io_out_1_req_bits_len,
  output        io_out_1_resp_ready,
  input         io_out_1_resp_valid,
  input  [63:0] io_out_1_resp_bits_rdata,
  input         io_to_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  _to_1_r_T = io_in_req_ready & io_in_req_valid; // @[Decoupled.scala 51:35]
  reg  to_1_r; // @[Reg.scala 35:20]
  assign io_in_req_ready = io_to_1 ? io_out_1_req_ready : io_out_0_req_ready; // @[Bus.scala 100:29]
  assign io_in_resp_valid = to_1_r ? io_out_1_resp_valid : io_out_0_resp_valid; // @[Bus.scala 104:30]
  assign io_in_resp_bits_rdata = to_1_r ? io_out_1_resp_bits_rdata : io_out_0_resp_bits_rdata; // @[Bus.scala 103:30]
  assign io_out_0_req_valid = io_in_req_valid & ~io_to_1; // @[Bus.scala 98:42]
  assign io_out_0_req_bits_addr = io_in_req_bits_addr; // @[Bus.scala 96:23]
  assign io_out_0_req_bits_wdata = io_in_req_bits_wdata; // @[Bus.scala 96:23]
  assign io_out_0_req_bits_wmask = io_in_req_bits_wmask; // @[Bus.scala 96:23]
  assign io_out_0_req_bits_wen = io_in_req_bits_wen; // @[Bus.scala 96:23]
  assign io_out_0_req_bits_len = io_in_req_bits_len; // @[Bus.scala 96:23]
  assign io_out_0_req_bits_lrsc = io_in_req_bits_lrsc; // @[Bus.scala 96:23]
  assign io_out_0_req_bits_amo = io_in_req_bits_amo; // @[Bus.scala 96:23]
  assign io_out_0_resp_ready = io_in_resp_ready; // @[Bus.scala 106:24]
  assign io_out_1_req_valid = io_in_req_valid & io_to_1; // @[Bus.scala 99:42]
  assign io_out_1_req_bits_addr = io_in_req_bits_addr; // @[Bus.scala 97:23]
  assign io_out_1_req_bits_wdata = io_in_req_bits_wdata; // @[Bus.scala 97:23]
  assign io_out_1_req_bits_wmask = io_in_req_bits_wmask; // @[Bus.scala 97:23]
  assign io_out_1_req_bits_wen = io_in_req_bits_wen; // @[Bus.scala 97:23]
  assign io_out_1_req_bits_len = io_in_req_bits_len; // @[Bus.scala 97:23]
  assign io_out_1_resp_ready = io_in_resp_ready; // @[Bus.scala 107:24]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 35:20]
      to_1_r <= 1'h0; // @[Reg.scala 35:20]
    end else if (_to_1_r_T) begin // @[Reg.scala 36:18]
      to_1_r <= io_to_1; // @[Reg.scala 36:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  to_1_r = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PipelineReg_1(
  input         clock,
  input         reset,
  input         io_in_uop_valid,
  input  [4:0]  io_in_uop_rd_index,
  input         io_in_uop_rd_wen,
  input  [63:0] io_in_rd_data,
  output        io_out_uop_valid,
  output [4:0]  io_out_uop_rd_index,
  output        io_out_uop_rd_wen,
  output [63:0] io_out_rd_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg  reg_uop_valid; // @[Reg.scala 35:20]
  reg [4:0] reg_uop_rd_index; // @[Reg.scala 35:20]
  reg  reg_uop_rd_wen; // @[Reg.scala 35:20]
  reg [63:0] reg_rd_data; // @[Reg.scala 35:20]
  assign io_out_uop_valid = reg_uop_valid; // @[DataType.scala 41:10]
  assign io_out_uop_rd_index = reg_uop_rd_index; // @[DataType.scala 41:10]
  assign io_out_uop_rd_wen = reg_uop_rd_wen; // @[DataType.scala 41:10]
  assign io_out_rd_data = reg_rd_data; // @[DataType.scala 41:10]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 35:20]
      reg_uop_valid <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      reg_uop_valid <= io_in_uop_valid;
    end
    if (reset) begin // @[Reg.scala 35:20]
      reg_uop_rd_index <= 5'h0; // @[Reg.scala 35:20]
    end else begin
      reg_uop_rd_index <= io_in_uop_rd_index;
    end
    if (reset) begin // @[Reg.scala 35:20]
      reg_uop_rd_wen <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      reg_uop_rd_wen <= io_in_uop_rd_wen;
    end
    if (reset) begin // @[Reg.scala 35:20]
      reg_rd_data <= 64'h0; // @[Reg.scala 35:20]
    end else begin
      reg_rd_data <= io_in_rd_data;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_uop_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  reg_uop_rd_index = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  reg_uop_rd_wen = _RAND_2[0:0];
  _RAND_3 = {2{`RANDOM}};
  reg_rd_data = _RAND_3[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Core(
  input         clock,
  input         reset,
  input         io_imem_req_ready,
  output        io_imem_req_valid,
  output [38:0] io_imem_req_bits_addr,
  output        io_imem_resp_ready,
  input         io_imem_resp_valid,
  input  [63:0] io_imem_resp_bits_rdata,
  input         io_dmem_req_ready,
  output        io_dmem_req_valid,
  output [38:0] io_dmem_req_bits_addr,
  output [63:0] io_dmem_req_bits_wdata,
  output [7:0]  io_dmem_req_bits_wmask,
  output        io_dmem_req_bits_wen,
  output [1:0]  io_dmem_req_bits_len,
  output        io_dmem_req_bits_lrsc,
  output [4:0]  io_dmem_req_bits_amo,
  output        io_dmem_resp_ready,
  input         io_dmem_resp_valid,
  input  [63:0] io_dmem_resp_bits_rdata,
  input         io_iptw_req_ready,
  output        io_iptw_req_valid,
  output [38:0] io_iptw_req_bits_addr,
  output        io_iptw_resp_ready,
  input         io_iptw_resp_valid,
  input  [63:0] io_iptw_resp_bits_rdata,
  input         io_dptw_req_ready,
  output        io_dptw_req_valid,
  output [38:0] io_dptw_req_bits_addr,
  output        io_dptw_resp_ready,
  input         io_dptw_resp_valid,
  input  [63:0] io_dptw_resp_bits_rdata,
  input         io_uncache_req_ready,
  output        io_uncache_req_valid,
  output [38:0] io_uncache_req_bits_addr,
  output [63:0] io_uncache_req_bits_wdata,
  output [7:0]  io_uncache_req_bits_wmask,
  output        io_uncache_req_bits_wen,
  output [1:0]  io_uncache_req_bits_len,
  output        io_uncache_resp_ready,
  input         io_uncache_resp_valid,
  input  [63:0] io_uncache_resp_bits_rdata,
  output        io_fence_i,
  input         io_intr_mtip,
  input         io_intr_msip,
  input         io_intr_meip,
  input         io_intr_seip
);
  wire  ifu_clock; // @[Core.scala 27:19]
  wire  ifu_reset; // @[Core.scala 27:19]
  wire  ifu_io_jmp_packet_valid; // @[Core.scala 27:19]
  wire [63:0] ifu_io_jmp_packet_target; // @[Core.scala 27:19]
  wire  ifu_io_jmp_packet_bp_update; // @[Core.scala 27:19]
  wire  ifu_io_jmp_packet_bp_taken; // @[Core.scala 27:19]
  wire [63:0] ifu_io_jmp_packet_bp_pc; // @[Core.scala 27:19]
  wire  ifu_io_imem_req_ready; // @[Core.scala 27:19]
  wire  ifu_io_imem_req_valid; // @[Core.scala 27:19]
  wire [38:0] ifu_io_imem_req_bits_addr; // @[Core.scala 27:19]
  wire  ifu_io_imem_resp_ready; // @[Core.scala 27:19]
  wire  ifu_io_imem_resp_valid; // @[Core.scala 27:19]
  wire [63:0] ifu_io_imem_resp_bits_rdata; // @[Core.scala 27:19]
  wire  ifu_io_imem_resp_bits_page_fault; // @[Core.scala 27:19]
  wire  ifu_io_imem_resp_bits_access_fault; // @[Core.scala 27:19]
  wire [63:0] ifu_io_out_pc; // @[Core.scala 27:19]
  wire [31:0] ifu_io_out_instr; // @[Core.scala 27:19]
  wire  ifu_io_out_valid; // @[Core.scala 27:19]
  wire  ifu_io_out_page_fault; // @[Core.scala 27:19]
  wire  ifu_io_out_access_fault; // @[Core.scala 27:19]
  wire [63:0] ifu_io_out_bp_npc; // @[Core.scala 27:19]
  wire  ifu_io_stall_b; // @[Core.scala 27:19]
  wire  imem_proxy_clock; // @[Core.scala 28:26]
  wire  imem_proxy_reset; // @[Core.scala 28:26]
  wire [1:0] imem_proxy_io_prv; // @[Core.scala 28:26]
  wire  imem_proxy_io_sv39_en; // @[Core.scala 28:26]
  wire [15:0] imem_proxy_io_satp_asid; // @[Core.scala 28:26]
  wire [43:0] imem_proxy_io_satp_ppn; // @[Core.scala 28:26]
  wire  imem_proxy_io_sfence_vma; // @[Core.scala 28:26]
  wire  imem_proxy_io_in_req_ready; // @[Core.scala 28:26]
  wire  imem_proxy_io_in_req_valid; // @[Core.scala 28:26]
  wire [38:0] imem_proxy_io_in_req_bits_addr; // @[Core.scala 28:26]
  wire  imem_proxy_io_in_resp_ready; // @[Core.scala 28:26]
  wire  imem_proxy_io_in_resp_valid; // @[Core.scala 28:26]
  wire [63:0] imem_proxy_io_in_resp_bits_rdata; // @[Core.scala 28:26]
  wire  imem_proxy_io_in_resp_bits_page_fault; // @[Core.scala 28:26]
  wire  imem_proxy_io_in_resp_bits_access_fault; // @[Core.scala 28:26]
  wire  imem_proxy_io_out_req_ready; // @[Core.scala 28:26]
  wire  imem_proxy_io_out_req_valid; // @[Core.scala 28:26]
  wire [38:0] imem_proxy_io_out_req_bits_addr; // @[Core.scala 28:26]
  wire  imem_proxy_io_out_resp_ready; // @[Core.scala 28:26]
  wire  imem_proxy_io_out_resp_valid; // @[Core.scala 28:26]
  wire [63:0] imem_proxy_io_out_resp_bits_rdata; // @[Core.scala 28:26]
  wire  imem_proxy_io_ptw_req_ready; // @[Core.scala 28:26]
  wire  imem_proxy_io_ptw_req_valid; // @[Core.scala 28:26]
  wire [38:0] imem_proxy_io_ptw_req_bits_addr; // @[Core.scala 28:26]
  wire  imem_proxy_io_ptw_resp_ready; // @[Core.scala 28:26]
  wire  imem_proxy_io_ptw_resp_valid; // @[Core.scala 28:26]
  wire [63:0] imem_proxy_io_ptw_resp_bits_rdata; // @[Core.scala 28:26]
  wire  instr_buffer_clock; // @[Core.scala 54:28]
  wire  instr_buffer_reset; // @[Core.scala 54:28]
  wire  instr_buffer_io_enq_ready; // @[Core.scala 54:28]
  wire  instr_buffer_io_enq_valid; // @[Core.scala 54:28]
  wire [63:0] instr_buffer_io_enq_bits_pc; // @[Core.scala 54:28]
  wire [31:0] instr_buffer_io_enq_bits_instr; // @[Core.scala 54:28]
  wire  instr_buffer_io_enq_bits_page_fault; // @[Core.scala 54:28]
  wire  instr_buffer_io_enq_bits_access_fault; // @[Core.scala 54:28]
  wire [63:0] instr_buffer_io_enq_bits_bp_npc; // @[Core.scala 54:28]
  wire  instr_buffer_io_deq_ready; // @[Core.scala 54:28]
  wire  instr_buffer_io_deq_valid; // @[Core.scala 54:28]
  wire [63:0] instr_buffer_io_deq_bits_pc; // @[Core.scala 54:28]
  wire [31:0] instr_buffer_io_deq_bits_instr; // @[Core.scala 54:28]
  wire  instr_buffer_io_deq_bits_page_fault; // @[Core.scala 54:28]
  wire  instr_buffer_io_deq_bits_access_fault; // @[Core.scala 54:28]
  wire [63:0] instr_buffer_io_deq_bits_bp_npc; // @[Core.scala 54:28]
  wire  instr_buffer_io_flush; // @[Core.scala 54:28]
  wire [63:0] decode_io_in_pc; // @[Core.scala 63:22]
  wire [31:0] decode_io_in_instr; // @[Core.scala 63:22]
  wire  decode_io_in_valid; // @[Core.scala 63:22]
  wire  decode_io_in_page_fault; // @[Core.scala 63:22]
  wire  decode_io_in_access_fault; // @[Core.scala 63:22]
  wire  decode_io_out_valid; // @[Core.scala 63:22]
  wire [2:0] decode_io_out_exc; // @[Core.scala 63:22]
  wire [63:0] decode_io_out_pc; // @[Core.scala 63:22]
  wire [63:0] decode_io_out_npc; // @[Core.scala 63:22]
  wire [31:0] decode_io_out_instr; // @[Core.scala 63:22]
  wire [2:0] decode_io_out_fu; // @[Core.scala 63:22]
  wire [3:0] decode_io_out_alu_op; // @[Core.scala 63:22]
  wire [1:0] decode_io_out_jmp_op; // @[Core.scala 63:22]
  wire [3:0] decode_io_out_mdu_op; // @[Core.scala 63:22]
  wire [4:0] decode_io_out_lsu_op; // @[Core.scala 63:22]
  wire [1:0] decode_io_out_mem_len; // @[Core.scala 63:22]
  wire [1:0] decode_io_out_csr_op; // @[Core.scala 63:22]
  wire [2:0] decode_io_out_sys_op; // @[Core.scala 63:22]
  wire [1:0] decode_io_out_rs1_src; // @[Core.scala 63:22]
  wire [1:0] decode_io_out_rs2_src; // @[Core.scala 63:22]
  wire [4:0] decode_io_out_rs1_index; // @[Core.scala 63:22]
  wire [4:0] decode_io_out_rs2_index; // @[Core.scala 63:22]
  wire [4:0] decode_io_out_rd_index; // @[Core.scala 63:22]
  wire  decode_io_out_rd_wen; // @[Core.scala 63:22]
  wire [31:0] decode_io_out_imm; // @[Core.scala 63:22]
  wire  decode_io_out_dw; // @[Core.scala 63:22]
  wire  rf_clock; // @[Core.scala 67:18]
  wire  rf_reset; // @[Core.scala 67:18]
  wire [4:0] rf_io_rs1_index; // @[Core.scala 67:18]
  wire [4:0] rf_io_rs2_index; // @[Core.scala 67:18]
  wire [63:0] rf_io_rs1_data; // @[Core.scala 67:18]
  wire [63:0] rf_io_rs2_data; // @[Core.scala 67:18]
  wire [4:0] rf_io_rd_index; // @[Core.scala 67:18]
  wire [63:0] rf_io_rd_data; // @[Core.scala 67:18]
  wire  rf_io_rd_wen; // @[Core.scala 67:18]
  wire  id_ex_clock; // @[Core.scala 74:35]
  wire  id_ex_reset; // @[Core.scala 74:35]
  wire  id_ex_io_in_uop_valid; // @[Core.scala 74:35]
  wire [2:0] id_ex_io_in_uop_exc; // @[Core.scala 74:35]
  wire [63:0] id_ex_io_in_uop_pc; // @[Core.scala 74:35]
  wire [63:0] id_ex_io_in_uop_npc; // @[Core.scala 74:35]
  wire [31:0] id_ex_io_in_uop_instr; // @[Core.scala 74:35]
  wire [2:0] id_ex_io_in_uop_fu; // @[Core.scala 74:35]
  wire [3:0] id_ex_io_in_uop_alu_op; // @[Core.scala 74:35]
  wire [1:0] id_ex_io_in_uop_jmp_op; // @[Core.scala 74:35]
  wire [3:0] id_ex_io_in_uop_mdu_op; // @[Core.scala 74:35]
  wire [4:0] id_ex_io_in_uop_lsu_op; // @[Core.scala 74:35]
  wire [1:0] id_ex_io_in_uop_mem_len; // @[Core.scala 74:35]
  wire [1:0] id_ex_io_in_uop_csr_op; // @[Core.scala 74:35]
  wire [2:0] id_ex_io_in_uop_sys_op; // @[Core.scala 74:35]
  wire [4:0] id_ex_io_in_uop_rd_index; // @[Core.scala 74:35]
  wire  id_ex_io_in_uop_rd_wen; // @[Core.scala 74:35]
  wire [31:0] id_ex_io_in_uop_imm; // @[Core.scala 74:35]
  wire  id_ex_io_in_uop_dw; // @[Core.scala 74:35]
  wire [63:0] id_ex_io_in_rs1_data; // @[Core.scala 74:35]
  wire [63:0] id_ex_io_in_rs2_data; // @[Core.scala 74:35]
  wire [63:0] id_ex_io_in_rs2_data_from_rf; // @[Core.scala 74:35]
  wire [63:0] id_ex_io_in_bp_npc; // @[Core.scala 74:35]
  wire  id_ex_io_out_uop_valid; // @[Core.scala 74:35]
  wire [2:0] id_ex_io_out_uop_exc; // @[Core.scala 74:35]
  wire [63:0] id_ex_io_out_uop_pc; // @[Core.scala 74:35]
  wire [63:0] id_ex_io_out_uop_npc; // @[Core.scala 74:35]
  wire [31:0] id_ex_io_out_uop_instr; // @[Core.scala 74:35]
  wire [2:0] id_ex_io_out_uop_fu; // @[Core.scala 74:35]
  wire [3:0] id_ex_io_out_uop_alu_op; // @[Core.scala 74:35]
  wire [1:0] id_ex_io_out_uop_jmp_op; // @[Core.scala 74:35]
  wire [3:0] id_ex_io_out_uop_mdu_op; // @[Core.scala 74:35]
  wire [4:0] id_ex_io_out_uop_lsu_op; // @[Core.scala 74:35]
  wire [1:0] id_ex_io_out_uop_mem_len; // @[Core.scala 74:35]
  wire [1:0] id_ex_io_out_uop_csr_op; // @[Core.scala 74:35]
  wire [2:0] id_ex_io_out_uop_sys_op; // @[Core.scala 74:35]
  wire [4:0] id_ex_io_out_uop_rd_index; // @[Core.scala 74:35]
  wire  id_ex_io_out_uop_rd_wen; // @[Core.scala 74:35]
  wire [31:0] id_ex_io_out_uop_imm; // @[Core.scala 74:35]
  wire  id_ex_io_out_uop_dw; // @[Core.scala 74:35]
  wire [63:0] id_ex_io_out_rs1_data; // @[Core.scala 74:35]
  wire [63:0] id_ex_io_out_rs2_data; // @[Core.scala 74:35]
  wire [63:0] id_ex_io_out_rs2_data_from_rf; // @[Core.scala 74:35]
  wire [63:0] id_ex_io_out_bp_npc; // @[Core.scala 74:35]
  wire  id_ex_io_en; // @[Core.scala 74:35]
  wire  id_ex_io_flush; // @[Core.scala 74:35]
  wire [3:0] alu_io_uop_alu_op; // @[Core.scala 85:19]
  wire [1:0] alu_io_uop_jmp_op; // @[Core.scala 85:19]
  wire  alu_io_uop_dw; // @[Core.scala 85:19]
  wire [63:0] alu_io_in1; // @[Core.scala 85:19]
  wire [63:0] alu_io_in2; // @[Core.scala 85:19]
  wire [63:0] alu_io_out; // @[Core.scala 85:19]
  wire [63:0] alu_io_adder_out; // @[Core.scala 85:19]
  wire  alu_io_cmp_out; // @[Core.scala 85:19]
  wire  lsu_clock; // @[Core.scala 108:19]
  wire  lsu_reset; // @[Core.scala 108:19]
  wire [4:0] lsu_io_uop_lsu_op; // @[Core.scala 108:19]
  wire [1:0] lsu_io_uop_mem_len; // @[Core.scala 108:19]
  wire  lsu_io_is_mem; // @[Core.scala 108:19]
  wire  lsu_io_is_store; // @[Core.scala 108:19]
  wire  lsu_io_is_amo; // @[Core.scala 108:19]
  wire [63:0] lsu_io_addr; // @[Core.scala 108:19]
  wire [63:0] lsu_io_wdata; // @[Core.scala 108:19]
  wire [63:0] lsu_io_rdata; // @[Core.scala 108:19]
  wire  lsu_io_valid; // @[Core.scala 108:19]
  wire [3:0] lsu_io_exc_code; // @[Core.scala 108:19]
  wire  lsu_io_dmem_req_ready; // @[Core.scala 108:19]
  wire  lsu_io_dmem_req_valid; // @[Core.scala 108:19]
  wire [38:0] lsu_io_dmem_req_bits_addr; // @[Core.scala 108:19]
  wire [63:0] lsu_io_dmem_req_bits_wdata; // @[Core.scala 108:19]
  wire [7:0] lsu_io_dmem_req_bits_wmask; // @[Core.scala 108:19]
  wire  lsu_io_dmem_req_bits_wen; // @[Core.scala 108:19]
  wire [1:0] lsu_io_dmem_req_bits_len; // @[Core.scala 108:19]
  wire  lsu_io_dmem_req_bits_lrsc; // @[Core.scala 108:19]
  wire [4:0] lsu_io_dmem_req_bits_amo; // @[Core.scala 108:19]
  wire  lsu_io_dmem_resp_ready; // @[Core.scala 108:19]
  wire  lsu_io_dmem_resp_valid; // @[Core.scala 108:19]
  wire [63:0] lsu_io_dmem_resp_bits_rdata; // @[Core.scala 108:19]
  wire  lsu_io_dmem_resp_bits_page_fault; // @[Core.scala 108:19]
  wire  lsu_io_dmem_resp_bits_access_fault; // @[Core.scala 108:19]
  wire  lsu_io_ready; // @[Core.scala 108:19]
  wire  mdu_clock; // @[Core.scala 116:19]
  wire  mdu_reset; // @[Core.scala 116:19]
  wire  mdu_io_uop_valid; // @[Core.scala 116:19]
  wire [3:0] mdu_io_uop_mdu_op; // @[Core.scala 116:19]
  wire  mdu_io_uop_dw; // @[Core.scala 116:19]
  wire  mdu_io_is_mdu; // @[Core.scala 116:19]
  wire [63:0] mdu_io_in1; // @[Core.scala 116:19]
  wire [63:0] mdu_io_in2; // @[Core.scala 116:19]
  wire [63:0] mdu_io_out; // @[Core.scala 116:19]
  wire  mdu_io_valid; // @[Core.scala 116:19]
  wire  mdu_io_ready; // @[Core.scala 116:19]
  wire  csr_clock; // @[Core.scala 122:19]
  wire  csr_reset; // @[Core.scala 122:19]
  wire  csr_io_uop_valid; // @[Core.scala 122:19]
  wire [2:0] csr_io_uop_exc; // @[Core.scala 122:19]
  wire [63:0] csr_io_uop_pc; // @[Core.scala 122:19]
  wire [63:0] csr_io_uop_npc; // @[Core.scala 122:19]
  wire [2:0] csr_io_uop_fu; // @[Core.scala 122:19]
  wire [2:0] csr_io_uop_sys_op; // @[Core.scala 122:19]
  wire [11:0] csr_io_rw_addr; // @[Core.scala 122:19]
  wire [1:0] csr_io_rw_cmd; // @[Core.scala 122:19]
  wire [63:0] csr_io_rw_wdata; // @[Core.scala 122:19]
  wire [63:0] csr_io_rw_rdata; // @[Core.scala 122:19]
  wire  csr_io_rw_valid; // @[Core.scala 122:19]
  wire [1:0] csr_io_prv; // @[Core.scala 122:19]
  wire  csr_io_mprv; // @[Core.scala 122:19]
  wire [1:0] csr_io_mpp; // @[Core.scala 122:19]
  wire  csr_io_sv39_en; // @[Core.scala 122:19]
  wire [15:0] csr_io_satp_asid; // @[Core.scala 122:19]
  wire [43:0] csr_io_satp_ppn; // @[Core.scala 122:19]
  wire  csr_io_sfence_vma; // @[Core.scala 122:19]
  wire  csr_io_fence_i; // @[Core.scala 122:19]
  wire  csr_io_jmp_packet_valid; // @[Core.scala 122:19]
  wire [63:0] csr_io_jmp_packet_target; // @[Core.scala 122:19]
  wire [63:0] csr_io_lsu_addr; // @[Core.scala 122:19]
  wire [3:0] csr_io_lsu_exc_code; // @[Core.scala 122:19]
  wire  csr_io_interrupt_mtip; // @[Core.scala 122:19]
  wire  csr_io_interrupt_msip; // @[Core.scala 122:19]
  wire  csr_io_interrupt_meip; // @[Core.scala 122:19]
  wire  csr_io_interrupt_seip; // @[Core.scala 122:19]
  wire  csr_io_is_int; // @[Core.scala 122:19]
  wire  csr_io_commit; // @[Core.scala 122:19]
  wire  dmem_proxy_clock; // @[Core.scala 142:26]
  wire  dmem_proxy_reset; // @[Core.scala 142:26]
  wire [1:0] dmem_proxy_io_prv; // @[Core.scala 142:26]
  wire  dmem_proxy_io_sv39_en; // @[Core.scala 142:26]
  wire [15:0] dmem_proxy_io_satp_asid; // @[Core.scala 142:26]
  wire [43:0] dmem_proxy_io_satp_ppn; // @[Core.scala 142:26]
  wire  dmem_proxy_io_sfence_vma; // @[Core.scala 142:26]
  wire  dmem_proxy_io_in_req_ready; // @[Core.scala 142:26]
  wire  dmem_proxy_io_in_req_valid; // @[Core.scala 142:26]
  wire [38:0] dmem_proxy_io_in_req_bits_addr; // @[Core.scala 142:26]
  wire [63:0] dmem_proxy_io_in_req_bits_wdata; // @[Core.scala 142:26]
  wire [7:0] dmem_proxy_io_in_req_bits_wmask; // @[Core.scala 142:26]
  wire  dmem_proxy_io_in_req_bits_wen; // @[Core.scala 142:26]
  wire [1:0] dmem_proxy_io_in_req_bits_len; // @[Core.scala 142:26]
  wire  dmem_proxy_io_in_req_bits_lrsc; // @[Core.scala 142:26]
  wire [4:0] dmem_proxy_io_in_req_bits_amo; // @[Core.scala 142:26]
  wire  dmem_proxy_io_in_resp_ready; // @[Core.scala 142:26]
  wire  dmem_proxy_io_in_resp_valid; // @[Core.scala 142:26]
  wire [63:0] dmem_proxy_io_in_resp_bits_rdata; // @[Core.scala 142:26]
  wire  dmem_proxy_io_in_resp_bits_page_fault; // @[Core.scala 142:26]
  wire  dmem_proxy_io_in_resp_bits_access_fault; // @[Core.scala 142:26]
  wire  dmem_proxy_io_out_req_ready; // @[Core.scala 142:26]
  wire  dmem_proxy_io_out_req_valid; // @[Core.scala 142:26]
  wire [38:0] dmem_proxy_io_out_req_bits_addr; // @[Core.scala 142:26]
  wire [63:0] dmem_proxy_io_out_req_bits_wdata; // @[Core.scala 142:26]
  wire [7:0] dmem_proxy_io_out_req_bits_wmask; // @[Core.scala 142:26]
  wire  dmem_proxy_io_out_req_bits_wen; // @[Core.scala 142:26]
  wire [1:0] dmem_proxy_io_out_req_bits_len; // @[Core.scala 142:26]
  wire  dmem_proxy_io_out_req_bits_lrsc; // @[Core.scala 142:26]
  wire [4:0] dmem_proxy_io_out_req_bits_amo; // @[Core.scala 142:26]
  wire  dmem_proxy_io_out_resp_ready; // @[Core.scala 142:26]
  wire  dmem_proxy_io_out_resp_valid; // @[Core.scala 142:26]
  wire [63:0] dmem_proxy_io_out_resp_bits_rdata; // @[Core.scala 142:26]
  wire  dmem_proxy_io_ptw_req_ready; // @[Core.scala 142:26]
  wire  dmem_proxy_io_ptw_req_valid; // @[Core.scala 142:26]
  wire [38:0] dmem_proxy_io_ptw_req_bits_addr; // @[Core.scala 142:26]
  wire  dmem_proxy_io_ptw_resp_ready; // @[Core.scala 142:26]
  wire  dmem_proxy_io_ptw_resp_valid; // @[Core.scala 142:26]
  wire [63:0] dmem_proxy_io_ptw_resp_bits_rdata; // @[Core.scala 142:26]
  wire  c2_xbar_clock; // @[Core.scala 164:23]
  wire  c2_xbar_reset; // @[Core.scala 164:23]
  wire  c2_xbar_io_in_req_ready; // @[Core.scala 164:23]
  wire  c2_xbar_io_in_req_valid; // @[Core.scala 164:23]
  wire [38:0] c2_xbar_io_in_req_bits_addr; // @[Core.scala 164:23]
  wire [63:0] c2_xbar_io_in_req_bits_wdata; // @[Core.scala 164:23]
  wire [7:0] c2_xbar_io_in_req_bits_wmask; // @[Core.scala 164:23]
  wire  c2_xbar_io_in_req_bits_wen; // @[Core.scala 164:23]
  wire [1:0] c2_xbar_io_in_req_bits_len; // @[Core.scala 164:23]
  wire  c2_xbar_io_in_req_bits_lrsc; // @[Core.scala 164:23]
  wire [4:0] c2_xbar_io_in_req_bits_amo; // @[Core.scala 164:23]
  wire  c2_xbar_io_in_resp_ready; // @[Core.scala 164:23]
  wire  c2_xbar_io_in_resp_valid; // @[Core.scala 164:23]
  wire [63:0] c2_xbar_io_in_resp_bits_rdata; // @[Core.scala 164:23]
  wire  c2_xbar_io_out_0_req_ready; // @[Core.scala 164:23]
  wire  c2_xbar_io_out_0_req_valid; // @[Core.scala 164:23]
  wire [38:0] c2_xbar_io_out_0_req_bits_addr; // @[Core.scala 164:23]
  wire [63:0] c2_xbar_io_out_0_req_bits_wdata; // @[Core.scala 164:23]
  wire [7:0] c2_xbar_io_out_0_req_bits_wmask; // @[Core.scala 164:23]
  wire  c2_xbar_io_out_0_req_bits_wen; // @[Core.scala 164:23]
  wire [1:0] c2_xbar_io_out_0_req_bits_len; // @[Core.scala 164:23]
  wire  c2_xbar_io_out_0_req_bits_lrsc; // @[Core.scala 164:23]
  wire [4:0] c2_xbar_io_out_0_req_bits_amo; // @[Core.scala 164:23]
  wire  c2_xbar_io_out_0_resp_ready; // @[Core.scala 164:23]
  wire  c2_xbar_io_out_0_resp_valid; // @[Core.scala 164:23]
  wire [63:0] c2_xbar_io_out_0_resp_bits_rdata; // @[Core.scala 164:23]
  wire  c2_xbar_io_out_1_req_ready; // @[Core.scala 164:23]
  wire  c2_xbar_io_out_1_req_valid; // @[Core.scala 164:23]
  wire [38:0] c2_xbar_io_out_1_req_bits_addr; // @[Core.scala 164:23]
  wire [63:0] c2_xbar_io_out_1_req_bits_wdata; // @[Core.scala 164:23]
  wire [7:0] c2_xbar_io_out_1_req_bits_wmask; // @[Core.scala 164:23]
  wire  c2_xbar_io_out_1_req_bits_wen; // @[Core.scala 164:23]
  wire [1:0] c2_xbar_io_out_1_req_bits_len; // @[Core.scala 164:23]
  wire  c2_xbar_io_out_1_resp_ready; // @[Core.scala 164:23]
  wire  c2_xbar_io_out_1_resp_valid; // @[Core.scala 164:23]
  wire [63:0] c2_xbar_io_out_1_resp_bits_rdata; // @[Core.scala 164:23]
  wire  c2_xbar_io_to_1; // @[Core.scala 164:23]
  wire  ex_wb_clock; // @[Core.scala 172:21]
  wire  ex_wb_reset; // @[Core.scala 172:21]
  wire  ex_wb_io_in_uop_valid; // @[Core.scala 172:21]
  wire [4:0] ex_wb_io_in_uop_rd_index; // @[Core.scala 172:21]
  wire  ex_wb_io_in_uop_rd_wen; // @[Core.scala 172:21]
  wire [63:0] ex_wb_io_in_rd_data; // @[Core.scala 172:21]
  wire  ex_wb_io_out_uop_valid; // @[Core.scala 172:21]
  wire [4:0] ex_wb_io_out_uop_rd_index; // @[Core.scala 172:21]
  wire  ex_wb_io_out_uop_rd_wen; // @[Core.scala 172:21]
  wire [63:0] ex_wb_io_out_rd_data; // @[Core.scala 172:21]
  wire  alu_jmp_packet_bp_update = id_ex_io_out_uop_valid & alu_io_uop_jmp_op != 2'h0; // @[Core.scala 96:54]
  wire  _alu_jmp_packet_target_T_5 = ~alu_io_uop_jmp_op[1] & alu_io_uop_jmp_op[0]; // @[Constant.scala 52:47]
  wire [31:0] _alu_jmp_packet_target_T_8 = id_ex_io_out_uop_imm[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _alu_jmp_packet_target_T_9 = {_alu_jmp_packet_target_T_8,id_ex_io_out_uop_imm}; // @[Cat.scala 33:92]
  wire [63:0] _alu_jmp_packet_target_T_11 = id_ex_io_out_uop_pc + _alu_jmp_packet_target_T_9; // @[Core.scala 93:45]
  wire [63:0] _alu_jmp_packet_target_T_12 = alu_io_cmp_out ? _alu_jmp_packet_target_T_11 : id_ex_io_out_uop_npc; // @[Core.scala 93:8]
  wire [63:0] alu_jmp_packet_target = _alu_jmp_packet_target_T_5 ? _alu_jmp_packet_target_T_12 : alu_io_adder_out; // @[Core.scala 91:31]
  wire  alu_jmp_packet_valid = alu_jmp_packet_bp_update & alu_jmp_packet_target != id_ex_io_out_bp_npc; // @[Core.scala 90:52]
  wire  sys_jmp_packet_valid = csr_io_jmp_packet_valid; // @[Core.scala 127:23 42:28]
  wire [63:0] sys_jmp_packet_target = csr_io_jmp_packet_target; // @[Core.scala 127:23 42:28]
  wire [63:0] alu_br_out = id_ex_io_out_uop_jmp_op[1] ? id_ex_io_out_uop_npc : alu_io_out; // @[Core.scala 100:23]
  wire  is_mem = id_ex_io_out_uop_fu == 3'h3 & id_ex_io_out_uop_valid; // @[Core.scala 102:58]
  wire  is_mdu = id_ex_io_out_uop_fu == 3'h2 & id_ex_io_out_uop_valid; // @[Core.scala 103:58]
  wire  is_csr = id_ex_io_out_uop_fu == 3'h4 & id_ex_io_out_uop_valid; // @[Core.scala 104:58]
  wire [1:0] prv = csr_io_prv; // @[Core.scala 128:23 19:24]
  wire  _ex_wb_io_in_uop_valid_T_3 = is_mdu & mdu_io_valid; // @[Core.scala 176:15]
  wire  _ex_wb_io_in_uop_valid_T_4 = is_mem & lsu_io_valid & lsu_io_exc_code == 4'h0 | _ex_wb_io_in_uop_valid_T_3; // @[Core.scala 175:59]
  wire  _ex_wb_io_in_uop_valid_T_5 = is_csr & csr_io_rw_valid; // @[Core.scala 177:15]
  wire  _ex_wb_io_in_uop_valid_T_6 = _ex_wb_io_in_uop_valid_T_4 | _ex_wb_io_in_uop_valid_T_5; // @[Core.scala 176:32]
  wire  _ex_wb_io_in_uop_valid_T_12 = ~is_mem & ~is_mdu & ~is_csr & id_ex_io_out_uop_valid; // @[Core.scala 178:38]
  wire  _ex_wb_io_in_uop_valid_T_13 = _ex_wb_io_in_uop_valid_T_6 | _ex_wb_io_in_uop_valid_T_12; // @[Core.scala 177:35]
  wire [63:0] _ex_wb_io_in_rd_data_T_1 = 3'h3 == id_ex_io_out_uop_fu ? lsu_io_rdata : alu_br_out; // @[Mux.scala 81:58]
  wire [63:0] _ex_wb_io_in_rd_data_T_3 = 3'h2 == id_ex_io_out_uop_fu ? mdu_io_out : _ex_wb_io_in_rd_data_T_1; // @[Mux.scala 81:58]
  wire  need_rs1 = decode_io_out_rs1_src == 2'h2; // @[Core.scala 202:40]
  wire  need_rs2 = decode_io_out_rs2_src == 2'h2; // @[Core.scala 203:40]
  wire  _need_rs2_from_rf_T_5 = ~decode_io_out_lsu_op[4] & decode_io_out_lsu_op[0]; // @[Constant.scala 82:45]
  wire  need_rs2_from_rf = _need_rs2_from_rf_T_5 | decode_io_out_lsu_op[4] | decode_io_out_fu == 3'h2; // @[Core.scala 205:66]
  wire  _T = need_rs1 & id_ex_io_out_uop_rd_wen; // @[Core.scala 208:14]
  wire  _T_2 = _T & decode_io_out_rs1_index == id_ex_io_out_uop_rd_index; // @[Core.scala 209:7]
  wire  _T_4 = _T_2 & decode_io_out_rs1_index != 5'h0; // @[Core.scala 210:7]
  wire [95:0] _id_rs1_data_T_1 = {32'h0,instr_buffer_io_deq_bits_pc}; // @[Cat.scala 33:92]
  wire [31:0] _id_rs1_data_T_4 = decode_io_out_imm[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _id_rs1_data_T_5 = {_id_rs1_data_T_4,decode_io_out_imm}; // @[Cat.scala 33:92]
  wire [95:0] _id_rs1_data_T_7 = 2'h1 == decode_io_out_rs1_src ? _id_rs1_data_T_1 : 96'h0; // @[Mux.scala 81:58]
  wire [95:0] _id_rs1_data_T_9 = 2'h2 == decode_io_out_rs1_src ? {{32'd0}, rf_io_rs1_data} : _id_rs1_data_T_7; // @[Mux.scala 81:58]
  wire [95:0] _id_rs1_data_T_11 = 2'h3 == decode_io_out_rs1_src ? {{32'd0}, _id_rs1_data_T_5} : _id_rs1_data_T_9; // @[Mux.scala 81:58]
  wire [95:0] _GEN_0 = _T_4 ? {{32'd0}, ex_wb_io_in_rd_data} : _id_rs1_data_T_11; // @[Core.scala 211:5 212:17 214:17]
  wire  _T_5 = need_rs2 & id_ex_io_out_uop_rd_wen; // @[Core.scala 226:14]
  wire  _T_6 = decode_io_out_rs2_index == id_ex_io_out_uop_rd_index; // @[Core.scala 227:34]
  wire  _T_7 = _T_5 & decode_io_out_rs2_index == id_ex_io_out_uop_rd_index; // @[Core.scala 227:7]
  wire  _T_8 = decode_io_out_rs2_index != 5'h0; // @[Core.scala 228:34]
  wire  _T_9 = _T_7 & decode_io_out_rs2_index != 5'h0; // @[Core.scala 228:7]
  wire [95:0] _id_rs2_data_T_7 = 2'h1 == decode_io_out_rs2_src ? _id_rs1_data_T_1 : 96'h0; // @[Mux.scala 81:58]
  wire [95:0] _id_rs2_data_T_9 = 2'h2 == decode_io_out_rs2_src ? {{32'd0}, rf_io_rs2_data} : _id_rs2_data_T_7; // @[Mux.scala 81:58]
  wire [95:0] _id_rs2_data_T_11 = 2'h3 == decode_io_out_rs2_src ? {{32'd0}, _id_rs1_data_T_5} : _id_rs2_data_T_9; // @[Mux.scala 81:58]
  wire [95:0] _GEN_1 = _T_9 ? {{32'd0}, ex_wb_io_in_rd_data} : _id_rs2_data_T_11; // @[Core.scala 229:5 230:17 232:17]
  wire  _T_10 = need_rs2_from_rf & id_ex_io_out_uop_rd_wen; // @[Core.scala 244:22]
  wire  _T_12 = _T_10 & _T_6; // @[Core.scala 245:7]
  wire  _T_14 = _T_12 & _T_8; // @[Core.scala 246:7]
  IFU ifu ( // @[Core.scala 27:19]
    .clock(ifu_clock),
    .reset(ifu_reset),
    .io_jmp_packet_valid(ifu_io_jmp_packet_valid),
    .io_jmp_packet_target(ifu_io_jmp_packet_target),
    .io_jmp_packet_bp_update(ifu_io_jmp_packet_bp_update),
    .io_jmp_packet_bp_taken(ifu_io_jmp_packet_bp_taken),
    .io_jmp_packet_bp_pc(ifu_io_jmp_packet_bp_pc),
    .io_imem_req_ready(ifu_io_imem_req_ready),
    .io_imem_req_valid(ifu_io_imem_req_valid),
    .io_imem_req_bits_addr(ifu_io_imem_req_bits_addr),
    .io_imem_resp_ready(ifu_io_imem_resp_ready),
    .io_imem_resp_valid(ifu_io_imem_resp_valid),
    .io_imem_resp_bits_rdata(ifu_io_imem_resp_bits_rdata),
    .io_imem_resp_bits_page_fault(ifu_io_imem_resp_bits_page_fault),
    .io_imem_resp_bits_access_fault(ifu_io_imem_resp_bits_access_fault),
    .io_out_pc(ifu_io_out_pc),
    .io_out_instr(ifu_io_out_instr),
    .io_out_valid(ifu_io_out_valid),
    .io_out_page_fault(ifu_io_out_page_fault),
    .io_out_access_fault(ifu_io_out_access_fault),
    .io_out_bp_npc(ifu_io_out_bp_npc),
    .io_stall_b(ifu_io_stall_b)
  );
  CachePortProxy imem_proxy ( // @[Core.scala 28:26]
    .clock(imem_proxy_clock),
    .reset(imem_proxy_reset),
    .io_prv(imem_proxy_io_prv),
    .io_sv39_en(imem_proxy_io_sv39_en),
    .io_satp_asid(imem_proxy_io_satp_asid),
    .io_satp_ppn(imem_proxy_io_satp_ppn),
    .io_sfence_vma(imem_proxy_io_sfence_vma),
    .io_in_req_ready(imem_proxy_io_in_req_ready),
    .io_in_req_valid(imem_proxy_io_in_req_valid),
    .io_in_req_bits_addr(imem_proxy_io_in_req_bits_addr),
    .io_in_resp_ready(imem_proxy_io_in_resp_ready),
    .io_in_resp_valid(imem_proxy_io_in_resp_valid),
    .io_in_resp_bits_rdata(imem_proxy_io_in_resp_bits_rdata),
    .io_in_resp_bits_page_fault(imem_proxy_io_in_resp_bits_page_fault),
    .io_in_resp_bits_access_fault(imem_proxy_io_in_resp_bits_access_fault),
    .io_out_req_ready(imem_proxy_io_out_req_ready),
    .io_out_req_valid(imem_proxy_io_out_req_valid),
    .io_out_req_bits_addr(imem_proxy_io_out_req_bits_addr),
    .io_out_resp_ready(imem_proxy_io_out_resp_ready),
    .io_out_resp_valid(imem_proxy_io_out_resp_valid),
    .io_out_resp_bits_rdata(imem_proxy_io_out_resp_bits_rdata),
    .io_ptw_req_ready(imem_proxy_io_ptw_req_ready),
    .io_ptw_req_valid(imem_proxy_io_ptw_req_valid),
    .io_ptw_req_bits_addr(imem_proxy_io_ptw_req_bits_addr),
    .io_ptw_resp_ready(imem_proxy_io_ptw_resp_ready),
    .io_ptw_resp_valid(imem_proxy_io_ptw_resp_valid),
    .io_ptw_resp_bits_rdata(imem_proxy_io_ptw_resp_bits_rdata)
  );
  Queue_2 instr_buffer ( // @[Core.scala 54:28]
    .clock(instr_buffer_clock),
    .reset(instr_buffer_reset),
    .io_enq_ready(instr_buffer_io_enq_ready),
    .io_enq_valid(instr_buffer_io_enq_valid),
    .io_enq_bits_pc(instr_buffer_io_enq_bits_pc),
    .io_enq_bits_instr(instr_buffer_io_enq_bits_instr),
    .io_enq_bits_page_fault(instr_buffer_io_enq_bits_page_fault),
    .io_enq_bits_access_fault(instr_buffer_io_enq_bits_access_fault),
    .io_enq_bits_bp_npc(instr_buffer_io_enq_bits_bp_npc),
    .io_deq_ready(instr_buffer_io_deq_ready),
    .io_deq_valid(instr_buffer_io_deq_valid),
    .io_deq_bits_pc(instr_buffer_io_deq_bits_pc),
    .io_deq_bits_instr(instr_buffer_io_deq_bits_instr),
    .io_deq_bits_page_fault(instr_buffer_io_deq_bits_page_fault),
    .io_deq_bits_access_fault(instr_buffer_io_deq_bits_access_fault),
    .io_deq_bits_bp_npc(instr_buffer_io_deq_bits_bp_npc),
    .io_flush(instr_buffer_io_flush)
  );
  Decode decode ( // @[Core.scala 63:22]
    .io_in_pc(decode_io_in_pc),
    .io_in_instr(decode_io_in_instr),
    .io_in_valid(decode_io_in_valid),
    .io_in_page_fault(decode_io_in_page_fault),
    .io_in_access_fault(decode_io_in_access_fault),
    .io_out_valid(decode_io_out_valid),
    .io_out_exc(decode_io_out_exc),
    .io_out_pc(decode_io_out_pc),
    .io_out_npc(decode_io_out_npc),
    .io_out_instr(decode_io_out_instr),
    .io_out_fu(decode_io_out_fu),
    .io_out_alu_op(decode_io_out_alu_op),
    .io_out_jmp_op(decode_io_out_jmp_op),
    .io_out_mdu_op(decode_io_out_mdu_op),
    .io_out_lsu_op(decode_io_out_lsu_op),
    .io_out_mem_len(decode_io_out_mem_len),
    .io_out_csr_op(decode_io_out_csr_op),
    .io_out_sys_op(decode_io_out_sys_op),
    .io_out_rs1_src(decode_io_out_rs1_src),
    .io_out_rs2_src(decode_io_out_rs2_src),
    .io_out_rs1_index(decode_io_out_rs1_index),
    .io_out_rs2_index(decode_io_out_rs2_index),
    .io_out_rd_index(decode_io_out_rd_index),
    .io_out_rd_wen(decode_io_out_rd_wen),
    .io_out_imm(decode_io_out_imm),
    .io_out_dw(decode_io_out_dw)
  );
  RegFile rf ( // @[Core.scala 67:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_rs1_index(rf_io_rs1_index),
    .io_rs2_index(rf_io_rs2_index),
    .io_rs1_data(rf_io_rs1_data),
    .io_rs2_data(rf_io_rs2_data),
    .io_rd_index(rf_io_rd_index),
    .io_rd_data(rf_io_rd_data),
    .io_rd_wen(rf_io_rd_wen)
  );
  PipelineReg id_ex ( // @[Core.scala 74:35]
    .clock(id_ex_clock),
    .reset(id_ex_reset),
    .io_in_uop_valid(id_ex_io_in_uop_valid),
    .io_in_uop_exc(id_ex_io_in_uop_exc),
    .io_in_uop_pc(id_ex_io_in_uop_pc),
    .io_in_uop_npc(id_ex_io_in_uop_npc),
    .io_in_uop_instr(id_ex_io_in_uop_instr),
    .io_in_uop_fu(id_ex_io_in_uop_fu),
    .io_in_uop_alu_op(id_ex_io_in_uop_alu_op),
    .io_in_uop_jmp_op(id_ex_io_in_uop_jmp_op),
    .io_in_uop_mdu_op(id_ex_io_in_uop_mdu_op),
    .io_in_uop_lsu_op(id_ex_io_in_uop_lsu_op),
    .io_in_uop_mem_len(id_ex_io_in_uop_mem_len),
    .io_in_uop_csr_op(id_ex_io_in_uop_csr_op),
    .io_in_uop_sys_op(id_ex_io_in_uop_sys_op),
    .io_in_uop_rd_index(id_ex_io_in_uop_rd_index),
    .io_in_uop_rd_wen(id_ex_io_in_uop_rd_wen),
    .io_in_uop_imm(id_ex_io_in_uop_imm),
    .io_in_uop_dw(id_ex_io_in_uop_dw),
    .io_in_rs1_data(id_ex_io_in_rs1_data),
    .io_in_rs2_data(id_ex_io_in_rs2_data),
    .io_in_rs2_data_from_rf(id_ex_io_in_rs2_data_from_rf),
    .io_in_bp_npc(id_ex_io_in_bp_npc),
    .io_out_uop_valid(id_ex_io_out_uop_valid),
    .io_out_uop_exc(id_ex_io_out_uop_exc),
    .io_out_uop_pc(id_ex_io_out_uop_pc),
    .io_out_uop_npc(id_ex_io_out_uop_npc),
    .io_out_uop_instr(id_ex_io_out_uop_instr),
    .io_out_uop_fu(id_ex_io_out_uop_fu),
    .io_out_uop_alu_op(id_ex_io_out_uop_alu_op),
    .io_out_uop_jmp_op(id_ex_io_out_uop_jmp_op),
    .io_out_uop_mdu_op(id_ex_io_out_uop_mdu_op),
    .io_out_uop_lsu_op(id_ex_io_out_uop_lsu_op),
    .io_out_uop_mem_len(id_ex_io_out_uop_mem_len),
    .io_out_uop_csr_op(id_ex_io_out_uop_csr_op),
    .io_out_uop_sys_op(id_ex_io_out_uop_sys_op),
    .io_out_uop_rd_index(id_ex_io_out_uop_rd_index),
    .io_out_uop_rd_wen(id_ex_io_out_uop_rd_wen),
    .io_out_uop_imm(id_ex_io_out_uop_imm),
    .io_out_uop_dw(id_ex_io_out_uop_dw),
    .io_out_rs1_data(id_ex_io_out_rs1_data),
    .io_out_rs2_data(id_ex_io_out_rs2_data),
    .io_out_rs2_data_from_rf(id_ex_io_out_rs2_data_from_rf),
    .io_out_bp_npc(id_ex_io_out_bp_npc),
    .io_en(id_ex_io_en),
    .io_flush(id_ex_io_flush)
  );
  ALU alu ( // @[Core.scala 85:19]
    .io_uop_alu_op(alu_io_uop_alu_op),
    .io_uop_jmp_op(alu_io_uop_jmp_op),
    .io_uop_dw(alu_io_uop_dw),
    .io_in1(alu_io_in1),
    .io_in2(alu_io_in2),
    .io_out(alu_io_out),
    .io_adder_out(alu_io_adder_out),
    .io_cmp_out(alu_io_cmp_out)
  );
  LSU lsu ( // @[Core.scala 108:19]
    .clock(lsu_clock),
    .reset(lsu_reset),
    .io_uop_lsu_op(lsu_io_uop_lsu_op),
    .io_uop_mem_len(lsu_io_uop_mem_len),
    .io_is_mem(lsu_io_is_mem),
    .io_is_store(lsu_io_is_store),
    .io_is_amo(lsu_io_is_amo),
    .io_addr(lsu_io_addr),
    .io_wdata(lsu_io_wdata),
    .io_rdata(lsu_io_rdata),
    .io_valid(lsu_io_valid),
    .io_exc_code(lsu_io_exc_code),
    .io_dmem_req_ready(lsu_io_dmem_req_ready),
    .io_dmem_req_valid(lsu_io_dmem_req_valid),
    .io_dmem_req_bits_addr(lsu_io_dmem_req_bits_addr),
    .io_dmem_req_bits_wdata(lsu_io_dmem_req_bits_wdata),
    .io_dmem_req_bits_wmask(lsu_io_dmem_req_bits_wmask),
    .io_dmem_req_bits_wen(lsu_io_dmem_req_bits_wen),
    .io_dmem_req_bits_len(lsu_io_dmem_req_bits_len),
    .io_dmem_req_bits_lrsc(lsu_io_dmem_req_bits_lrsc),
    .io_dmem_req_bits_amo(lsu_io_dmem_req_bits_amo),
    .io_dmem_resp_ready(lsu_io_dmem_resp_ready),
    .io_dmem_resp_valid(lsu_io_dmem_resp_valid),
    .io_dmem_resp_bits_rdata(lsu_io_dmem_resp_bits_rdata),
    .io_dmem_resp_bits_page_fault(lsu_io_dmem_resp_bits_page_fault),
    .io_dmem_resp_bits_access_fault(lsu_io_dmem_resp_bits_access_fault),
    .io_ready(lsu_io_ready)
  );
  MDU mdu ( // @[Core.scala 116:19]
    .clock(mdu_clock),
    .reset(mdu_reset),
    .io_uop_valid(mdu_io_uop_valid),
    .io_uop_mdu_op(mdu_io_uop_mdu_op),
    .io_uop_dw(mdu_io_uop_dw),
    .io_is_mdu(mdu_io_is_mdu),
    .io_in1(mdu_io_in1),
    .io_in2(mdu_io_in2),
    .io_out(mdu_io_out),
    .io_valid(mdu_io_valid),
    .io_ready(mdu_io_ready)
  );
  CSR csr ( // @[Core.scala 122:19]
    .clock(csr_clock),
    .reset(csr_reset),
    .io_uop_valid(csr_io_uop_valid),
    .io_uop_exc(csr_io_uop_exc),
    .io_uop_pc(csr_io_uop_pc),
    .io_uop_npc(csr_io_uop_npc),
    .io_uop_fu(csr_io_uop_fu),
    .io_uop_sys_op(csr_io_uop_sys_op),
    .io_rw_addr(csr_io_rw_addr),
    .io_rw_cmd(csr_io_rw_cmd),
    .io_rw_wdata(csr_io_rw_wdata),
    .io_rw_rdata(csr_io_rw_rdata),
    .io_rw_valid(csr_io_rw_valid),
    .io_prv(csr_io_prv),
    .io_mprv(csr_io_mprv),
    .io_mpp(csr_io_mpp),
    .io_sv39_en(csr_io_sv39_en),
    .io_satp_asid(csr_io_satp_asid),
    .io_satp_ppn(csr_io_satp_ppn),
    .io_sfence_vma(csr_io_sfence_vma),
    .io_fence_i(csr_io_fence_i),
    .io_jmp_packet_valid(csr_io_jmp_packet_valid),
    .io_jmp_packet_target(csr_io_jmp_packet_target),
    .io_lsu_addr(csr_io_lsu_addr),
    .io_lsu_exc_code(csr_io_lsu_exc_code),
    .io_interrupt_mtip(csr_io_interrupt_mtip),
    .io_interrupt_msip(csr_io_interrupt_msip),
    .io_interrupt_meip(csr_io_interrupt_meip),
    .io_interrupt_seip(csr_io_interrupt_seip),
    .io_is_int(csr_io_is_int),
    .io_commit(csr_io_commit)
  );
  CachePortProxy_1 dmem_proxy ( // @[Core.scala 142:26]
    .clock(dmem_proxy_clock),
    .reset(dmem_proxy_reset),
    .io_prv(dmem_proxy_io_prv),
    .io_sv39_en(dmem_proxy_io_sv39_en),
    .io_satp_asid(dmem_proxy_io_satp_asid),
    .io_satp_ppn(dmem_proxy_io_satp_ppn),
    .io_sfence_vma(dmem_proxy_io_sfence_vma),
    .io_in_req_ready(dmem_proxy_io_in_req_ready),
    .io_in_req_valid(dmem_proxy_io_in_req_valid),
    .io_in_req_bits_addr(dmem_proxy_io_in_req_bits_addr),
    .io_in_req_bits_wdata(dmem_proxy_io_in_req_bits_wdata),
    .io_in_req_bits_wmask(dmem_proxy_io_in_req_bits_wmask),
    .io_in_req_bits_wen(dmem_proxy_io_in_req_bits_wen),
    .io_in_req_bits_len(dmem_proxy_io_in_req_bits_len),
    .io_in_req_bits_lrsc(dmem_proxy_io_in_req_bits_lrsc),
    .io_in_req_bits_amo(dmem_proxy_io_in_req_bits_amo),
    .io_in_resp_ready(dmem_proxy_io_in_resp_ready),
    .io_in_resp_valid(dmem_proxy_io_in_resp_valid),
    .io_in_resp_bits_rdata(dmem_proxy_io_in_resp_bits_rdata),
    .io_in_resp_bits_page_fault(dmem_proxy_io_in_resp_bits_page_fault),
    .io_in_resp_bits_access_fault(dmem_proxy_io_in_resp_bits_access_fault),
    .io_out_req_ready(dmem_proxy_io_out_req_ready),
    .io_out_req_valid(dmem_proxy_io_out_req_valid),
    .io_out_req_bits_addr(dmem_proxy_io_out_req_bits_addr),
    .io_out_req_bits_wdata(dmem_proxy_io_out_req_bits_wdata),
    .io_out_req_bits_wmask(dmem_proxy_io_out_req_bits_wmask),
    .io_out_req_bits_wen(dmem_proxy_io_out_req_bits_wen),
    .io_out_req_bits_len(dmem_proxy_io_out_req_bits_len),
    .io_out_req_bits_lrsc(dmem_proxy_io_out_req_bits_lrsc),
    .io_out_req_bits_amo(dmem_proxy_io_out_req_bits_amo),
    .io_out_resp_ready(dmem_proxy_io_out_resp_ready),
    .io_out_resp_valid(dmem_proxy_io_out_resp_valid),
    .io_out_resp_bits_rdata(dmem_proxy_io_out_resp_bits_rdata),
    .io_ptw_req_ready(dmem_proxy_io_ptw_req_ready),
    .io_ptw_req_valid(dmem_proxy_io_ptw_req_valid),
    .io_ptw_req_bits_addr(dmem_proxy_io_ptw_req_bits_addr),
    .io_ptw_resp_ready(dmem_proxy_io_ptw_resp_ready),
    .io_ptw_resp_valid(dmem_proxy_io_ptw_resp_valid),
    .io_ptw_resp_bits_rdata(dmem_proxy_io_ptw_resp_bits_rdata)
  );
  CachePortXBar1to2 c2_xbar ( // @[Core.scala 164:23]
    .clock(c2_xbar_clock),
    .reset(c2_xbar_reset),
    .io_in_req_ready(c2_xbar_io_in_req_ready),
    .io_in_req_valid(c2_xbar_io_in_req_valid),
    .io_in_req_bits_addr(c2_xbar_io_in_req_bits_addr),
    .io_in_req_bits_wdata(c2_xbar_io_in_req_bits_wdata),
    .io_in_req_bits_wmask(c2_xbar_io_in_req_bits_wmask),
    .io_in_req_bits_wen(c2_xbar_io_in_req_bits_wen),
    .io_in_req_bits_len(c2_xbar_io_in_req_bits_len),
    .io_in_req_bits_lrsc(c2_xbar_io_in_req_bits_lrsc),
    .io_in_req_bits_amo(c2_xbar_io_in_req_bits_amo),
    .io_in_resp_ready(c2_xbar_io_in_resp_ready),
    .io_in_resp_valid(c2_xbar_io_in_resp_valid),
    .io_in_resp_bits_rdata(c2_xbar_io_in_resp_bits_rdata),
    .io_out_0_req_ready(c2_xbar_io_out_0_req_ready),
    .io_out_0_req_valid(c2_xbar_io_out_0_req_valid),
    .io_out_0_req_bits_addr(c2_xbar_io_out_0_req_bits_addr),
    .io_out_0_req_bits_wdata(c2_xbar_io_out_0_req_bits_wdata),
    .io_out_0_req_bits_wmask(c2_xbar_io_out_0_req_bits_wmask),
    .io_out_0_req_bits_wen(c2_xbar_io_out_0_req_bits_wen),
    .io_out_0_req_bits_len(c2_xbar_io_out_0_req_bits_len),
    .io_out_0_req_bits_lrsc(c2_xbar_io_out_0_req_bits_lrsc),
    .io_out_0_req_bits_amo(c2_xbar_io_out_0_req_bits_amo),
    .io_out_0_resp_ready(c2_xbar_io_out_0_resp_ready),
    .io_out_0_resp_valid(c2_xbar_io_out_0_resp_valid),
    .io_out_0_resp_bits_rdata(c2_xbar_io_out_0_resp_bits_rdata),
    .io_out_1_req_ready(c2_xbar_io_out_1_req_ready),
    .io_out_1_req_valid(c2_xbar_io_out_1_req_valid),
    .io_out_1_req_bits_addr(c2_xbar_io_out_1_req_bits_addr),
    .io_out_1_req_bits_wdata(c2_xbar_io_out_1_req_bits_wdata),
    .io_out_1_req_bits_wmask(c2_xbar_io_out_1_req_bits_wmask),
    .io_out_1_req_bits_wen(c2_xbar_io_out_1_req_bits_wen),
    .io_out_1_req_bits_len(c2_xbar_io_out_1_req_bits_len),
    .io_out_1_resp_ready(c2_xbar_io_out_1_resp_ready),
    .io_out_1_resp_valid(c2_xbar_io_out_1_resp_valid),
    .io_out_1_resp_bits_rdata(c2_xbar_io_out_1_resp_bits_rdata),
    .io_to_1(c2_xbar_io_to_1)
  );
  PipelineReg_1 ex_wb ( // @[Core.scala 172:21]
    .clock(ex_wb_clock),
    .reset(ex_wb_reset),
    .io_in_uop_valid(ex_wb_io_in_uop_valid),
    .io_in_uop_rd_index(ex_wb_io_in_uop_rd_index),
    .io_in_uop_rd_wen(ex_wb_io_in_uop_rd_wen),
    .io_in_rd_data(ex_wb_io_in_rd_data),
    .io_out_uop_valid(ex_wb_io_out_uop_valid),
    .io_out_uop_rd_index(ex_wb_io_out_uop_rd_index),
    .io_out_uop_rd_wen(ex_wb_io_out_uop_rd_wen),
    .io_out_rd_data(ex_wb_io_out_rd_data)
  );
  assign io_imem_req_valid = imem_proxy_io_out_req_valid; // @[Core.scala 33:28]
  assign io_imem_req_bits_addr = imem_proxy_io_out_req_bits_addr; // @[Core.scala 33:28]
  assign io_imem_resp_ready = imem_proxy_io_out_resp_ready; // @[Core.scala 33:28]
  assign io_dmem_req_valid = c2_xbar_io_out_0_req_valid; // @[Core.scala 169:20]
  assign io_dmem_req_bits_addr = c2_xbar_io_out_0_req_bits_addr; // @[Core.scala 169:20]
  assign io_dmem_req_bits_wdata = c2_xbar_io_out_0_req_bits_wdata; // @[Core.scala 169:20]
  assign io_dmem_req_bits_wmask = c2_xbar_io_out_0_req_bits_wmask; // @[Core.scala 169:20]
  assign io_dmem_req_bits_wen = c2_xbar_io_out_0_req_bits_wen; // @[Core.scala 169:20]
  assign io_dmem_req_bits_len = c2_xbar_io_out_0_req_bits_len; // @[Core.scala 169:20]
  assign io_dmem_req_bits_lrsc = c2_xbar_io_out_0_req_bits_lrsc; // @[Core.scala 169:20]
  assign io_dmem_req_bits_amo = c2_xbar_io_out_0_req_bits_amo; // @[Core.scala 169:20]
  assign io_dmem_resp_ready = c2_xbar_io_out_0_resp_ready; // @[Core.scala 169:20]
  assign io_iptw_req_valid = imem_proxy_io_ptw_req_valid; // @[Core.scala 34:28]
  assign io_iptw_req_bits_addr = imem_proxy_io_ptw_req_bits_addr; // @[Core.scala 34:28]
  assign io_iptw_resp_ready = imem_proxy_io_ptw_resp_ready; // @[Core.scala 34:28]
  assign io_dptw_req_valid = dmem_proxy_io_ptw_req_valid; // @[Core.scala 166:20]
  assign io_dptw_req_bits_addr = dmem_proxy_io_ptw_req_bits_addr; // @[Core.scala 166:20]
  assign io_dptw_resp_ready = dmem_proxy_io_ptw_resp_ready; // @[Core.scala 166:20]
  assign io_uncache_req_valid = c2_xbar_io_out_1_req_valid; // @[Core.scala 170:20]
  assign io_uncache_req_bits_addr = c2_xbar_io_out_1_req_bits_addr; // @[Core.scala 170:20]
  assign io_uncache_req_bits_wdata = c2_xbar_io_out_1_req_bits_wdata; // @[Core.scala 170:20]
  assign io_uncache_req_bits_wmask = c2_xbar_io_out_1_req_bits_wmask; // @[Core.scala 170:20]
  assign io_uncache_req_bits_wen = c2_xbar_io_out_1_req_bits_wen; // @[Core.scala 170:20]
  assign io_uncache_req_bits_len = c2_xbar_io_out_1_req_bits_len; // @[Core.scala 170:20]
  assign io_uncache_resp_ready = c2_xbar_io_out_1_resp_ready; // @[Core.scala 170:20]
  assign io_fence_i = csr_io_fence_i; // @[Core.scala 136:23]
  assign ifu_clock = clock;
  assign ifu_reset = reset;
  assign ifu_io_jmp_packet_valid = alu_jmp_packet_valid | sys_jmp_packet_valid; // @[Core.scala 43:55]
  assign ifu_io_jmp_packet_target = sys_jmp_packet_valid ? sys_jmp_packet_target : alu_jmp_packet_target; // @[Core.scala 44:37]
  assign ifu_io_jmp_packet_bp_update = id_ex_io_out_uop_valid & alu_io_uop_jmp_op != 2'h0; // @[Core.scala 96:54]
  assign ifu_io_jmp_packet_bp_taken = _alu_jmp_packet_target_T_5 ? alu_io_cmp_out : alu_io_uop_jmp_op[1]; // @[Core.scala 97:34]
  assign ifu_io_jmp_packet_bp_pc = id_ex_io_out_uop_pc; // @[Core.scala 41:28 98:28]
  assign ifu_io_imem_req_ready = imem_proxy_io_in_req_ready; // @[Core.scala 32:28]
  assign ifu_io_imem_resp_valid = imem_proxy_io_in_resp_valid; // @[Core.scala 32:28]
  assign ifu_io_imem_resp_bits_rdata = imem_proxy_io_in_resp_bits_rdata; // @[Core.scala 32:28]
  assign ifu_io_imem_resp_bits_page_fault = imem_proxy_io_in_resp_bits_page_fault; // @[Core.scala 32:28]
  assign ifu_io_imem_resp_bits_access_fault = imem_proxy_io_in_resp_bits_access_fault; // @[Core.scala 32:28]
  assign ifu_io_stall_b = instr_buffer_io_enq_ready; // @[Core.scala 55:29]
  assign imem_proxy_clock = clock;
  assign imem_proxy_reset = reset;
  assign imem_proxy_io_prv = csr_io_prv; // @[Core.scala 128:23 19:24]
  assign imem_proxy_io_sv39_en = csr_io_sv39_en; // @[Core.scala 129:23 20:24]
  assign imem_proxy_io_satp_asid = csr_io_satp_asid; // @[Core.scala 130:23 21:24]
  assign imem_proxy_io_satp_ppn = csr_io_satp_ppn; // @[Core.scala 131:23 22:24]
  assign imem_proxy_io_sfence_vma = csr_io_sfence_vma; // @[Core.scala 132:23 23:24]
  assign imem_proxy_io_in_req_valid = ifu_io_imem_req_valid; // @[Core.scala 32:28]
  assign imem_proxy_io_in_req_bits_addr = ifu_io_imem_req_bits_addr; // @[Core.scala 32:28]
  assign imem_proxy_io_in_resp_ready = ifu_io_imem_resp_ready; // @[Core.scala 32:28]
  assign imem_proxy_io_out_req_ready = io_imem_req_ready; // @[Core.scala 33:28]
  assign imem_proxy_io_out_resp_valid = io_imem_resp_valid; // @[Core.scala 33:28]
  assign imem_proxy_io_out_resp_bits_rdata = io_imem_resp_bits_rdata; // @[Core.scala 33:28]
  assign imem_proxy_io_ptw_req_ready = io_iptw_req_ready; // @[Core.scala 34:28]
  assign imem_proxy_io_ptw_resp_valid = io_iptw_resp_valid; // @[Core.scala 34:28]
  assign imem_proxy_io_ptw_resp_bits_rdata = io_iptw_resp_bits_rdata; // @[Core.scala 34:28]
  assign instr_buffer_clock = clock;
  assign instr_buffer_reset = reset;
  assign instr_buffer_io_enq_valid = ifu_io_out_valid; // @[Core.scala 57:29]
  assign instr_buffer_io_enq_bits_pc = ifu_io_out_pc; // @[Core.scala 56:29]
  assign instr_buffer_io_enq_bits_instr = ifu_io_out_instr; // @[Core.scala 56:29]
  assign instr_buffer_io_enq_bits_page_fault = ifu_io_out_page_fault; // @[Core.scala 56:29]
  assign instr_buffer_io_enq_bits_access_fault = ifu_io_out_access_fault; // @[Core.scala 56:29]
  assign instr_buffer_io_enq_bits_bp_npc = ifu_io_out_bp_npc; // @[Core.scala 56:29]
  assign instr_buffer_io_deq_ready = lsu_io_ready & mdu_io_ready; // @[Core.scala 255:27]
  assign instr_buffer_io_flush = alu_jmp_packet_valid | sys_jmp_packet_valid; // @[Core.scala 256:35]
  assign decode_io_in_pc = instr_buffer_io_deq_bits_pc; // @[Core.scala 64:22]
  assign decode_io_in_instr = instr_buffer_io_deq_bits_instr; // @[Core.scala 64:22]
  assign decode_io_in_valid = instr_buffer_io_deq_ready & instr_buffer_io_deq_valid; // @[Decoupled.scala 51:35]
  assign decode_io_in_page_fault = instr_buffer_io_deq_bits_page_fault; // @[Core.scala 64:22]
  assign decode_io_in_access_fault = instr_buffer_io_deq_bits_access_fault; // @[Core.scala 64:22]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_rs1_index = decode_io_out_rs1_index; // @[Core.scala 68:19]
  assign rf_io_rs2_index = decode_io_out_rs2_index; // @[Core.scala 69:19]
  assign rf_io_rd_index = ex_wb_io_out_uop_rd_index; // @[Core.scala 197:18]
  assign rf_io_rd_data = ex_wb_io_out_rd_data; // @[Core.scala 198:18]
  assign rf_io_rd_wen = ex_wb_io_out_uop_valid & ex_wb_io_out_uop_rd_wen; // @[Core.scala 196:38]
  assign id_ex_clock = clock;
  assign id_ex_reset = reset;
  assign id_ex_io_in_uop_valid = decode_io_out_valid; // @[Core.scala 75:32]
  assign id_ex_io_in_uop_exc = decode_io_out_exc; // @[Core.scala 75:32]
  assign id_ex_io_in_uop_pc = decode_io_out_pc; // @[Core.scala 75:32]
  assign id_ex_io_in_uop_npc = decode_io_out_npc; // @[Core.scala 75:32]
  assign id_ex_io_in_uop_instr = decode_io_out_instr; // @[Core.scala 75:32]
  assign id_ex_io_in_uop_fu = decode_io_out_fu; // @[Core.scala 75:32]
  assign id_ex_io_in_uop_alu_op = decode_io_out_alu_op; // @[Core.scala 75:32]
  assign id_ex_io_in_uop_jmp_op = decode_io_out_jmp_op; // @[Core.scala 75:32]
  assign id_ex_io_in_uop_mdu_op = decode_io_out_mdu_op; // @[Core.scala 75:32]
  assign id_ex_io_in_uop_lsu_op = decode_io_out_lsu_op; // @[Core.scala 75:32]
  assign id_ex_io_in_uop_mem_len = decode_io_out_mem_len; // @[Core.scala 75:32]
  assign id_ex_io_in_uop_csr_op = decode_io_out_csr_op; // @[Core.scala 75:32]
  assign id_ex_io_in_uop_sys_op = decode_io_out_sys_op; // @[Core.scala 75:32]
  assign id_ex_io_in_uop_rd_index = decode_io_out_rd_index; // @[Core.scala 75:32]
  assign id_ex_io_in_uop_rd_wen = decode_io_out_rd_wen; // @[Core.scala 75:32]
  assign id_ex_io_in_uop_imm = decode_io_out_imm; // @[Core.scala 75:32]
  assign id_ex_io_in_uop_dw = decode_io_out_dw; // @[Core.scala 75:32]
  assign id_ex_io_in_rs1_data = _GEN_0[63:0]; // @[Core.scala 71:33]
  assign id_ex_io_in_rs2_data = _GEN_1[63:0]; // @[Core.scala 72:33]
  assign id_ex_io_in_rs2_data_from_rf = _T_14 ? ex_wb_io_in_rd_data : rf_io_rs2_data; // @[Core.scala 247:5 248:25 250:25]
  assign id_ex_io_in_bp_npc = instr_buffer_io_deq_bits_bp_npc; // @[Core.scala 79:32]
  assign id_ex_io_en = lsu_io_ready & mdu_io_ready; // @[Core.scala 255:27]
  assign id_ex_io_flush = alu_jmp_packet_valid | sys_jmp_packet_valid; // @[Core.scala 256:35]
  assign alu_io_uop_alu_op = id_ex_io_out_uop_alu_op; // @[Core.scala 86:14]
  assign alu_io_uop_jmp_op = id_ex_io_out_uop_jmp_op; // @[Core.scala 86:14]
  assign alu_io_uop_dw = id_ex_io_out_uop_dw; // @[Core.scala 86:14]
  assign alu_io_in1 = id_ex_io_out_rs1_data; // @[Core.scala 87:14]
  assign alu_io_in2 = id_ex_io_out_rs2_data; // @[Core.scala 88:14]
  assign lsu_clock = clock;
  assign lsu_reset = reset;
  assign lsu_io_uop_lsu_op = id_ex_io_out_uop_lsu_op; // @[Core.scala 109:19]
  assign lsu_io_uop_mem_len = id_ex_io_out_uop_mem_len; // @[Core.scala 109:19]
  assign lsu_io_is_mem = id_ex_io_out_uop_fu == 3'h3 & id_ex_io_out_uop_valid; // @[Core.scala 102:58]
  assign lsu_io_is_store = ~id_ex_io_out_uop_lsu_op[4] & id_ex_io_out_uop_lsu_op[0]; // @[Constant.scala 82:45]
  assign lsu_io_is_amo = id_ex_io_out_uop_lsu_op[4]; // @[Constant.scala 81:33]
  assign lsu_io_addr = id_ex_io_out_uop_jmp_op[1] ? id_ex_io_out_uop_npc : alu_io_out; // @[Core.scala 100:23]
  assign lsu_io_wdata = id_ex_io_out_rs2_data_from_rf; // @[Core.scala 114:19]
  assign lsu_io_dmem_req_ready = dmem_proxy_io_in_req_ready; // @[Core.scala 165:20]
  assign lsu_io_dmem_resp_valid = dmem_proxy_io_in_resp_valid; // @[Core.scala 165:20]
  assign lsu_io_dmem_resp_bits_rdata = dmem_proxy_io_in_resp_bits_rdata; // @[Core.scala 165:20]
  assign lsu_io_dmem_resp_bits_page_fault = dmem_proxy_io_in_resp_bits_page_fault; // @[Core.scala 165:20]
  assign lsu_io_dmem_resp_bits_access_fault = dmem_proxy_io_in_resp_bits_access_fault; // @[Core.scala 165:20]
  assign mdu_clock = clock;
  assign mdu_reset = reset;
  assign mdu_io_uop_valid = id_ex_io_out_uop_valid; // @[Core.scala 117:17]
  assign mdu_io_uop_mdu_op = id_ex_io_out_uop_mdu_op; // @[Core.scala 117:17]
  assign mdu_io_uop_dw = id_ex_io_out_uop_dw; // @[Core.scala 117:17]
  assign mdu_io_is_mdu = id_ex_io_out_uop_fu == 3'h2 & id_ex_io_out_uop_valid; // @[Core.scala 103:58]
  assign mdu_io_in1 = id_ex_io_out_rs1_data; // @[Core.scala 119:17]
  assign mdu_io_in2 = id_ex_io_out_rs2_data_from_rf; // @[Core.scala 120:17]
  assign csr_clock = clock;
  assign csr_reset = reset;
  assign csr_io_uop_valid = id_ex_io_out_uop_valid; // @[Core.scala 123:23]
  assign csr_io_uop_exc = id_ex_io_out_uop_exc; // @[Core.scala 123:23]
  assign csr_io_uop_pc = id_ex_io_out_uop_pc; // @[Core.scala 123:23]
  assign csr_io_uop_npc = id_ex_io_out_uop_npc; // @[Core.scala 123:23]
  assign csr_io_uop_fu = id_ex_io_out_uop_fu; // @[Core.scala 123:23]
  assign csr_io_uop_sys_op = id_ex_io_out_uop_sys_op; // @[Core.scala 123:23]
  assign csr_io_rw_addr = id_ex_io_out_uop_instr[31:20]; // @[Core.scala 124:48]
  assign csr_io_rw_cmd = id_ex_io_out_uop_csr_op; // @[Core.scala 125:23]
  assign csr_io_rw_wdata = id_ex_io_out_rs1_data; // @[Core.scala 126:23]
  assign csr_io_lsu_addr = lsu_io_addr; // @[Core.scala 133:23]
  assign csr_io_lsu_exc_code = lsu_io_exc_code; // @[Core.scala 134:23]
  assign csr_io_interrupt_mtip = io_intr_mtip; // @[Core.scala 135:23]
  assign csr_io_interrupt_msip = io_intr_msip; // @[Core.scala 135:23]
  assign csr_io_interrupt_meip = io_intr_meip; // @[Core.scala 135:23]
  assign csr_io_interrupt_seip = io_intr_seip; // @[Core.scala 135:23]
  assign csr_io_commit = ex_wb_io_out_uop_valid; // @[Core.scala 262:17]
  assign dmem_proxy_clock = clock;
  assign dmem_proxy_reset = reset;
  assign dmem_proxy_io_prv = csr_io_mprv ? csr_io_mpp : prv; // @[Core.scala 146:34]
  assign dmem_proxy_io_sv39_en = csr_io_sv39_en; // @[Core.scala 129:23 20:24]
  assign dmem_proxy_io_satp_asid = csr_io_satp_asid; // @[Core.scala 130:23 21:24]
  assign dmem_proxy_io_satp_ppn = csr_io_satp_ppn; // @[Core.scala 131:23 22:24]
  assign dmem_proxy_io_sfence_vma = csr_io_sfence_vma; // @[Core.scala 132:23 23:24]
  assign dmem_proxy_io_in_req_valid = lsu_io_dmem_req_valid; // @[Core.scala 165:20]
  assign dmem_proxy_io_in_req_bits_addr = lsu_io_dmem_req_bits_addr; // @[Core.scala 165:20]
  assign dmem_proxy_io_in_req_bits_wdata = lsu_io_dmem_req_bits_wdata; // @[Core.scala 165:20]
  assign dmem_proxy_io_in_req_bits_wmask = lsu_io_dmem_req_bits_wmask; // @[Core.scala 165:20]
  assign dmem_proxy_io_in_req_bits_wen = lsu_io_dmem_req_bits_wen; // @[Core.scala 165:20]
  assign dmem_proxy_io_in_req_bits_len = lsu_io_dmem_req_bits_len; // @[Core.scala 165:20]
  assign dmem_proxy_io_in_req_bits_lrsc = lsu_io_dmem_req_bits_lrsc; // @[Core.scala 165:20]
  assign dmem_proxy_io_in_req_bits_amo = lsu_io_dmem_req_bits_amo; // @[Core.scala 165:20]
  assign dmem_proxy_io_in_resp_ready = lsu_io_dmem_resp_ready; // @[Core.scala 165:20]
  assign dmem_proxy_io_out_req_ready = c2_xbar_io_in_req_ready; // @[Core.scala 167:20]
  assign dmem_proxy_io_out_resp_valid = c2_xbar_io_in_resp_valid; // @[Core.scala 167:20]
  assign dmem_proxy_io_out_resp_bits_rdata = c2_xbar_io_in_resp_bits_rdata; // @[Core.scala 167:20]
  assign dmem_proxy_io_ptw_req_ready = io_dptw_req_ready; // @[Core.scala 166:20]
  assign dmem_proxy_io_ptw_resp_valid = io_dptw_resp_valid; // @[Core.scala 166:20]
  assign dmem_proxy_io_ptw_resp_bits_rdata = io_dptw_resp_bits_rdata; // @[Core.scala 166:20]
  assign c2_xbar_clock = clock;
  assign c2_xbar_reset = reset;
  assign c2_xbar_io_in_req_valid = dmem_proxy_io_out_req_valid; // @[Core.scala 167:20]
  assign c2_xbar_io_in_req_bits_addr = dmem_proxy_io_out_req_bits_addr; // @[Core.scala 167:20]
  assign c2_xbar_io_in_req_bits_wdata = dmem_proxy_io_out_req_bits_wdata; // @[Core.scala 167:20]
  assign c2_xbar_io_in_req_bits_wmask = dmem_proxy_io_out_req_bits_wmask; // @[Core.scala 167:20]
  assign c2_xbar_io_in_req_bits_wen = dmem_proxy_io_out_req_bits_wen; // @[Core.scala 167:20]
  assign c2_xbar_io_in_req_bits_len = dmem_proxy_io_out_req_bits_len; // @[Core.scala 167:20]
  assign c2_xbar_io_in_req_bits_lrsc = dmem_proxy_io_out_req_bits_lrsc; // @[Core.scala 167:20]
  assign c2_xbar_io_in_req_bits_amo = dmem_proxy_io_out_req_bits_amo; // @[Core.scala 167:20]
  assign c2_xbar_io_in_resp_ready = dmem_proxy_io_out_resp_ready; // @[Core.scala 167:20]
  assign c2_xbar_io_out_0_req_ready = io_dmem_req_ready; // @[Core.scala 169:20]
  assign c2_xbar_io_out_0_resp_valid = io_dmem_resp_valid; // @[Core.scala 169:20]
  assign c2_xbar_io_out_0_resp_bits_rdata = io_dmem_resp_bits_rdata; // @[Core.scala 169:20]
  assign c2_xbar_io_out_1_req_ready = io_uncache_req_ready; // @[Core.scala 170:20]
  assign c2_xbar_io_out_1_resp_valid = io_uncache_resp_valid; // @[Core.scala 170:20]
  assign c2_xbar_io_out_1_resp_bits_rdata = io_uncache_resp_bits_rdata; // @[Core.scala 170:20]
  assign c2_xbar_io_to_1 = ~dmem_proxy_io_out_req_bits_addr[31]; // @[Core.scala 168:23]
  assign ex_wb_clock = clock;
  assign ex_wb_reset = reset;
  assign ex_wb_io_in_uop_valid = _ex_wb_io_in_uop_valid_T_13 & ~csr_io_is_int; // @[Core.scala 179:5]
  assign ex_wb_io_in_uop_rd_index = id_ex_io_out_uop_rd_index; // @[Core.scala 173:19]
  assign ex_wb_io_in_uop_rd_wen = id_ex_io_out_uop_rd_wen; // @[Core.scala 173:19]
  assign ex_wb_io_in_rd_data = 3'h4 == id_ex_io_out_uop_fu ? csr_io_rw_rdata : _ex_wb_io_in_rd_data_T_3; // @[Mux.scala 81:58]
endmodule
module RRArbiter(
  input         clock,
  input         io_in_0_valid,
  input  [38:0] io_in_0_bits_addr,
  input  [63:0] io_in_0_bits_wdata,
  input  [7:0]  io_in_0_bits_wmask,
  input         io_in_0_bits_wen,
  input  [1:0]  io_in_0_bits_len,
  input         io_in_0_bits_lrsc,
  input  [4:0]  io_in_0_bits_amo,
  input         io_in_1_valid,
  input  [38:0] io_in_1_bits_addr,
  input         io_in_2_valid,
  input  [38:0] io_in_2_bits_addr,
  input         io_out_ready,
  output        io_out_valid,
  output [38:0] io_out_bits_addr,
  output [63:0] io_out_bits_wdata,
  output [7:0]  io_out_bits_wmask,
  output        io_out_bits_wen,
  output [1:0]  io_out_bits_len,
  output        io_out_bits_lrsc,
  output [4:0]  io_out_bits_amo,
  output [1:0]  io_chosen
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  _GEN_1 = 2'h1 == io_chosen ? io_in_1_valid : io_in_0_valid; // @[Arbiter.scala 55:{16,16}]
  wire [38:0] _GEN_4 = 2'h1 == io_chosen ? io_in_1_bits_addr : io_in_0_bits_addr; // @[Arbiter.scala 56:{15,15}]
  wire [63:0] _GEN_7 = 2'h1 == io_chosen ? 64'h0 : io_in_0_bits_wdata; // @[Arbiter.scala 56:{15,15}]
  wire [7:0] _GEN_10 = 2'h1 == io_chosen ? 8'h0 : io_in_0_bits_wmask; // @[Arbiter.scala 56:{15,15}]
  wire  _GEN_13 = 2'h1 == io_chosen ? 1'h0 : io_in_0_bits_wen; // @[Arbiter.scala 56:{15,15}]
  wire [1:0] _GEN_16 = 2'h1 == io_chosen ? 2'h0 : io_in_0_bits_len; // @[Arbiter.scala 56:{15,15}]
  wire  _GEN_19 = 2'h1 == io_chosen ? 1'h0 : io_in_0_bits_lrsc; // @[Arbiter.scala 56:{15,15}]
  wire [4:0] _GEN_22 = 2'h1 == io_chosen ? 5'h0 : io_in_0_bits_amo; // @[Arbiter.scala 56:{15,15}]
  wire  _ctrl_validMask_grantMask_lastGrant_T = io_out_ready & io_out_valid; // @[Decoupled.scala 51:35]
  reg [1:0] lastGrant; // @[Reg.scala 19:16]
  wire  grantMask_1 = 2'h1 > lastGrant; // @[Arbiter.scala 81:49]
  wire  grantMask_2 = 2'h2 > lastGrant; // @[Arbiter.scala 81:49]
  wire  validMask_1 = io_in_1_valid & grantMask_1; // @[Arbiter.scala 82:76]
  wire  validMask_2 = io_in_2_valid & grantMask_2; // @[Arbiter.scala 82:76]
  wire [1:0] _GEN_25 = io_in_1_valid ? 2'h1 : 2'h2; // @[Arbiter.scala 91:{26,35} 89:41]
  wire [1:0] _GEN_26 = io_in_0_valid ? 2'h0 : _GEN_25; // @[Arbiter.scala 91:{26,35}]
  wire [1:0] _GEN_27 = validMask_2 ? 2'h2 : _GEN_26; // @[Arbiter.scala 93:{24,33}]
  assign io_out_valid = 2'h2 == io_chosen ? io_in_2_valid : _GEN_1; // @[Arbiter.scala 55:{16,16}]
  assign io_out_bits_addr = 2'h2 == io_chosen ? io_in_2_bits_addr : _GEN_4; // @[Arbiter.scala 56:{15,15}]
  assign io_out_bits_wdata = 2'h2 == io_chosen ? 64'h0 : _GEN_7; // @[Arbiter.scala 56:{15,15}]
  assign io_out_bits_wmask = 2'h2 == io_chosen ? 8'h0 : _GEN_10; // @[Arbiter.scala 56:{15,15}]
  assign io_out_bits_wen = 2'h2 == io_chosen ? 1'h0 : _GEN_13; // @[Arbiter.scala 56:{15,15}]
  assign io_out_bits_len = 2'h2 == io_chosen ? 2'h0 : _GEN_16; // @[Arbiter.scala 56:{15,15}]
  assign io_out_bits_lrsc = 2'h2 == io_chosen ? 1'h0 : _GEN_19; // @[Arbiter.scala 56:{15,15}]
  assign io_out_bits_amo = 2'h2 == io_chosen ? 5'h0 : _GEN_22; // @[Arbiter.scala 56:{15,15}]
  assign io_chosen = validMask_1 ? 2'h1 : _GEN_27; // @[Arbiter.scala 93:{24,33}]
  always @(posedge clock) begin
    if (_ctrl_validMask_grantMask_lastGrant_T) begin // @[Reg.scala 20:18]
      lastGrant <= io_chosen; // @[Reg.scala 20:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lastGrant = _RAND_0[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_3(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [1:0] io_enq_bits,
  input        io_deq_ready,
  output       io_deq_valid,
  output [1:0] io_deq_bits
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] ram [0:3]; // @[Decoupled.scala 273:95]
  wire  ram_io_deq_bits_MPORT_en; // @[Decoupled.scala 273:95]
  wire [1:0] ram_io_deq_bits_MPORT_addr; // @[Decoupled.scala 273:95]
  wire [1:0] ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_MPORT_data; // @[Decoupled.scala 273:95]
  wire [1:0] ram_MPORT_addr; // @[Decoupled.scala 273:95]
  wire  ram_MPORT_mask; // @[Decoupled.scala 273:95]
  wire  ram_MPORT_en; // @[Decoupled.scala 273:95]
  reg [1:0] enq_ptr_value; // @[Counter.scala 61:40]
  reg [1:0] deq_ptr_value; // @[Counter.scala 61:40]
  reg  maybe_full; // @[Decoupled.scala 276:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 277:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 278:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 279:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  wire [1:0] _value_T_1 = enq_ptr_value + 2'h1; // @[Counter.scala 77:24]
  wire [1:0] _value_T_3 = deq_ptr_value + 2'h1; // @[Counter.scala 77:24]
  assign ram_io_deq_bits_MPORT_en = 1'h1;
  assign ram_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 273:95]
  assign ram_MPORT_data = io_enq_bits;
  assign ram_MPORT_addr = enq_ptr_value;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 303:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 302:19]
  assign io_deq_bits = ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 310:17]
  always @(posedge clock) begin
    if (ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[Decoupled.scala 273:95]
    end
    if (reset) begin // @[Counter.scala 61:40]
      enq_ptr_value <= 2'h0; // @[Counter.scala 61:40]
    end else if (do_enq) begin // @[Decoupled.scala 286:16]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Counter.scala 61:40]
      deq_ptr_value <= 2'h0; // @[Counter.scala 61:40]
    end else if (do_deq) begin // @[Decoupled.scala 290:16]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 77:15]
    end
    if (reset) begin // @[Decoupled.scala 276:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 276:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 293:27]
      maybe_full <= do_enq; // @[Decoupled.scala 294:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram[initvar] = _RAND_0[1:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enq_ptr_value = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  deq_ptr_value = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CachePortXBarNto1(
  input         clock,
  input         reset,
  output        io_in_0_req_ready,
  input         io_in_0_req_valid,
  input  [38:0] io_in_0_req_bits_addr,
  input  [63:0] io_in_0_req_bits_wdata,
  input  [7:0]  io_in_0_req_bits_wmask,
  input         io_in_0_req_bits_wen,
  input  [1:0]  io_in_0_req_bits_len,
  input         io_in_0_req_bits_lrsc,
  input  [4:0]  io_in_0_req_bits_amo,
  input         io_in_0_resp_ready,
  output        io_in_0_resp_valid,
  output [63:0] io_in_0_resp_bits_rdata,
  output        io_in_1_req_ready,
  input         io_in_1_req_valid,
  input  [38:0] io_in_1_req_bits_addr,
  input         io_in_1_resp_ready,
  output        io_in_1_resp_valid,
  output [63:0] io_in_1_resp_bits_rdata,
  output        io_in_2_req_ready,
  input         io_in_2_req_valid,
  input  [38:0] io_in_2_req_bits_addr,
  input         io_in_2_resp_ready,
  output        io_in_2_resp_valid,
  output [63:0] io_in_2_resp_bits_rdata,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [38:0] io_out_req_bits_addr,
  output [63:0] io_out_req_bits_wdata,
  output [7:0]  io_out_req_bits_wmask,
  output        io_out_req_bits_wen,
  output [1:0]  io_out_req_bits_len,
  output        io_out_req_bits_lrsc,
  output [4:0]  io_out_req_bits_amo,
  output        io_out_resp_ready,
  input         io_out_resp_valid,
  input  [63:0] io_out_resp_bits_rdata
);
  wire  arbiter_clock; // @[Bus.scala 47:23]
  wire  arbiter_io_in_0_valid; // @[Bus.scala 47:23]
  wire [38:0] arbiter_io_in_0_bits_addr; // @[Bus.scala 47:23]
  wire [63:0] arbiter_io_in_0_bits_wdata; // @[Bus.scala 47:23]
  wire [7:0] arbiter_io_in_0_bits_wmask; // @[Bus.scala 47:23]
  wire  arbiter_io_in_0_bits_wen; // @[Bus.scala 47:23]
  wire [1:0] arbiter_io_in_0_bits_len; // @[Bus.scala 47:23]
  wire  arbiter_io_in_0_bits_lrsc; // @[Bus.scala 47:23]
  wire [4:0] arbiter_io_in_0_bits_amo; // @[Bus.scala 47:23]
  wire  arbiter_io_in_1_valid; // @[Bus.scala 47:23]
  wire [38:0] arbiter_io_in_1_bits_addr; // @[Bus.scala 47:23]
  wire  arbiter_io_in_2_valid; // @[Bus.scala 47:23]
  wire [38:0] arbiter_io_in_2_bits_addr; // @[Bus.scala 47:23]
  wire  arbiter_io_out_ready; // @[Bus.scala 47:23]
  wire  arbiter_io_out_valid; // @[Bus.scala 47:23]
  wire [38:0] arbiter_io_out_bits_addr; // @[Bus.scala 47:23]
  wire [63:0] arbiter_io_out_bits_wdata; // @[Bus.scala 47:23]
  wire [7:0] arbiter_io_out_bits_wmask; // @[Bus.scala 47:23]
  wire  arbiter_io_out_bits_wen; // @[Bus.scala 47:23]
  wire [1:0] arbiter_io_out_bits_len; // @[Bus.scala 47:23]
  wire  arbiter_io_out_bits_lrsc; // @[Bus.scala 47:23]
  wire [4:0] arbiter_io_out_bits_amo; // @[Bus.scala 47:23]
  wire [1:0] arbiter_io_chosen; // @[Bus.scala 47:23]
  wire  id_queue_clock; // @[Bus.scala 54:24]
  wire  id_queue_reset; // @[Bus.scala 54:24]
  wire  id_queue_io_enq_ready; // @[Bus.scala 54:24]
  wire  id_queue_io_enq_valid; // @[Bus.scala 54:24]
  wire [1:0] id_queue_io_enq_bits; // @[Bus.scala 54:24]
  wire  id_queue_io_deq_ready; // @[Bus.scala 54:24]
  wire  id_queue_io_deq_valid; // @[Bus.scala 54:24]
  wire [1:0] id_queue_io_deq_bits; // @[Bus.scala 54:24]
  wire  _GEN_0 = id_queue_io_deq_valid & id_queue_io_deq_bits == 2'h0 & io_in_0_resp_ready; // @[Bus.scala 75:25 78:67 79:27]
  wire  _GEN_2 = id_queue_io_deq_valid & id_queue_io_deq_bits == 2'h1 ? io_in_1_resp_ready : _GEN_0; // @[Bus.scala 78:67 79:27]
  RRArbiter arbiter ( // @[Bus.scala 47:23]
    .clock(arbiter_clock),
    .io_in_0_valid(arbiter_io_in_0_valid),
    .io_in_0_bits_addr(arbiter_io_in_0_bits_addr),
    .io_in_0_bits_wdata(arbiter_io_in_0_bits_wdata),
    .io_in_0_bits_wmask(arbiter_io_in_0_bits_wmask),
    .io_in_0_bits_wen(arbiter_io_in_0_bits_wen),
    .io_in_0_bits_len(arbiter_io_in_0_bits_len),
    .io_in_0_bits_lrsc(arbiter_io_in_0_bits_lrsc),
    .io_in_0_bits_amo(arbiter_io_in_0_bits_amo),
    .io_in_1_valid(arbiter_io_in_1_valid),
    .io_in_1_bits_addr(arbiter_io_in_1_bits_addr),
    .io_in_2_valid(arbiter_io_in_2_valid),
    .io_in_2_bits_addr(arbiter_io_in_2_bits_addr),
    .io_out_ready(arbiter_io_out_ready),
    .io_out_valid(arbiter_io_out_valid),
    .io_out_bits_addr(arbiter_io_out_bits_addr),
    .io_out_bits_wdata(arbiter_io_out_bits_wdata),
    .io_out_bits_wmask(arbiter_io_out_bits_wmask),
    .io_out_bits_wen(arbiter_io_out_bits_wen),
    .io_out_bits_len(arbiter_io_out_bits_len),
    .io_out_bits_lrsc(arbiter_io_out_bits_lrsc),
    .io_out_bits_amo(arbiter_io_out_bits_amo),
    .io_chosen(arbiter_io_chosen)
  );
  Queue_3 id_queue ( // @[Bus.scala 54:24]
    .clock(id_queue_clock),
    .reset(id_queue_reset),
    .io_enq_ready(id_queue_io_enq_ready),
    .io_enq_valid(id_queue_io_enq_valid),
    .io_enq_bits(id_queue_io_enq_bits),
    .io_deq_ready(id_queue_io_deq_ready),
    .io_deq_valid(id_queue_io_deq_valid),
    .io_deq_bits(id_queue_io_deq_bits)
  );
  assign io_in_0_req_ready = arbiter_io_chosen == 2'h0 & io_out_req_ready & id_queue_io_enq_ready; // @[Bus.scala 61:75]
  assign io_in_0_resp_valid = id_queue_io_deq_valid & id_queue_io_deq_bits == 2'h0 & io_out_resp_valid; // @[Bus.scala 74:25 78:67 80:27]
  assign io_in_0_resp_bits_rdata = io_out_resp_bits_rdata; // @[Bus.scala 73:25]
  assign io_in_1_req_ready = arbiter_io_chosen == 2'h1 & io_out_req_ready & id_queue_io_enq_ready; // @[Bus.scala 61:75]
  assign io_in_1_resp_valid = id_queue_io_deq_valid & id_queue_io_deq_bits == 2'h1 & io_out_resp_valid; // @[Bus.scala 74:25 78:67 80:27]
  assign io_in_1_resp_bits_rdata = io_out_resp_bits_rdata; // @[Bus.scala 73:25]
  assign io_in_2_req_ready = arbiter_io_chosen == 2'h2 & io_out_req_ready & id_queue_io_enq_ready; // @[Bus.scala 61:75]
  assign io_in_2_resp_valid = id_queue_io_deq_valid & id_queue_io_deq_bits == 2'h2 & io_out_resp_valid; // @[Bus.scala 74:25 78:67 80:27]
  assign io_in_2_resp_bits_rdata = io_out_resp_bits_rdata; // @[Bus.scala 73:25]
  assign io_out_req_valid = arbiter_io_out_valid; // @[Bus.scala 66:15]
  assign io_out_req_bits_addr = arbiter_io_out_bits_addr; // @[Bus.scala 65:15]
  assign io_out_req_bits_wdata = arbiter_io_out_bits_wdata; // @[Bus.scala 65:15]
  assign io_out_req_bits_wmask = arbiter_io_out_bits_wmask; // @[Bus.scala 65:15]
  assign io_out_req_bits_wen = arbiter_io_out_bits_wen; // @[Bus.scala 65:15]
  assign io_out_req_bits_len = arbiter_io_out_bits_len; // @[Bus.scala 65:15]
  assign io_out_req_bits_lrsc = arbiter_io_out_bits_lrsc; // @[Bus.scala 65:15]
  assign io_out_req_bits_amo = arbiter_io_out_bits_amo; // @[Bus.scala 65:15]
  assign io_out_resp_ready = id_queue_io_deq_valid & id_queue_io_deq_bits == 2'h2 ? io_in_2_resp_ready : _GEN_2; // @[Bus.scala 78:67 79:27]
  assign arbiter_clock = clock;
  assign arbiter_io_in_0_valid = io_in_0_req_valid; // @[Bus.scala 50:22]
  assign arbiter_io_in_0_bits_addr = io_in_0_req_bits_addr; // @[Bus.scala 50:22]
  assign arbiter_io_in_0_bits_wdata = io_in_0_req_bits_wdata; // @[Bus.scala 50:22]
  assign arbiter_io_in_0_bits_wmask = io_in_0_req_bits_wmask; // @[Bus.scala 50:22]
  assign arbiter_io_in_0_bits_wen = io_in_0_req_bits_wen; // @[Bus.scala 50:22]
  assign arbiter_io_in_0_bits_len = io_in_0_req_bits_len; // @[Bus.scala 50:22]
  assign arbiter_io_in_0_bits_lrsc = io_in_0_req_bits_lrsc; // @[Bus.scala 50:22]
  assign arbiter_io_in_0_bits_amo = io_in_0_req_bits_amo; // @[Bus.scala 50:22]
  assign arbiter_io_in_1_valid = io_in_1_req_valid; // @[Bus.scala 50:22]
  assign arbiter_io_in_1_bits_addr = io_in_1_req_bits_addr; // @[Bus.scala 50:22]
  assign arbiter_io_in_2_valid = io_in_2_req_valid; // @[Bus.scala 50:22]
  assign arbiter_io_in_2_bits_addr = io_in_2_req_bits_addr; // @[Bus.scala 50:22]
  assign arbiter_io_out_ready = io_out_req_ready; // @[Bus.scala 67:15]
  assign id_queue_clock = clock;
  assign id_queue_reset = reset;
  assign id_queue_io_enq_valid = io_out_req_ready & io_out_req_valid; // @[Decoupled.scala 51:35]
  assign id_queue_io_enq_bits = arbiter_io_chosen; // @[Bus.scala 56:25]
  assign id_queue_io_deq_ready = io_out_resp_ready & io_out_resp_valid; // @[Decoupled.scala 51:35]
endmodule
module SoCImp(
  input          clock,
  input          reset,
  input          auto_out_a_ready,
  output         auto_out_a_valid,
  output [2:0]   auto_out_a_bits_opcode,
  output [2:0]   auto_out_a_bits_param,
  output [2:0]   auto_out_a_bits_size,
  output [3:0]   auto_out_a_bits_source,
  output [31:0]  auto_out_a_bits_address,
  output [31:0]  auto_out_a_bits_mask,
  output [255:0] auto_out_a_bits_data,
  output         auto_out_b_ready,
  input          auto_out_b_valid,
  input  [2:0]   auto_out_b_bits_size,
  input  [3:0]   auto_out_b_bits_source,
  input  [31:0]  auto_out_b_bits_address,
  input          auto_out_c_ready,
  output         auto_out_c_valid,
  output [2:0]   auto_out_c_bits_opcode,
  output [2:0]   auto_out_c_bits_param,
  output [2:0]   auto_out_c_bits_size,
  output [3:0]   auto_out_c_bits_source,
  output [31:0]  auto_out_c_bits_address,
  output [255:0] auto_out_c_bits_data,
  output         auto_out_d_ready,
  input          auto_out_d_valid,
  input  [2:0]   auto_out_d_bits_opcode,
  input  [2:0]   auto_out_d_bits_size,
  input  [3:0]   auto_out_d_bits_source,
  input  [5:0]   auto_out_d_bits_sink,
  input  [255:0] auto_out_d_bits_data,
  input          auto_out_e_ready,
  output         auto_out_e_valid,
  output [5:0]   auto_out_e_bits_sink,
  input          io_intr_mtip,
  input          io_intr_msip,
  input          io_intr_meip,
  input          io_intr_seip
);
  wire  icache_clock; // @[SoC.scala 27:27]
  wire  icache_reset; // @[SoC.scala 27:27]
  wire  icache_auto_out_a_ready; // @[SoC.scala 27:27]
  wire  icache_auto_out_a_valid; // @[SoC.scala 27:27]
  wire [1:0] icache_auto_out_a_bits_source; // @[SoC.scala 27:27]
  wire [31:0] icache_auto_out_a_bits_address; // @[SoC.scala 27:27]
  wire  icache_auto_out_d_ready; // @[SoC.scala 27:27]
  wire  icache_auto_out_d_valid; // @[SoC.scala 27:27]
  wire [255:0] icache_auto_out_d_bits_data; // @[SoC.scala 27:27]
  wire  icache_io_cache_req_ready; // @[SoC.scala 27:27]
  wire  icache_io_cache_req_valid; // @[SoC.scala 27:27]
  wire [38:0] icache_io_cache_req_bits_addr; // @[SoC.scala 27:27]
  wire  icache_io_cache_resp_ready; // @[SoC.scala 27:27]
  wire  icache_io_cache_resp_valid; // @[SoC.scala 27:27]
  wire [63:0] icache_io_cache_resp_bits_rdata; // @[SoC.scala 27:27]
  wire  icache_io_fence_i; // @[SoC.scala 27:27]
  wire  dcache_clock; // @[SoC.scala 28:27]
  wire  dcache_reset; // @[SoC.scala 28:27]
  wire  dcache_auto_out_a_ready; // @[SoC.scala 28:27]
  wire  dcache_auto_out_a_valid; // @[SoC.scala 28:27]
  wire [1:0] dcache_auto_out_a_bits_source; // @[SoC.scala 28:27]
  wire [31:0] dcache_auto_out_a_bits_address; // @[SoC.scala 28:27]
  wire  dcache_auto_out_b_ready; // @[SoC.scala 28:27]
  wire  dcache_auto_out_b_valid; // @[SoC.scala 28:27]
  wire [2:0] dcache_auto_out_b_bits_size; // @[SoC.scala 28:27]
  wire [1:0] dcache_auto_out_b_bits_source; // @[SoC.scala 28:27]
  wire [31:0] dcache_auto_out_b_bits_address; // @[SoC.scala 28:27]
  wire  dcache_auto_out_c_ready; // @[SoC.scala 28:27]
  wire  dcache_auto_out_c_valid; // @[SoC.scala 28:27]
  wire [2:0] dcache_auto_out_c_bits_opcode; // @[SoC.scala 28:27]
  wire [2:0] dcache_auto_out_c_bits_param; // @[SoC.scala 28:27]
  wire [2:0] dcache_auto_out_c_bits_size; // @[SoC.scala 28:27]
  wire [1:0] dcache_auto_out_c_bits_source; // @[SoC.scala 28:27]
  wire [31:0] dcache_auto_out_c_bits_address; // @[SoC.scala 28:27]
  wire [255:0] dcache_auto_out_c_bits_data; // @[SoC.scala 28:27]
  wire  dcache_auto_out_d_ready; // @[SoC.scala 28:27]
  wire  dcache_auto_out_d_valid; // @[SoC.scala 28:27]
  wire [5:0] dcache_auto_out_d_bits_sink; // @[SoC.scala 28:27]
  wire [255:0] dcache_auto_out_d_bits_data; // @[SoC.scala 28:27]
  wire  dcache_auto_out_e_ready; // @[SoC.scala 28:27]
  wire  dcache_auto_out_e_valid; // @[SoC.scala 28:27]
  wire [5:0] dcache_auto_out_e_bits_sink; // @[SoC.scala 28:27]
  wire  dcache_io_cache_req_ready; // @[SoC.scala 28:27]
  wire  dcache_io_cache_req_valid; // @[SoC.scala 28:27]
  wire [38:0] dcache_io_cache_req_bits_addr; // @[SoC.scala 28:27]
  wire [63:0] dcache_io_cache_req_bits_wdata; // @[SoC.scala 28:27]
  wire [7:0] dcache_io_cache_req_bits_wmask; // @[SoC.scala 28:27]
  wire  dcache_io_cache_req_bits_wen; // @[SoC.scala 28:27]
  wire [1:0] dcache_io_cache_req_bits_len; // @[SoC.scala 28:27]
  wire  dcache_io_cache_req_bits_lrsc; // @[SoC.scala 28:27]
  wire [4:0] dcache_io_cache_req_bits_amo; // @[SoC.scala 28:27]
  wire  dcache_io_cache_resp_ready; // @[SoC.scala 28:27]
  wire  dcache_io_cache_resp_valid; // @[SoC.scala 28:27]
  wire [63:0] dcache_io_cache_resp_bits_rdata; // @[SoC.scala 28:27]
  wire  uncache_clock; // @[SoC.scala 29:27]
  wire  uncache_reset; // @[SoC.scala 29:27]
  wire  uncache_auto_out_a_ready; // @[SoC.scala 29:27]
  wire  uncache_auto_out_a_valid; // @[SoC.scala 29:27]
  wire [2:0] uncache_auto_out_a_bits_opcode; // @[SoC.scala 29:27]
  wire [2:0] uncache_auto_out_a_bits_size; // @[SoC.scala 29:27]
  wire [1:0] uncache_auto_out_a_bits_source; // @[SoC.scala 29:27]
  wire [31:0] uncache_auto_out_a_bits_address; // @[SoC.scala 29:27]
  wire [7:0] uncache_auto_out_a_bits_mask; // @[SoC.scala 29:27]
  wire [63:0] uncache_auto_out_a_bits_data; // @[SoC.scala 29:27]
  wire  uncache_auto_out_d_ready; // @[SoC.scala 29:27]
  wire  uncache_auto_out_d_valid; // @[SoC.scala 29:27]
  wire [63:0] uncache_auto_out_d_bits_data; // @[SoC.scala 29:27]
  wire  uncache_io_in_req_ready; // @[SoC.scala 29:27]
  wire  uncache_io_in_req_valid; // @[SoC.scala 29:27]
  wire [38:0] uncache_io_in_req_bits_addr; // @[SoC.scala 29:27]
  wire [63:0] uncache_io_in_req_bits_wdata; // @[SoC.scala 29:27]
  wire [7:0] uncache_io_in_req_bits_wmask; // @[SoC.scala 29:27]
  wire  uncache_io_in_req_bits_wen; // @[SoC.scala 29:27]
  wire [1:0] uncache_io_in_req_bits_len; // @[SoC.scala 29:27]
  wire  uncache_io_in_resp_ready; // @[SoC.scala 29:27]
  wire  uncache_io_in_resp_valid; // @[SoC.scala 29:27]
  wire [63:0] uncache_io_in_resp_bits_rdata; // @[SoC.scala 29:27]
  wire  xbar_clock; // @[SoC.scala 30:27]
  wire  xbar_reset; // @[SoC.scala 30:27]
  wire  xbar_auto_in_2_a_ready; // @[SoC.scala 30:27]
  wire  xbar_auto_in_2_a_valid; // @[SoC.scala 30:27]
  wire [1:0] xbar_auto_in_2_a_bits_source; // @[SoC.scala 30:27]
  wire [31:0] xbar_auto_in_2_a_bits_address; // @[SoC.scala 30:27]
  wire  xbar_auto_in_2_b_ready; // @[SoC.scala 30:27]
  wire  xbar_auto_in_2_b_valid; // @[SoC.scala 30:27]
  wire [2:0] xbar_auto_in_2_b_bits_size; // @[SoC.scala 30:27]
  wire [1:0] xbar_auto_in_2_b_bits_source; // @[SoC.scala 30:27]
  wire [31:0] xbar_auto_in_2_b_bits_address; // @[SoC.scala 30:27]
  wire  xbar_auto_in_2_c_ready; // @[SoC.scala 30:27]
  wire  xbar_auto_in_2_c_valid; // @[SoC.scala 30:27]
  wire [2:0] xbar_auto_in_2_c_bits_opcode; // @[SoC.scala 30:27]
  wire [2:0] xbar_auto_in_2_c_bits_param; // @[SoC.scala 30:27]
  wire [2:0] xbar_auto_in_2_c_bits_size; // @[SoC.scala 30:27]
  wire [1:0] xbar_auto_in_2_c_bits_source; // @[SoC.scala 30:27]
  wire [31:0] xbar_auto_in_2_c_bits_address; // @[SoC.scala 30:27]
  wire [255:0] xbar_auto_in_2_c_bits_data; // @[SoC.scala 30:27]
  wire  xbar_auto_in_2_d_ready; // @[SoC.scala 30:27]
  wire  xbar_auto_in_2_d_valid; // @[SoC.scala 30:27]
  wire [5:0] xbar_auto_in_2_d_bits_sink; // @[SoC.scala 30:27]
  wire [255:0] xbar_auto_in_2_d_bits_data; // @[SoC.scala 30:27]
  wire  xbar_auto_in_2_e_ready; // @[SoC.scala 30:27]
  wire  xbar_auto_in_2_e_valid; // @[SoC.scala 30:27]
  wire [5:0] xbar_auto_in_2_e_bits_sink; // @[SoC.scala 30:27]
  wire  xbar_auto_in_1_a_ready; // @[SoC.scala 30:27]
  wire  xbar_auto_in_1_a_valid; // @[SoC.scala 30:27]
  wire [2:0] xbar_auto_in_1_a_bits_opcode; // @[SoC.scala 30:27]
  wire [2:0] xbar_auto_in_1_a_bits_size; // @[SoC.scala 30:27]
  wire [1:0] xbar_auto_in_1_a_bits_source; // @[SoC.scala 30:27]
  wire [31:0] xbar_auto_in_1_a_bits_address; // @[SoC.scala 30:27]
  wire [31:0] xbar_auto_in_1_a_bits_mask; // @[SoC.scala 30:27]
  wire [255:0] xbar_auto_in_1_a_bits_data; // @[SoC.scala 30:27]
  wire  xbar_auto_in_1_d_ready; // @[SoC.scala 30:27]
  wire  xbar_auto_in_1_d_valid; // @[SoC.scala 30:27]
  wire [2:0] xbar_auto_in_1_d_bits_opcode; // @[SoC.scala 30:27]
  wire [2:0] xbar_auto_in_1_d_bits_size; // @[SoC.scala 30:27]
  wire [1:0] xbar_auto_in_1_d_bits_source; // @[SoC.scala 30:27]
  wire [255:0] xbar_auto_in_1_d_bits_data; // @[SoC.scala 30:27]
  wire  xbar_auto_in_0_a_ready; // @[SoC.scala 30:27]
  wire  xbar_auto_in_0_a_valid; // @[SoC.scala 30:27]
  wire [1:0] xbar_auto_in_0_a_bits_source; // @[SoC.scala 30:27]
  wire [31:0] xbar_auto_in_0_a_bits_address; // @[SoC.scala 30:27]
  wire  xbar_auto_in_0_d_ready; // @[SoC.scala 30:27]
  wire  xbar_auto_in_0_d_valid; // @[SoC.scala 30:27]
  wire [255:0] xbar_auto_in_0_d_bits_data; // @[SoC.scala 30:27]
  wire  xbar_auto_out_a_ready; // @[SoC.scala 30:27]
  wire  xbar_auto_out_a_valid; // @[SoC.scala 30:27]
  wire [2:0] xbar_auto_out_a_bits_opcode; // @[SoC.scala 30:27]
  wire [2:0] xbar_auto_out_a_bits_param; // @[SoC.scala 30:27]
  wire [2:0] xbar_auto_out_a_bits_size; // @[SoC.scala 30:27]
  wire [3:0] xbar_auto_out_a_bits_source; // @[SoC.scala 30:27]
  wire [31:0] xbar_auto_out_a_bits_address; // @[SoC.scala 30:27]
  wire [31:0] xbar_auto_out_a_bits_mask; // @[SoC.scala 30:27]
  wire [255:0] xbar_auto_out_a_bits_data; // @[SoC.scala 30:27]
  wire  xbar_auto_out_b_ready; // @[SoC.scala 30:27]
  wire  xbar_auto_out_b_valid; // @[SoC.scala 30:27]
  wire [2:0] xbar_auto_out_b_bits_size; // @[SoC.scala 30:27]
  wire [3:0] xbar_auto_out_b_bits_source; // @[SoC.scala 30:27]
  wire [31:0] xbar_auto_out_b_bits_address; // @[SoC.scala 30:27]
  wire  xbar_auto_out_c_ready; // @[SoC.scala 30:27]
  wire  xbar_auto_out_c_valid; // @[SoC.scala 30:27]
  wire [2:0] xbar_auto_out_c_bits_opcode; // @[SoC.scala 30:27]
  wire [2:0] xbar_auto_out_c_bits_param; // @[SoC.scala 30:27]
  wire [2:0] xbar_auto_out_c_bits_size; // @[SoC.scala 30:27]
  wire [3:0] xbar_auto_out_c_bits_source; // @[SoC.scala 30:27]
  wire [31:0] xbar_auto_out_c_bits_address; // @[SoC.scala 30:27]
  wire [255:0] xbar_auto_out_c_bits_data; // @[SoC.scala 30:27]
  wire  xbar_auto_out_d_ready; // @[SoC.scala 30:27]
  wire  xbar_auto_out_d_valid; // @[SoC.scala 30:27]
  wire [2:0] xbar_auto_out_d_bits_opcode; // @[SoC.scala 30:27]
  wire [2:0] xbar_auto_out_d_bits_size; // @[SoC.scala 30:27]
  wire [3:0] xbar_auto_out_d_bits_source; // @[SoC.scala 30:27]
  wire [5:0] xbar_auto_out_d_bits_sink; // @[SoC.scala 30:27]
  wire [255:0] xbar_auto_out_d_bits_data; // @[SoC.scala 30:27]
  wire  xbar_auto_out_e_ready; // @[SoC.scala 30:27]
  wire  xbar_auto_out_e_valid; // @[SoC.scala 30:27]
  wire [5:0] xbar_auto_out_e_bits_sink; // @[SoC.scala 30:27]
  wire  widget_clock; // @[WidthWidget.scala 220:28]
  wire  widget_reset; // @[WidthWidget.scala 220:28]
  wire  widget_auto_in_a_ready; // @[WidthWidget.scala 220:28]
  wire  widget_auto_in_a_valid; // @[WidthWidget.scala 220:28]
  wire [2:0] widget_auto_in_a_bits_opcode; // @[WidthWidget.scala 220:28]
  wire [2:0] widget_auto_in_a_bits_size; // @[WidthWidget.scala 220:28]
  wire [1:0] widget_auto_in_a_bits_source; // @[WidthWidget.scala 220:28]
  wire [31:0] widget_auto_in_a_bits_address; // @[WidthWidget.scala 220:28]
  wire [7:0] widget_auto_in_a_bits_mask; // @[WidthWidget.scala 220:28]
  wire [63:0] widget_auto_in_a_bits_data; // @[WidthWidget.scala 220:28]
  wire  widget_auto_in_d_ready; // @[WidthWidget.scala 220:28]
  wire  widget_auto_in_d_valid; // @[WidthWidget.scala 220:28]
  wire [63:0] widget_auto_in_d_bits_data; // @[WidthWidget.scala 220:28]
  wire  widget_auto_out_a_ready; // @[WidthWidget.scala 220:28]
  wire  widget_auto_out_a_valid; // @[WidthWidget.scala 220:28]
  wire [2:0] widget_auto_out_a_bits_opcode; // @[WidthWidget.scala 220:28]
  wire [2:0] widget_auto_out_a_bits_size; // @[WidthWidget.scala 220:28]
  wire [1:0] widget_auto_out_a_bits_source; // @[WidthWidget.scala 220:28]
  wire [31:0] widget_auto_out_a_bits_address; // @[WidthWidget.scala 220:28]
  wire [31:0] widget_auto_out_a_bits_mask; // @[WidthWidget.scala 220:28]
  wire [255:0] widget_auto_out_a_bits_data; // @[WidthWidget.scala 220:28]
  wire  widget_auto_out_d_ready; // @[WidthWidget.scala 220:28]
  wire  widget_auto_out_d_valid; // @[WidthWidget.scala 220:28]
  wire [2:0] widget_auto_out_d_bits_opcode; // @[WidthWidget.scala 220:28]
  wire [2:0] widget_auto_out_d_bits_size; // @[WidthWidget.scala 220:28]
  wire [1:0] widget_auto_out_d_bits_source; // @[WidthWidget.scala 220:28]
  wire [255:0] widget_auto_out_d_bits_data; // @[WidthWidget.scala 220:28]
  wire  core_clock; // @[SoC.scala 40:22]
  wire  core_reset; // @[SoC.scala 40:22]
  wire  core_io_imem_req_ready; // @[SoC.scala 40:22]
  wire  core_io_imem_req_valid; // @[SoC.scala 40:22]
  wire [38:0] core_io_imem_req_bits_addr; // @[SoC.scala 40:22]
  wire  core_io_imem_resp_ready; // @[SoC.scala 40:22]
  wire  core_io_imem_resp_valid; // @[SoC.scala 40:22]
  wire [63:0] core_io_imem_resp_bits_rdata; // @[SoC.scala 40:22]
  wire  core_io_dmem_req_ready; // @[SoC.scala 40:22]
  wire  core_io_dmem_req_valid; // @[SoC.scala 40:22]
  wire [38:0] core_io_dmem_req_bits_addr; // @[SoC.scala 40:22]
  wire [63:0] core_io_dmem_req_bits_wdata; // @[SoC.scala 40:22]
  wire [7:0] core_io_dmem_req_bits_wmask; // @[SoC.scala 40:22]
  wire  core_io_dmem_req_bits_wen; // @[SoC.scala 40:22]
  wire [1:0] core_io_dmem_req_bits_len; // @[SoC.scala 40:22]
  wire  core_io_dmem_req_bits_lrsc; // @[SoC.scala 40:22]
  wire [4:0] core_io_dmem_req_bits_amo; // @[SoC.scala 40:22]
  wire  core_io_dmem_resp_ready; // @[SoC.scala 40:22]
  wire  core_io_dmem_resp_valid; // @[SoC.scala 40:22]
  wire [63:0] core_io_dmem_resp_bits_rdata; // @[SoC.scala 40:22]
  wire  core_io_iptw_req_ready; // @[SoC.scala 40:22]
  wire  core_io_iptw_req_valid; // @[SoC.scala 40:22]
  wire [38:0] core_io_iptw_req_bits_addr; // @[SoC.scala 40:22]
  wire  core_io_iptw_resp_ready; // @[SoC.scala 40:22]
  wire  core_io_iptw_resp_valid; // @[SoC.scala 40:22]
  wire [63:0] core_io_iptw_resp_bits_rdata; // @[SoC.scala 40:22]
  wire  core_io_dptw_req_ready; // @[SoC.scala 40:22]
  wire  core_io_dptw_req_valid; // @[SoC.scala 40:22]
  wire [38:0] core_io_dptw_req_bits_addr; // @[SoC.scala 40:22]
  wire  core_io_dptw_resp_ready; // @[SoC.scala 40:22]
  wire  core_io_dptw_resp_valid; // @[SoC.scala 40:22]
  wire [63:0] core_io_dptw_resp_bits_rdata; // @[SoC.scala 40:22]
  wire  core_io_uncache_req_ready; // @[SoC.scala 40:22]
  wire  core_io_uncache_req_valid; // @[SoC.scala 40:22]
  wire [38:0] core_io_uncache_req_bits_addr; // @[SoC.scala 40:22]
  wire [63:0] core_io_uncache_req_bits_wdata; // @[SoC.scala 40:22]
  wire [7:0] core_io_uncache_req_bits_wmask; // @[SoC.scala 40:22]
  wire  core_io_uncache_req_bits_wen; // @[SoC.scala 40:22]
  wire [1:0] core_io_uncache_req_bits_len; // @[SoC.scala 40:22]
  wire  core_io_uncache_resp_ready; // @[SoC.scala 40:22]
  wire  core_io_uncache_resp_valid; // @[SoC.scala 40:22]
  wire [63:0] core_io_uncache_resp_bits_rdata; // @[SoC.scala 40:22]
  wire  core_io_fence_i; // @[SoC.scala 40:22]
  wire  core_io_intr_mtip; // @[SoC.scala 40:22]
  wire  core_io_intr_msip; // @[SoC.scala 40:22]
  wire  core_io_intr_meip; // @[SoC.scala 40:22]
  wire  core_io_intr_seip; // @[SoC.scala 40:22]
  wire  xbar_1_clock; // @[SoC.scala 50:22]
  wire  xbar_1_reset; // @[SoC.scala 50:22]
  wire  xbar_1_io_in_0_req_ready; // @[SoC.scala 50:22]
  wire  xbar_1_io_in_0_req_valid; // @[SoC.scala 50:22]
  wire [38:0] xbar_1_io_in_0_req_bits_addr; // @[SoC.scala 50:22]
  wire [63:0] xbar_1_io_in_0_req_bits_wdata; // @[SoC.scala 50:22]
  wire [7:0] xbar_1_io_in_0_req_bits_wmask; // @[SoC.scala 50:22]
  wire  xbar_1_io_in_0_req_bits_wen; // @[SoC.scala 50:22]
  wire [1:0] xbar_1_io_in_0_req_bits_len; // @[SoC.scala 50:22]
  wire  xbar_1_io_in_0_req_bits_lrsc; // @[SoC.scala 50:22]
  wire [4:0] xbar_1_io_in_0_req_bits_amo; // @[SoC.scala 50:22]
  wire  xbar_1_io_in_0_resp_ready; // @[SoC.scala 50:22]
  wire  xbar_1_io_in_0_resp_valid; // @[SoC.scala 50:22]
  wire [63:0] xbar_1_io_in_0_resp_bits_rdata; // @[SoC.scala 50:22]
  wire  xbar_1_io_in_1_req_ready; // @[SoC.scala 50:22]
  wire  xbar_1_io_in_1_req_valid; // @[SoC.scala 50:22]
  wire [38:0] xbar_1_io_in_1_req_bits_addr; // @[SoC.scala 50:22]
  wire  xbar_1_io_in_1_resp_ready; // @[SoC.scala 50:22]
  wire  xbar_1_io_in_1_resp_valid; // @[SoC.scala 50:22]
  wire [63:0] xbar_1_io_in_1_resp_bits_rdata; // @[SoC.scala 50:22]
  wire  xbar_1_io_in_2_req_ready; // @[SoC.scala 50:22]
  wire  xbar_1_io_in_2_req_valid; // @[SoC.scala 50:22]
  wire [38:0] xbar_1_io_in_2_req_bits_addr; // @[SoC.scala 50:22]
  wire  xbar_1_io_in_2_resp_ready; // @[SoC.scala 50:22]
  wire  xbar_1_io_in_2_resp_valid; // @[SoC.scala 50:22]
  wire [63:0] xbar_1_io_in_2_resp_bits_rdata; // @[SoC.scala 50:22]
  wire  xbar_1_io_out_req_ready; // @[SoC.scala 50:22]
  wire  xbar_1_io_out_req_valid; // @[SoC.scala 50:22]
  wire [38:0] xbar_1_io_out_req_bits_addr; // @[SoC.scala 50:22]
  wire [63:0] xbar_1_io_out_req_bits_wdata; // @[SoC.scala 50:22]
  wire [7:0] xbar_1_io_out_req_bits_wmask; // @[SoC.scala 50:22]
  wire  xbar_1_io_out_req_bits_wen; // @[SoC.scala 50:22]
  wire [1:0] xbar_1_io_out_req_bits_len; // @[SoC.scala 50:22]
  wire  xbar_1_io_out_req_bits_lrsc; // @[SoC.scala 50:22]
  wire [4:0] xbar_1_io_out_req_bits_amo; // @[SoC.scala 50:22]
  wire  xbar_1_io_out_resp_ready; // @[SoC.scala 50:22]
  wire  xbar_1_io_out_resp_valid; // @[SoC.scala 50:22]
  wire [63:0] xbar_1_io_out_resp_bits_rdata; // @[SoC.scala 50:22]
  ICache icache ( // @[SoC.scala 27:27]
    .clock(icache_clock),
    .reset(icache_reset),
    .auto_out_a_ready(icache_auto_out_a_ready),
    .auto_out_a_valid(icache_auto_out_a_valid),
    .auto_out_a_bits_source(icache_auto_out_a_bits_source),
    .auto_out_a_bits_address(icache_auto_out_a_bits_address),
    .auto_out_d_ready(icache_auto_out_d_ready),
    .auto_out_d_valid(icache_auto_out_d_valid),
    .auto_out_d_bits_data(icache_auto_out_d_bits_data),
    .io_cache_req_ready(icache_io_cache_req_ready),
    .io_cache_req_valid(icache_io_cache_req_valid),
    .io_cache_req_bits_addr(icache_io_cache_req_bits_addr),
    .io_cache_resp_ready(icache_io_cache_resp_ready),
    .io_cache_resp_valid(icache_io_cache_resp_valid),
    .io_cache_resp_bits_rdata(icache_io_cache_resp_bits_rdata),
    .io_fence_i(icache_io_fence_i)
  );
  DCache dcache ( // @[SoC.scala 28:27]
    .clock(dcache_clock),
    .reset(dcache_reset),
    .auto_out_a_ready(dcache_auto_out_a_ready),
    .auto_out_a_valid(dcache_auto_out_a_valid),
    .auto_out_a_bits_source(dcache_auto_out_a_bits_source),
    .auto_out_a_bits_address(dcache_auto_out_a_bits_address),
    .auto_out_b_ready(dcache_auto_out_b_ready),
    .auto_out_b_valid(dcache_auto_out_b_valid),
    .auto_out_b_bits_size(dcache_auto_out_b_bits_size),
    .auto_out_b_bits_source(dcache_auto_out_b_bits_source),
    .auto_out_b_bits_address(dcache_auto_out_b_bits_address),
    .auto_out_c_ready(dcache_auto_out_c_ready),
    .auto_out_c_valid(dcache_auto_out_c_valid),
    .auto_out_c_bits_opcode(dcache_auto_out_c_bits_opcode),
    .auto_out_c_bits_param(dcache_auto_out_c_bits_param),
    .auto_out_c_bits_size(dcache_auto_out_c_bits_size),
    .auto_out_c_bits_source(dcache_auto_out_c_bits_source),
    .auto_out_c_bits_address(dcache_auto_out_c_bits_address),
    .auto_out_c_bits_data(dcache_auto_out_c_bits_data),
    .auto_out_d_ready(dcache_auto_out_d_ready),
    .auto_out_d_valid(dcache_auto_out_d_valid),
    .auto_out_d_bits_sink(dcache_auto_out_d_bits_sink),
    .auto_out_d_bits_data(dcache_auto_out_d_bits_data),
    .auto_out_e_ready(dcache_auto_out_e_ready),
    .auto_out_e_valid(dcache_auto_out_e_valid),
    .auto_out_e_bits_sink(dcache_auto_out_e_bits_sink),
    .io_cache_req_ready(dcache_io_cache_req_ready),
    .io_cache_req_valid(dcache_io_cache_req_valid),
    .io_cache_req_bits_addr(dcache_io_cache_req_bits_addr),
    .io_cache_req_bits_wdata(dcache_io_cache_req_bits_wdata),
    .io_cache_req_bits_wmask(dcache_io_cache_req_bits_wmask),
    .io_cache_req_bits_wen(dcache_io_cache_req_bits_wen),
    .io_cache_req_bits_len(dcache_io_cache_req_bits_len),
    .io_cache_req_bits_lrsc(dcache_io_cache_req_bits_lrsc),
    .io_cache_req_bits_amo(dcache_io_cache_req_bits_amo),
    .io_cache_resp_ready(dcache_io_cache_resp_ready),
    .io_cache_resp_valid(dcache_io_cache_resp_valid),
    .io_cache_resp_bits_rdata(dcache_io_cache_resp_bits_rdata)
  );
  Uncache uncache ( // @[SoC.scala 29:27]
    .clock(uncache_clock),
    .reset(uncache_reset),
    .auto_out_a_ready(uncache_auto_out_a_ready),
    .auto_out_a_valid(uncache_auto_out_a_valid),
    .auto_out_a_bits_opcode(uncache_auto_out_a_bits_opcode),
    .auto_out_a_bits_size(uncache_auto_out_a_bits_size),
    .auto_out_a_bits_source(uncache_auto_out_a_bits_source),
    .auto_out_a_bits_address(uncache_auto_out_a_bits_address),
    .auto_out_a_bits_mask(uncache_auto_out_a_bits_mask),
    .auto_out_a_bits_data(uncache_auto_out_a_bits_data),
    .auto_out_d_ready(uncache_auto_out_d_ready),
    .auto_out_d_valid(uncache_auto_out_d_valid),
    .auto_out_d_bits_data(uncache_auto_out_d_bits_data),
    .io_in_req_ready(uncache_io_in_req_ready),
    .io_in_req_valid(uncache_io_in_req_valid),
    .io_in_req_bits_addr(uncache_io_in_req_bits_addr),
    .io_in_req_bits_wdata(uncache_io_in_req_bits_wdata),
    .io_in_req_bits_wmask(uncache_io_in_req_bits_wmask),
    .io_in_req_bits_wen(uncache_io_in_req_bits_wen),
    .io_in_req_bits_len(uncache_io_in_req_bits_len),
    .io_in_resp_ready(uncache_io_in_resp_ready),
    .io_in_resp_valid(uncache_io_in_resp_valid),
    .io_in_resp_bits_rdata(uncache_io_in_resp_bits_rdata)
  );
  TLXbar xbar ( // @[SoC.scala 30:27]
    .clock(xbar_clock),
    .reset(xbar_reset),
    .auto_in_2_a_ready(xbar_auto_in_2_a_ready),
    .auto_in_2_a_valid(xbar_auto_in_2_a_valid),
    .auto_in_2_a_bits_source(xbar_auto_in_2_a_bits_source),
    .auto_in_2_a_bits_address(xbar_auto_in_2_a_bits_address),
    .auto_in_2_b_ready(xbar_auto_in_2_b_ready),
    .auto_in_2_b_valid(xbar_auto_in_2_b_valid),
    .auto_in_2_b_bits_size(xbar_auto_in_2_b_bits_size),
    .auto_in_2_b_bits_source(xbar_auto_in_2_b_bits_source),
    .auto_in_2_b_bits_address(xbar_auto_in_2_b_bits_address),
    .auto_in_2_c_ready(xbar_auto_in_2_c_ready),
    .auto_in_2_c_valid(xbar_auto_in_2_c_valid),
    .auto_in_2_c_bits_opcode(xbar_auto_in_2_c_bits_opcode),
    .auto_in_2_c_bits_param(xbar_auto_in_2_c_bits_param),
    .auto_in_2_c_bits_size(xbar_auto_in_2_c_bits_size),
    .auto_in_2_c_bits_source(xbar_auto_in_2_c_bits_source),
    .auto_in_2_c_bits_address(xbar_auto_in_2_c_bits_address),
    .auto_in_2_c_bits_data(xbar_auto_in_2_c_bits_data),
    .auto_in_2_d_ready(xbar_auto_in_2_d_ready),
    .auto_in_2_d_valid(xbar_auto_in_2_d_valid),
    .auto_in_2_d_bits_sink(xbar_auto_in_2_d_bits_sink),
    .auto_in_2_d_bits_data(xbar_auto_in_2_d_bits_data),
    .auto_in_2_e_ready(xbar_auto_in_2_e_ready),
    .auto_in_2_e_valid(xbar_auto_in_2_e_valid),
    .auto_in_2_e_bits_sink(xbar_auto_in_2_e_bits_sink),
    .auto_in_1_a_ready(xbar_auto_in_1_a_ready),
    .auto_in_1_a_valid(xbar_auto_in_1_a_valid),
    .auto_in_1_a_bits_opcode(xbar_auto_in_1_a_bits_opcode),
    .auto_in_1_a_bits_size(xbar_auto_in_1_a_bits_size),
    .auto_in_1_a_bits_source(xbar_auto_in_1_a_bits_source),
    .auto_in_1_a_bits_address(xbar_auto_in_1_a_bits_address),
    .auto_in_1_a_bits_mask(xbar_auto_in_1_a_bits_mask),
    .auto_in_1_a_bits_data(xbar_auto_in_1_a_bits_data),
    .auto_in_1_d_ready(xbar_auto_in_1_d_ready),
    .auto_in_1_d_valid(xbar_auto_in_1_d_valid),
    .auto_in_1_d_bits_opcode(xbar_auto_in_1_d_bits_opcode),
    .auto_in_1_d_bits_size(xbar_auto_in_1_d_bits_size),
    .auto_in_1_d_bits_source(xbar_auto_in_1_d_bits_source),
    .auto_in_1_d_bits_data(xbar_auto_in_1_d_bits_data),
    .auto_in_0_a_ready(xbar_auto_in_0_a_ready),
    .auto_in_0_a_valid(xbar_auto_in_0_a_valid),
    .auto_in_0_a_bits_source(xbar_auto_in_0_a_bits_source),
    .auto_in_0_a_bits_address(xbar_auto_in_0_a_bits_address),
    .auto_in_0_d_ready(xbar_auto_in_0_d_ready),
    .auto_in_0_d_valid(xbar_auto_in_0_d_valid),
    .auto_in_0_d_bits_data(xbar_auto_in_0_d_bits_data),
    .auto_out_a_ready(xbar_auto_out_a_ready),
    .auto_out_a_valid(xbar_auto_out_a_valid),
    .auto_out_a_bits_opcode(xbar_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(xbar_auto_out_a_bits_param),
    .auto_out_a_bits_size(xbar_auto_out_a_bits_size),
    .auto_out_a_bits_source(xbar_auto_out_a_bits_source),
    .auto_out_a_bits_address(xbar_auto_out_a_bits_address),
    .auto_out_a_bits_mask(xbar_auto_out_a_bits_mask),
    .auto_out_a_bits_data(xbar_auto_out_a_bits_data),
    .auto_out_b_ready(xbar_auto_out_b_ready),
    .auto_out_b_valid(xbar_auto_out_b_valid),
    .auto_out_b_bits_size(xbar_auto_out_b_bits_size),
    .auto_out_b_bits_source(xbar_auto_out_b_bits_source),
    .auto_out_b_bits_address(xbar_auto_out_b_bits_address),
    .auto_out_c_ready(xbar_auto_out_c_ready),
    .auto_out_c_valid(xbar_auto_out_c_valid),
    .auto_out_c_bits_opcode(xbar_auto_out_c_bits_opcode),
    .auto_out_c_bits_param(xbar_auto_out_c_bits_param),
    .auto_out_c_bits_size(xbar_auto_out_c_bits_size),
    .auto_out_c_bits_source(xbar_auto_out_c_bits_source),
    .auto_out_c_bits_address(xbar_auto_out_c_bits_address),
    .auto_out_c_bits_data(xbar_auto_out_c_bits_data),
    .auto_out_d_ready(xbar_auto_out_d_ready),
    .auto_out_d_valid(xbar_auto_out_d_valid),
    .auto_out_d_bits_opcode(xbar_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(xbar_auto_out_d_bits_size),
    .auto_out_d_bits_source(xbar_auto_out_d_bits_source),
    .auto_out_d_bits_sink(xbar_auto_out_d_bits_sink),
    .auto_out_d_bits_data(xbar_auto_out_d_bits_data),
    .auto_out_e_ready(xbar_auto_out_e_ready),
    .auto_out_e_valid(xbar_auto_out_e_valid),
    .auto_out_e_bits_sink(xbar_auto_out_e_bits_sink)
  );
  TLWidthWidget widget ( // @[WidthWidget.scala 220:28]
    .clock(widget_clock),
    .reset(widget_reset),
    .auto_in_a_ready(widget_auto_in_a_ready),
    .auto_in_a_valid(widget_auto_in_a_valid),
    .auto_in_a_bits_opcode(widget_auto_in_a_bits_opcode),
    .auto_in_a_bits_size(widget_auto_in_a_bits_size),
    .auto_in_a_bits_source(widget_auto_in_a_bits_source),
    .auto_in_a_bits_address(widget_auto_in_a_bits_address),
    .auto_in_a_bits_mask(widget_auto_in_a_bits_mask),
    .auto_in_a_bits_data(widget_auto_in_a_bits_data),
    .auto_in_d_ready(widget_auto_in_d_ready),
    .auto_in_d_valid(widget_auto_in_d_valid),
    .auto_in_d_bits_data(widget_auto_in_d_bits_data),
    .auto_out_a_ready(widget_auto_out_a_ready),
    .auto_out_a_valid(widget_auto_out_a_valid),
    .auto_out_a_bits_opcode(widget_auto_out_a_bits_opcode),
    .auto_out_a_bits_size(widget_auto_out_a_bits_size),
    .auto_out_a_bits_source(widget_auto_out_a_bits_source),
    .auto_out_a_bits_address(widget_auto_out_a_bits_address),
    .auto_out_a_bits_mask(widget_auto_out_a_bits_mask),
    .auto_out_a_bits_data(widget_auto_out_a_bits_data),
    .auto_out_d_ready(widget_auto_out_d_ready),
    .auto_out_d_valid(widget_auto_out_d_valid),
    .auto_out_d_bits_opcode(widget_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(widget_auto_out_d_bits_size),
    .auto_out_d_bits_source(widget_auto_out_d_bits_source),
    .auto_out_d_bits_data(widget_auto_out_d_bits_data)
  );
  Core core ( // @[SoC.scala 40:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_imem_req_ready(core_io_imem_req_ready),
    .io_imem_req_valid(core_io_imem_req_valid),
    .io_imem_req_bits_addr(core_io_imem_req_bits_addr),
    .io_imem_resp_ready(core_io_imem_resp_ready),
    .io_imem_resp_valid(core_io_imem_resp_valid),
    .io_imem_resp_bits_rdata(core_io_imem_resp_bits_rdata),
    .io_dmem_req_ready(core_io_dmem_req_ready),
    .io_dmem_req_valid(core_io_dmem_req_valid),
    .io_dmem_req_bits_addr(core_io_dmem_req_bits_addr),
    .io_dmem_req_bits_wdata(core_io_dmem_req_bits_wdata),
    .io_dmem_req_bits_wmask(core_io_dmem_req_bits_wmask),
    .io_dmem_req_bits_wen(core_io_dmem_req_bits_wen),
    .io_dmem_req_bits_len(core_io_dmem_req_bits_len),
    .io_dmem_req_bits_lrsc(core_io_dmem_req_bits_lrsc),
    .io_dmem_req_bits_amo(core_io_dmem_req_bits_amo),
    .io_dmem_resp_ready(core_io_dmem_resp_ready),
    .io_dmem_resp_valid(core_io_dmem_resp_valid),
    .io_dmem_resp_bits_rdata(core_io_dmem_resp_bits_rdata),
    .io_iptw_req_ready(core_io_iptw_req_ready),
    .io_iptw_req_valid(core_io_iptw_req_valid),
    .io_iptw_req_bits_addr(core_io_iptw_req_bits_addr),
    .io_iptw_resp_ready(core_io_iptw_resp_ready),
    .io_iptw_resp_valid(core_io_iptw_resp_valid),
    .io_iptw_resp_bits_rdata(core_io_iptw_resp_bits_rdata),
    .io_dptw_req_ready(core_io_dptw_req_ready),
    .io_dptw_req_valid(core_io_dptw_req_valid),
    .io_dptw_req_bits_addr(core_io_dptw_req_bits_addr),
    .io_dptw_resp_ready(core_io_dptw_resp_ready),
    .io_dptw_resp_valid(core_io_dptw_resp_valid),
    .io_dptw_resp_bits_rdata(core_io_dptw_resp_bits_rdata),
    .io_uncache_req_ready(core_io_uncache_req_ready),
    .io_uncache_req_valid(core_io_uncache_req_valid),
    .io_uncache_req_bits_addr(core_io_uncache_req_bits_addr),
    .io_uncache_req_bits_wdata(core_io_uncache_req_bits_wdata),
    .io_uncache_req_bits_wmask(core_io_uncache_req_bits_wmask),
    .io_uncache_req_bits_wen(core_io_uncache_req_bits_wen),
    .io_uncache_req_bits_len(core_io_uncache_req_bits_len),
    .io_uncache_resp_ready(core_io_uncache_resp_ready),
    .io_uncache_resp_valid(core_io_uncache_resp_valid),
    .io_uncache_resp_bits_rdata(core_io_uncache_resp_bits_rdata),
    .io_fence_i(core_io_fence_i),
    .io_intr_mtip(core_io_intr_mtip),
    .io_intr_msip(core_io_intr_msip),
    .io_intr_meip(core_io_intr_meip),
    .io_intr_seip(core_io_intr_seip)
  );
  CachePortXBarNto1 xbar_1 ( // @[SoC.scala 50:22]
    .clock(xbar_1_clock),
    .reset(xbar_1_reset),
    .io_in_0_req_ready(xbar_1_io_in_0_req_ready),
    .io_in_0_req_valid(xbar_1_io_in_0_req_valid),
    .io_in_0_req_bits_addr(xbar_1_io_in_0_req_bits_addr),
    .io_in_0_req_bits_wdata(xbar_1_io_in_0_req_bits_wdata),
    .io_in_0_req_bits_wmask(xbar_1_io_in_0_req_bits_wmask),
    .io_in_0_req_bits_wen(xbar_1_io_in_0_req_bits_wen),
    .io_in_0_req_bits_len(xbar_1_io_in_0_req_bits_len),
    .io_in_0_req_bits_lrsc(xbar_1_io_in_0_req_bits_lrsc),
    .io_in_0_req_bits_amo(xbar_1_io_in_0_req_bits_amo),
    .io_in_0_resp_ready(xbar_1_io_in_0_resp_ready),
    .io_in_0_resp_valid(xbar_1_io_in_0_resp_valid),
    .io_in_0_resp_bits_rdata(xbar_1_io_in_0_resp_bits_rdata),
    .io_in_1_req_ready(xbar_1_io_in_1_req_ready),
    .io_in_1_req_valid(xbar_1_io_in_1_req_valid),
    .io_in_1_req_bits_addr(xbar_1_io_in_1_req_bits_addr),
    .io_in_1_resp_ready(xbar_1_io_in_1_resp_ready),
    .io_in_1_resp_valid(xbar_1_io_in_1_resp_valid),
    .io_in_1_resp_bits_rdata(xbar_1_io_in_1_resp_bits_rdata),
    .io_in_2_req_ready(xbar_1_io_in_2_req_ready),
    .io_in_2_req_valid(xbar_1_io_in_2_req_valid),
    .io_in_2_req_bits_addr(xbar_1_io_in_2_req_bits_addr),
    .io_in_2_resp_ready(xbar_1_io_in_2_resp_ready),
    .io_in_2_resp_valid(xbar_1_io_in_2_resp_valid),
    .io_in_2_resp_bits_rdata(xbar_1_io_in_2_resp_bits_rdata),
    .io_out_req_ready(xbar_1_io_out_req_ready),
    .io_out_req_valid(xbar_1_io_out_req_valid),
    .io_out_req_bits_addr(xbar_1_io_out_req_bits_addr),
    .io_out_req_bits_wdata(xbar_1_io_out_req_bits_wdata),
    .io_out_req_bits_wmask(xbar_1_io_out_req_bits_wmask),
    .io_out_req_bits_wen(xbar_1_io_out_req_bits_wen),
    .io_out_req_bits_len(xbar_1_io_out_req_bits_len),
    .io_out_req_bits_lrsc(xbar_1_io_out_req_bits_lrsc),
    .io_out_req_bits_amo(xbar_1_io_out_req_bits_amo),
    .io_out_resp_ready(xbar_1_io_out_resp_ready),
    .io_out_resp_valid(xbar_1_io_out_resp_valid),
    .io_out_resp_bits_rdata(xbar_1_io_out_resp_bits_rdata)
  );
  assign auto_out_a_valid = xbar_auto_out_a_valid; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_out_a_bits_opcode = xbar_auto_out_a_bits_opcode; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_out_a_bits_param = xbar_auto_out_a_bits_param; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_out_a_bits_size = xbar_auto_out_a_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_out_a_bits_source = xbar_auto_out_a_bits_source; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_out_a_bits_address = xbar_auto_out_a_bits_address; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_out_a_bits_mask = xbar_auto_out_a_bits_mask; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_out_a_bits_data = xbar_auto_out_a_bits_data; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_out_b_ready = xbar_auto_out_b_ready; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_out_c_valid = xbar_auto_out_c_valid; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_out_c_bits_opcode = xbar_auto_out_c_bits_opcode; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_out_c_bits_param = xbar_auto_out_c_bits_param; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_out_c_bits_size = xbar_auto_out_c_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_out_c_bits_source = xbar_auto_out_c_bits_source; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_out_c_bits_address = xbar_auto_out_c_bits_address; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_out_c_bits_data = xbar_auto_out_c_bits_data; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_out_d_ready = xbar_auto_out_d_ready; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_out_e_valid = xbar_auto_out_e_valid; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign auto_out_e_bits_sink = xbar_auto_out_e_bits_sink; // @[Nodes.scala 1215:84 LazyModule.scala 353:16]
  assign icache_clock = clock;
  assign icache_reset = reset;
  assign icache_auto_out_a_ready = xbar_auto_in_0_a_ready; // @[LazyModule.scala 355:16]
  assign icache_auto_out_d_valid = xbar_auto_in_0_d_valid; // @[LazyModule.scala 355:16]
  assign icache_auto_out_d_bits_data = xbar_auto_in_0_d_bits_data; // @[LazyModule.scala 355:16]
  assign icache_io_cache_req_valid = core_io_imem_req_valid; // @[SoC.scala 46:30]
  assign icache_io_cache_req_bits_addr = core_io_imem_req_bits_addr; // @[SoC.scala 46:30]
  assign icache_io_cache_resp_ready = core_io_imem_resp_ready; // @[SoC.scala 46:30]
  assign icache_io_fence_i = core_io_fence_i; // @[SoC.scala 47:30]
  assign dcache_clock = clock;
  assign dcache_reset = reset;
  assign dcache_auto_out_a_ready = xbar_auto_in_2_a_ready; // @[LazyModule.scala 355:16]
  assign dcache_auto_out_b_valid = xbar_auto_in_2_b_valid; // @[LazyModule.scala 355:16]
  assign dcache_auto_out_b_bits_size = xbar_auto_in_2_b_bits_size; // @[LazyModule.scala 355:16]
  assign dcache_auto_out_b_bits_source = xbar_auto_in_2_b_bits_source; // @[LazyModule.scala 355:16]
  assign dcache_auto_out_b_bits_address = xbar_auto_in_2_b_bits_address; // @[LazyModule.scala 355:16]
  assign dcache_auto_out_c_ready = xbar_auto_in_2_c_ready; // @[LazyModule.scala 355:16]
  assign dcache_auto_out_d_valid = xbar_auto_in_2_d_valid; // @[LazyModule.scala 355:16]
  assign dcache_auto_out_d_bits_sink = xbar_auto_in_2_d_bits_sink; // @[LazyModule.scala 355:16]
  assign dcache_auto_out_d_bits_data = xbar_auto_in_2_d_bits_data; // @[LazyModule.scala 355:16]
  assign dcache_auto_out_e_ready = xbar_auto_in_2_e_ready; // @[LazyModule.scala 355:16]
  assign dcache_io_cache_req_valid = xbar_1_io_out_req_valid; // @[SoC.scala 54:28]
  assign dcache_io_cache_req_bits_addr = xbar_1_io_out_req_bits_addr; // @[SoC.scala 54:28]
  assign dcache_io_cache_req_bits_wdata = xbar_1_io_out_req_bits_wdata; // @[SoC.scala 54:28]
  assign dcache_io_cache_req_bits_wmask = xbar_1_io_out_req_bits_wmask; // @[SoC.scala 54:28]
  assign dcache_io_cache_req_bits_wen = xbar_1_io_out_req_bits_wen; // @[SoC.scala 54:28]
  assign dcache_io_cache_req_bits_len = xbar_1_io_out_req_bits_len; // @[SoC.scala 54:28]
  assign dcache_io_cache_req_bits_lrsc = xbar_1_io_out_req_bits_lrsc; // @[SoC.scala 54:28]
  assign dcache_io_cache_req_bits_amo = xbar_1_io_out_req_bits_amo; // @[SoC.scala 54:28]
  assign dcache_io_cache_resp_ready = xbar_1_io_out_resp_ready; // @[SoC.scala 54:28]
  assign uncache_clock = clock;
  assign uncache_reset = reset;
  assign uncache_auto_out_a_ready = widget_auto_in_a_ready; // @[LazyModule.scala 355:16]
  assign uncache_auto_out_d_valid = widget_auto_in_d_valid; // @[LazyModule.scala 355:16]
  assign uncache_auto_out_d_bits_data = widget_auto_in_d_bits_data; // @[LazyModule.scala 355:16]
  assign uncache_io_in_req_valid = core_io_uncache_req_valid; // @[SoC.scala 57:26]
  assign uncache_io_in_req_bits_addr = core_io_uncache_req_bits_addr; // @[SoC.scala 57:26]
  assign uncache_io_in_req_bits_wdata = core_io_uncache_req_bits_wdata; // @[SoC.scala 57:26]
  assign uncache_io_in_req_bits_wmask = core_io_uncache_req_bits_wmask; // @[SoC.scala 57:26]
  assign uncache_io_in_req_bits_wen = core_io_uncache_req_bits_wen; // @[SoC.scala 57:26]
  assign uncache_io_in_req_bits_len = core_io_uncache_req_bits_len; // @[SoC.scala 57:26]
  assign uncache_io_in_resp_ready = core_io_uncache_resp_ready; // @[SoC.scala 57:26]
  assign xbar_clock = clock;
  assign xbar_reset = reset;
  assign xbar_auto_in_2_a_valid = dcache_auto_out_a_valid; // @[LazyModule.scala 355:16]
  assign xbar_auto_in_2_a_bits_source = dcache_auto_out_a_bits_source; // @[LazyModule.scala 355:16]
  assign xbar_auto_in_2_a_bits_address = dcache_auto_out_a_bits_address; // @[LazyModule.scala 355:16]
  assign xbar_auto_in_2_b_ready = dcache_auto_out_b_ready; // @[LazyModule.scala 355:16]
  assign xbar_auto_in_2_c_valid = dcache_auto_out_c_valid; // @[LazyModule.scala 355:16]
  assign xbar_auto_in_2_c_bits_opcode = dcache_auto_out_c_bits_opcode; // @[LazyModule.scala 355:16]
  assign xbar_auto_in_2_c_bits_param = dcache_auto_out_c_bits_param; // @[LazyModule.scala 355:16]
  assign xbar_auto_in_2_c_bits_size = dcache_auto_out_c_bits_size; // @[LazyModule.scala 355:16]
  assign xbar_auto_in_2_c_bits_source = dcache_auto_out_c_bits_source; // @[LazyModule.scala 355:16]
  assign xbar_auto_in_2_c_bits_address = dcache_auto_out_c_bits_address; // @[LazyModule.scala 355:16]
  assign xbar_auto_in_2_c_bits_data = dcache_auto_out_c_bits_data; // @[LazyModule.scala 355:16]
  assign xbar_auto_in_2_d_ready = dcache_auto_out_d_ready; // @[LazyModule.scala 355:16]
  assign xbar_auto_in_2_e_valid = dcache_auto_out_e_valid; // @[LazyModule.scala 355:16]
  assign xbar_auto_in_2_e_bits_sink = dcache_auto_out_e_bits_sink; // @[LazyModule.scala 355:16]
  assign xbar_auto_in_1_a_valid = widget_auto_out_a_valid; // @[LazyModule.scala 353:16]
  assign xbar_auto_in_1_a_bits_opcode = widget_auto_out_a_bits_opcode; // @[LazyModule.scala 353:16]
  assign xbar_auto_in_1_a_bits_size = widget_auto_out_a_bits_size; // @[LazyModule.scala 353:16]
  assign xbar_auto_in_1_a_bits_source = widget_auto_out_a_bits_source; // @[LazyModule.scala 353:16]
  assign xbar_auto_in_1_a_bits_address = widget_auto_out_a_bits_address; // @[LazyModule.scala 353:16]
  assign xbar_auto_in_1_a_bits_mask = widget_auto_out_a_bits_mask; // @[LazyModule.scala 353:16]
  assign xbar_auto_in_1_a_bits_data = widget_auto_out_a_bits_data; // @[LazyModule.scala 353:16]
  assign xbar_auto_in_1_d_ready = widget_auto_out_d_ready; // @[LazyModule.scala 353:16]
  assign xbar_auto_in_0_a_valid = icache_auto_out_a_valid; // @[LazyModule.scala 355:16]
  assign xbar_auto_in_0_a_bits_source = icache_auto_out_a_bits_source; // @[LazyModule.scala 355:16]
  assign xbar_auto_in_0_a_bits_address = icache_auto_out_a_bits_address; // @[LazyModule.scala 355:16]
  assign xbar_auto_in_0_d_ready = icache_auto_out_d_ready; // @[LazyModule.scala 355:16]
  assign xbar_auto_out_a_ready = auto_out_a_ready; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign xbar_auto_out_b_valid = auto_out_b_valid; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign xbar_auto_out_b_bits_size = auto_out_b_bits_size; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign xbar_auto_out_b_bits_source = auto_out_b_bits_source; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign xbar_auto_out_b_bits_address = auto_out_b_bits_address; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign xbar_auto_out_c_ready = auto_out_c_ready; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign xbar_auto_out_d_valid = auto_out_d_valid; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign xbar_auto_out_d_bits_opcode = auto_out_d_bits_opcode; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign xbar_auto_out_d_bits_size = auto_out_d_bits_size; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign xbar_auto_out_d_bits_source = auto_out_d_bits_source; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign xbar_auto_out_d_bits_sink = auto_out_d_bits_sink; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign xbar_auto_out_d_bits_data = auto_out_d_bits_data; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign xbar_auto_out_e_ready = auto_out_e_ready; // @[Nodes.scala 1212:84 LazyModule.scala 368:12]
  assign widget_clock = clock;
  assign widget_reset = reset;
  assign widget_auto_in_a_valid = uncache_auto_out_a_valid; // @[LazyModule.scala 355:16]
  assign widget_auto_in_a_bits_opcode = uncache_auto_out_a_bits_opcode; // @[LazyModule.scala 355:16]
  assign widget_auto_in_a_bits_size = uncache_auto_out_a_bits_size; // @[LazyModule.scala 355:16]
  assign widget_auto_in_a_bits_source = uncache_auto_out_a_bits_source; // @[LazyModule.scala 355:16]
  assign widget_auto_in_a_bits_address = uncache_auto_out_a_bits_address; // @[LazyModule.scala 355:16]
  assign widget_auto_in_a_bits_mask = uncache_auto_out_a_bits_mask; // @[LazyModule.scala 355:16]
  assign widget_auto_in_a_bits_data = uncache_auto_out_a_bits_data; // @[LazyModule.scala 355:16]
  assign widget_auto_in_d_ready = uncache_auto_out_d_ready; // @[LazyModule.scala 355:16]
  assign widget_auto_out_a_ready = xbar_auto_in_1_a_ready; // @[LazyModule.scala 353:16]
  assign widget_auto_out_d_valid = xbar_auto_in_1_d_valid; // @[LazyModule.scala 353:16]
  assign widget_auto_out_d_bits_opcode = xbar_auto_in_1_d_bits_opcode; // @[LazyModule.scala 353:16]
  assign widget_auto_out_d_bits_size = xbar_auto_in_1_d_bits_size; // @[LazyModule.scala 353:16]
  assign widget_auto_out_d_bits_source = xbar_auto_in_1_d_bits_source; // @[LazyModule.scala 353:16]
  assign widget_auto_out_d_bits_data = xbar_auto_in_1_d_bits_data; // @[LazyModule.scala 353:16]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_imem_req_ready = icache_io_cache_req_ready; // @[SoC.scala 46:30]
  assign core_io_imem_resp_valid = icache_io_cache_resp_valid; // @[SoC.scala 46:30]
  assign core_io_imem_resp_bits_rdata = icache_io_cache_resp_bits_rdata; // @[SoC.scala 46:30]
  assign core_io_dmem_req_ready = xbar_1_io_in_0_req_ready; // @[SoC.scala 51:28]
  assign core_io_dmem_resp_valid = xbar_1_io_in_0_resp_valid; // @[SoC.scala 51:28]
  assign core_io_dmem_resp_bits_rdata = xbar_1_io_in_0_resp_bits_rdata; // @[SoC.scala 51:28]
  assign core_io_iptw_req_ready = xbar_1_io_in_1_req_ready; // @[SoC.scala 52:28]
  assign core_io_iptw_resp_valid = xbar_1_io_in_1_resp_valid; // @[SoC.scala 52:28]
  assign core_io_iptw_resp_bits_rdata = xbar_1_io_in_1_resp_bits_rdata; // @[SoC.scala 52:28]
  assign core_io_dptw_req_ready = xbar_1_io_in_2_req_ready; // @[SoC.scala 53:28]
  assign core_io_dptw_resp_valid = xbar_1_io_in_2_resp_valid; // @[SoC.scala 53:28]
  assign core_io_dptw_resp_bits_rdata = xbar_1_io_in_2_resp_bits_rdata; // @[SoC.scala 53:28]
  assign core_io_uncache_req_ready = uncache_io_in_req_ready; // @[SoC.scala 57:26]
  assign core_io_uncache_resp_valid = uncache_io_in_resp_valid; // @[SoC.scala 57:26]
  assign core_io_uncache_resp_bits_rdata = uncache_io_in_resp_bits_rdata; // @[SoC.scala 57:26]
  assign core_io_intr_mtip = io_intr_mtip; // @[SoC.scala 43:18]
  assign core_io_intr_msip = io_intr_msip; // @[SoC.scala 43:18]
  assign core_io_intr_meip = io_intr_meip; // @[SoC.scala 43:18]
  assign core_io_intr_seip = io_intr_seip; // @[SoC.scala 43:18]
  assign xbar_1_clock = clock;
  assign xbar_1_reset = reset;
  assign xbar_1_io_in_0_req_valid = core_io_dmem_req_valid; // @[SoC.scala 51:28]
  assign xbar_1_io_in_0_req_bits_addr = core_io_dmem_req_bits_addr; // @[SoC.scala 51:28]
  assign xbar_1_io_in_0_req_bits_wdata = core_io_dmem_req_bits_wdata; // @[SoC.scala 51:28]
  assign xbar_1_io_in_0_req_bits_wmask = core_io_dmem_req_bits_wmask; // @[SoC.scala 51:28]
  assign xbar_1_io_in_0_req_bits_wen = core_io_dmem_req_bits_wen; // @[SoC.scala 51:28]
  assign xbar_1_io_in_0_req_bits_len = core_io_dmem_req_bits_len; // @[SoC.scala 51:28]
  assign xbar_1_io_in_0_req_bits_lrsc = core_io_dmem_req_bits_lrsc; // @[SoC.scala 51:28]
  assign xbar_1_io_in_0_req_bits_amo = core_io_dmem_req_bits_amo; // @[SoC.scala 51:28]
  assign xbar_1_io_in_0_resp_ready = core_io_dmem_resp_ready; // @[SoC.scala 51:28]
  assign xbar_1_io_in_1_req_valid = core_io_iptw_req_valid; // @[SoC.scala 52:28]
  assign xbar_1_io_in_1_req_bits_addr = core_io_iptw_req_bits_addr; // @[SoC.scala 52:28]
  assign xbar_1_io_in_1_resp_ready = core_io_iptw_resp_ready; // @[SoC.scala 52:28]
  assign xbar_1_io_in_2_req_valid = core_io_dptw_req_valid; // @[SoC.scala 53:28]
  assign xbar_1_io_in_2_req_bits_addr = core_io_dptw_req_bits_addr; // @[SoC.scala 53:28]
  assign xbar_1_io_in_2_resp_ready = core_io_dptw_resp_ready; // @[SoC.scala 53:28]
  assign xbar_1_io_out_req_ready = dcache_io_cache_req_ready; // @[SoC.scala 54:28]
  assign xbar_1_io_out_resp_valid = dcache_io_cache_resp_valid; // @[SoC.scala 54:28]
  assign xbar_1_io_out_resp_bits_rdata = dcache_io_cache_resp_bits_rdata; // @[SoC.scala 54:28]
endmodule
module HellaPeekingArbiter(
  input          clock,
  input          reset,
  output         io_in_0_ready,
  input          io_in_0_valid,
  input  [31:0]  io_in_0_bits_union,
  output         io_in_1_ready,
  input          io_in_1_valid,
  input  [2:0]   io_in_1_bits_opcode,
  input  [2:0]   io_in_1_bits_param,
  input  [2:0]   io_in_1_bits_size,
  input  [3:0]   io_in_1_bits_source,
  input  [31:0]  io_in_1_bits_address,
  input  [255:0] io_in_1_bits_data,
  output         io_in_2_ready,
  input          io_in_2_valid,
  input  [2:0]   io_in_2_bits_opcode,
  input  [2:0]   io_in_2_bits_param,
  input  [2:0]   io_in_2_bits_size,
  input  [3:0]   io_in_2_bits_source,
  input  [31:0]  io_in_2_bits_address,
  input  [255:0] io_in_2_bits_data,
  input  [31:0]  io_in_2_bits_union,
  input          io_out_ready,
  output         io_out_valid,
  output [2:0]   io_out_bits_chanId,
  output [2:0]   io_out_bits_opcode,
  output [2:0]   io_out_bits_param,
  output [2:0]   io_out_bits_size,
  output [3:0]   io_out_bits_source,
  output [31:0]  io_out_bits_address,
  output [255:0] io_out_bits_data,
  output [31:0]  io_out_bits_union,
  output         io_out_bits_last
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] lockIdx; // @[Arbiters.scala 26:24]
  reg  locked; // @[Arbiters.scala 27:23]
  wire [1:0] _choice_T = io_in_1_valid ? 2'h1 : 2'h2; // @[Mux.scala 47:70]
  wire [1:0] choice = io_in_0_valid ? 2'h0 : _choice_T; // @[Mux.scala 47:70]
  wire [1:0] chosen = locked ? lockIdx : choice; // @[Arbiters.scala 37:19]
  wire  _GEN_1 = 2'h1 == chosen ? io_in_1_valid : io_in_0_valid; // @[Arbiters.scala 43:{16,16}]
  wire [2:0] _GEN_4 = 2'h1 == chosen ? 3'h2 : 3'h4; // @[Arbiters.scala 44:{15,15}]
  wire [2:0] _GEN_7 = 2'h1 == chosen ? io_in_1_bits_opcode : 3'h0; // @[Arbiters.scala 44:{15,15}]
  wire [2:0] _GEN_10 = 2'h1 == chosen ? io_in_1_bits_param : 3'h0; // @[Arbiters.scala 44:{15,15}]
  wire [2:0] _GEN_13 = 2'h1 == chosen ? io_in_1_bits_size : 3'h0; // @[Arbiters.scala 44:{15,15}]
  wire [3:0] _GEN_16 = 2'h1 == chosen ? io_in_1_bits_source : 4'h0; // @[Arbiters.scala 44:{15,15}]
  wire [31:0] _GEN_19 = 2'h1 == chosen ? io_in_1_bits_address : 32'h0; // @[Arbiters.scala 44:{15,15}]
  wire [255:0] _GEN_22 = 2'h1 == chosen ? io_in_1_bits_data : 256'h0; // @[Arbiters.scala 44:{15,15}]
  wire [31:0] _GEN_28 = 2'h1 == chosen ? 32'h0 : io_in_0_bits_union; // @[Arbiters.scala 44:{15,15}]
  wire  _T = io_out_ready & io_out_valid; // @[Decoupled.scala 51:35]
  wire  _GEN_34 = ~locked | locked; // @[Arbiters.scala 60:50 62:14 27:23]
  assign io_in_0_ready = io_out_ready & chosen == 2'h0; // @[Arbiters.scala 40:36]
  assign io_in_1_ready = io_out_ready & chosen == 2'h1; // @[Arbiters.scala 40:36]
  assign io_in_2_ready = io_out_ready & chosen == 2'h2; // @[Arbiters.scala 40:36]
  assign io_out_valid = 2'h2 == chosen ? io_in_2_valid : _GEN_1; // @[Arbiters.scala 43:{16,16}]
  assign io_out_bits_chanId = 2'h2 == chosen ? 3'h0 : _GEN_4; // @[Arbiters.scala 44:{15,15}]
  assign io_out_bits_opcode = 2'h2 == chosen ? io_in_2_bits_opcode : _GEN_7; // @[Arbiters.scala 44:{15,15}]
  assign io_out_bits_param = 2'h2 == chosen ? io_in_2_bits_param : _GEN_10; // @[Arbiters.scala 44:{15,15}]
  assign io_out_bits_size = 2'h2 == chosen ? io_in_2_bits_size : _GEN_13; // @[Arbiters.scala 44:{15,15}]
  assign io_out_bits_source = 2'h2 == chosen ? io_in_2_bits_source : _GEN_16; // @[Arbiters.scala 44:{15,15}]
  assign io_out_bits_address = 2'h2 == chosen ? io_in_2_bits_address : _GEN_19; // @[Arbiters.scala 44:{15,15}]
  assign io_out_bits_data = 2'h2 == chosen ? io_in_2_bits_data : _GEN_22; // @[Arbiters.scala 44:{15,15}]
  assign io_out_bits_union = 2'h2 == chosen ? io_in_2_bits_union : _GEN_28; // @[Arbiters.scala 44:{15,15}]
  assign io_out_bits_last = 1'h1; // @[Arbiters.scala 44:{15,15}]
  always @(posedge clock) begin
    if (reset) begin // @[Arbiters.scala 26:24]
      lockIdx <= 2'h0; // @[Arbiters.scala 26:24]
    end else if (_T) begin // @[Arbiters.scala 59:22]
      if (~locked) begin // @[Arbiters.scala 60:50]
        if (io_in_0_valid) begin // @[Mux.scala 47:70]
          lockIdx <= 2'h0;
        end else begin
          lockIdx <= _choice_T;
        end
      end
    end
    if (reset) begin // @[Arbiters.scala 27:23]
      locked <= 1'h0; // @[Arbiters.scala 27:23]
    end else if (_T) begin // @[Arbiters.scala 59:22]
      if (io_out_bits_last) begin // @[Arbiters.scala 65:35]
        locked <= 1'h0; // @[Arbiters.scala 66:14]
      end else begin
        locked <= _GEN_34;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lockIdx = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  locked = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module GenericSerializer(
  input          clock,
  input          reset,
  output         io_in_ready,
  input          io_in_valid,
  input  [2:0]   io_in_bits_chanId,
  input  [2:0]   io_in_bits_opcode,
  input  [2:0]   io_in_bits_param,
  input  [2:0]   io_in_bits_size,
  input  [3:0]   io_in_bits_source,
  input  [31:0]  io_in_bits_address,
  input  [255:0] io_in_bits_data,
  input  [31:0]  io_in_bits_union,
  input          io_out_ready,
  output         io_out_valid,
  output [7:0]   io_out_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [351:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [337:0] data; // @[Serdes.scala 173:22]
  reg  sending; // @[Serdes.scala 175:38]
  wire  _T = io_out_ready & io_out_valid; // @[Decoupled.scala 51:35]
  reg [5:0] sendCount; // @[Counter.scala 61:40]
  wire  wrap_wrap = sendCount == 6'h2a; // @[Counter.scala 73:24]
  wire [5:0] _wrap_value_T_1 = sendCount + 6'h1; // @[Counter.scala 77:24]
  wire  sendDone = _T & wrap_wrap; // @[Counter.scala 118:{16,23} 117:24]
  wire  _T_1 = io_in_ready & io_in_valid; // @[Decoupled.scala 51:35]
  wire [337:0] _data_T = {io_in_bits_chanId,io_in_bits_opcode,io_in_bits_param,io_in_bits_size,io_in_bits_source,
    io_in_bits_address,io_in_bits_data,1'h0,io_in_bits_union,1'h1}; // @[Serdes.scala 183:27]
  wire  _GEN_4 = _T_1 | sending; // @[Serdes.scala 182:20 184:13 175:38]
  wire [337:0] _data_T_1 = {{8'd0}, data[337:8]}; // @[Serdes.scala 187:36]
  assign io_in_ready = ~sending; // @[Serdes.scala 178:19]
  assign io_out_valid = sending; // @[Serdes.scala 179:16]
  assign io_out_bits = data[7:0]; // @[Serdes.scala 180:23]
  always @(posedge clock) begin
    if (_T) begin // @[Serdes.scala 187:21]
      data <= _data_T_1; // @[Serdes.scala 187:28]
    end else if (_T_1) begin // @[Serdes.scala 182:20]
      data <= _data_T; // @[Serdes.scala 183:13]
    end
    if (reset) begin // @[Serdes.scala 175:38]
      sending <= 1'h0; // @[Serdes.scala 175:38]
    end else if (sendDone) begin // @[Serdes.scala 189:18]
      sending <= 1'h0; // @[Serdes.scala 189:28]
    end else begin
      sending <= _GEN_4;
    end
    if (reset) begin // @[Counter.scala 61:40]
      sendCount <= 6'h0; // @[Counter.scala 61:40]
    end else if (_T) begin // @[Counter.scala 118:16]
      if (wrap_wrap) begin // @[Counter.scala 87:20]
        sendCount <= 6'h0; // @[Counter.scala 87:28]
      end else begin
        sendCount <= _wrap_value_T_1; // @[Counter.scala 77:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {11{`RANDOM}};
  data = _RAND_0[337:0];
  _RAND_1 = {1{`RANDOM}};
  sending = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  sendCount = _RAND_2[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module GenericDeserializer(
  input          clock,
  input          reset,
  output         io_in_ready,
  input          io_in_valid,
  input  [7:0]   io_in_bits,
  input          io_out_ready,
  output         io_out_valid,
  output [2:0]   io_out_bits_chanId,
  output [2:0]   io_out_bits_opcode,
  output [2:0]   io_out_bits_size,
  output [3:0]   io_out_bits_source,
  output [31:0]  io_out_bits_address,
  output [255:0] io_out_bits_data,
  output [31:0]  io_out_bits_union
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] data_0; // @[Serdes.scala 200:22]
  reg [7:0] data_1; // @[Serdes.scala 200:22]
  reg [7:0] data_2; // @[Serdes.scala 200:22]
  reg [7:0] data_3; // @[Serdes.scala 200:22]
  reg [7:0] data_4; // @[Serdes.scala 200:22]
  reg [7:0] data_5; // @[Serdes.scala 200:22]
  reg [7:0] data_6; // @[Serdes.scala 200:22]
  reg [7:0] data_7; // @[Serdes.scala 200:22]
  reg [7:0] data_8; // @[Serdes.scala 200:22]
  reg [7:0] data_9; // @[Serdes.scala 200:22]
  reg [7:0] data_10; // @[Serdes.scala 200:22]
  reg [7:0] data_11; // @[Serdes.scala 200:22]
  reg [7:0] data_12; // @[Serdes.scala 200:22]
  reg [7:0] data_13; // @[Serdes.scala 200:22]
  reg [7:0] data_14; // @[Serdes.scala 200:22]
  reg [7:0] data_15; // @[Serdes.scala 200:22]
  reg [7:0] data_16; // @[Serdes.scala 200:22]
  reg [7:0] data_17; // @[Serdes.scala 200:22]
  reg [7:0] data_18; // @[Serdes.scala 200:22]
  reg [7:0] data_19; // @[Serdes.scala 200:22]
  reg [7:0] data_20; // @[Serdes.scala 200:22]
  reg [7:0] data_21; // @[Serdes.scala 200:22]
  reg [7:0] data_22; // @[Serdes.scala 200:22]
  reg [7:0] data_23; // @[Serdes.scala 200:22]
  reg [7:0] data_24; // @[Serdes.scala 200:22]
  reg [7:0] data_25; // @[Serdes.scala 200:22]
  reg [7:0] data_26; // @[Serdes.scala 200:22]
  reg [7:0] data_27; // @[Serdes.scala 200:22]
  reg [7:0] data_28; // @[Serdes.scala 200:22]
  reg [7:0] data_29; // @[Serdes.scala 200:22]
  reg [7:0] data_30; // @[Serdes.scala 200:22]
  reg [7:0] data_31; // @[Serdes.scala 200:22]
  reg [7:0] data_32; // @[Serdes.scala 200:22]
  reg [7:0] data_33; // @[Serdes.scala 200:22]
  reg [7:0] data_34; // @[Serdes.scala 200:22]
  reg [7:0] data_35; // @[Serdes.scala 200:22]
  reg [7:0] data_36; // @[Serdes.scala 200:22]
  reg [7:0] data_37; // @[Serdes.scala 200:22]
  reg [7:0] data_38; // @[Serdes.scala 200:22]
  reg [7:0] data_39; // @[Serdes.scala 200:22]
  reg [7:0] data_40; // @[Serdes.scala 200:22]
  reg [7:0] data_41; // @[Serdes.scala 200:22]
  reg [7:0] data_42; // @[Serdes.scala 200:22]
  reg  receiving; // @[Serdes.scala 202:38]
  wire  _T = io_in_ready & io_in_valid; // @[Decoupled.scala 51:35]
  reg [5:0] recvCount; // @[Counter.scala 61:40]
  wire  wrap_wrap = recvCount == 6'h2a; // @[Counter.scala 73:24]
  wire [5:0] _wrap_value_T_1 = recvCount + 6'h1; // @[Counter.scala 77:24]
  wire  recvDone = _T & wrap_wrap; // @[Counter.scala 118:{16,23} 117:24]
  wire [79:0] io_out_bits_lo_lo = {data_9,data_8,data_7,data_6,data_5,data_4,data_3,data_2,data_1,data_0}; // @[Serdes.scala 207:24]
  wire [39:0] io_out_bits_lo_hi_lo = {data_14,data_13,data_12,data_11,data_10}; // @[Serdes.scala 207:24]
  wire [167:0] io_out_bits_lo = {data_20,data_19,data_18,data_17,data_16,data_15,io_out_bits_lo_hi_lo,io_out_bits_lo_lo}
    ; // @[Serdes.scala 207:24]
  wire [39:0] io_out_bits_hi_lo_lo = {data_25,data_24,data_23,data_22,data_21}; // @[Serdes.scala 207:24]
  wire [87:0] io_out_bits_hi_lo = {data_31,data_30,data_29,data_28,data_27,data_26,io_out_bits_hi_lo_lo}; // @[Serdes.scala 207:24]
  wire [39:0] io_out_bits_hi_hi_lo = {data_36,data_35,data_34,data_33,data_32}; // @[Serdes.scala 207:24]
  wire [343:0] _io_out_bits_T = {data_42,data_41,data_40,data_39,data_38,data_37,io_out_bits_hi_hi_lo,io_out_bits_hi_lo,
    io_out_bits_lo}; // @[Serdes.scala 207:24]
  wire  _GEN_89 = recvDone ? 1'h0 : receiving; // @[Serdes.scala 213:{18,30} 202:38]
  wire  _T_2 = io_out_ready & io_out_valid; // @[Decoupled.scala 51:35]
  wire  _GEN_90 = _T_2 | _GEN_89; // @[Serdes.scala 215:{21,33}]
  assign io_in_ready = receiving; // @[Serdes.scala 205:16]
  assign io_out_valid = ~receiving; // @[Serdes.scala 206:19]
  assign io_out_bits_chanId = _io_out_bits_T[337:335]; // @[Serdes.scala 207:39]
  assign io_out_bits_opcode = _io_out_bits_T[334:332]; // @[Serdes.scala 207:39]
  assign io_out_bits_size = _io_out_bits_T[328:326]; // @[Serdes.scala 207:39]
  assign io_out_bits_source = _io_out_bits_T[325:322]; // @[Serdes.scala 207:39]
  assign io_out_bits_address = _io_out_bits_T[321:290]; // @[Serdes.scala 207:39]
  assign io_out_bits_data = _io_out_bits_T[289:34]; // @[Serdes.scala 207:39]
  assign io_out_bits_union = _io_out_bits_T[32:1]; // @[Serdes.scala 207:39]
  always @(posedge clock) begin
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h0 == recvCount) begin // @[Serdes.scala 210:21]
        data_0 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h1 == recvCount) begin // @[Serdes.scala 210:21]
        data_1 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h2 == recvCount) begin // @[Serdes.scala 210:21]
        data_2 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h3 == recvCount) begin // @[Serdes.scala 210:21]
        data_3 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h4 == recvCount) begin // @[Serdes.scala 210:21]
        data_4 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h5 == recvCount) begin // @[Serdes.scala 210:21]
        data_5 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h6 == recvCount) begin // @[Serdes.scala 210:21]
        data_6 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h7 == recvCount) begin // @[Serdes.scala 210:21]
        data_7 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h8 == recvCount) begin // @[Serdes.scala 210:21]
        data_8 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h9 == recvCount) begin // @[Serdes.scala 210:21]
        data_9 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'ha == recvCount) begin // @[Serdes.scala 210:21]
        data_10 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'hb == recvCount) begin // @[Serdes.scala 210:21]
        data_11 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'hc == recvCount) begin // @[Serdes.scala 210:21]
        data_12 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'hd == recvCount) begin // @[Serdes.scala 210:21]
        data_13 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'he == recvCount) begin // @[Serdes.scala 210:21]
        data_14 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'hf == recvCount) begin // @[Serdes.scala 210:21]
        data_15 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h10 == recvCount) begin // @[Serdes.scala 210:21]
        data_16 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h11 == recvCount) begin // @[Serdes.scala 210:21]
        data_17 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h12 == recvCount) begin // @[Serdes.scala 210:21]
        data_18 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h13 == recvCount) begin // @[Serdes.scala 210:21]
        data_19 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h14 == recvCount) begin // @[Serdes.scala 210:21]
        data_20 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h15 == recvCount) begin // @[Serdes.scala 210:21]
        data_21 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h16 == recvCount) begin // @[Serdes.scala 210:21]
        data_22 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h17 == recvCount) begin // @[Serdes.scala 210:21]
        data_23 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h18 == recvCount) begin // @[Serdes.scala 210:21]
        data_24 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h19 == recvCount) begin // @[Serdes.scala 210:21]
        data_25 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h1a == recvCount) begin // @[Serdes.scala 210:21]
        data_26 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h1b == recvCount) begin // @[Serdes.scala 210:21]
        data_27 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h1c == recvCount) begin // @[Serdes.scala 210:21]
        data_28 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h1d == recvCount) begin // @[Serdes.scala 210:21]
        data_29 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h1e == recvCount) begin // @[Serdes.scala 210:21]
        data_30 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h1f == recvCount) begin // @[Serdes.scala 210:21]
        data_31 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h20 == recvCount) begin // @[Serdes.scala 210:21]
        data_32 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h21 == recvCount) begin // @[Serdes.scala 210:21]
        data_33 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h22 == recvCount) begin // @[Serdes.scala 210:21]
        data_34 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h23 == recvCount) begin // @[Serdes.scala 210:21]
        data_35 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h24 == recvCount) begin // @[Serdes.scala 210:21]
        data_36 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h25 == recvCount) begin // @[Serdes.scala 210:21]
        data_37 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h26 == recvCount) begin // @[Serdes.scala 210:21]
        data_38 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h27 == recvCount) begin // @[Serdes.scala 210:21]
        data_39 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h28 == recvCount) begin // @[Serdes.scala 210:21]
        data_40 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h29 == recvCount) begin // @[Serdes.scala 210:21]
        data_41 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    if (_T) begin // @[Serdes.scala 209:20]
      if (6'h2a == recvCount) begin // @[Serdes.scala 210:21]
        data_42 <= io_in_bits; // @[Serdes.scala 210:21]
      end
    end
    receiving <= reset | _GEN_90; // @[Serdes.scala 202:{38,38}]
    if (reset) begin // @[Counter.scala 61:40]
      recvCount <= 6'h0; // @[Counter.scala 61:40]
    end else if (_T) begin // @[Counter.scala 118:16]
      if (wrap_wrap) begin // @[Counter.scala 87:20]
        recvCount <= 6'h0; // @[Counter.scala 87:28]
      end else begin
        recvCount <= _wrap_value_T_1; // @[Counter.scala 77:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  data_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  data_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  data_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  data_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  data_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  data_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  data_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  data_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  data_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  data_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  data_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  data_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  data_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  data_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  data_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  data_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  data_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  data_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  data_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  data_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  data_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  data_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  data_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  data_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  data_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  data_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  data_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  data_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  data_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  data_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  data_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  data_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  data_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  data_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  data_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  data_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  data_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  data_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  data_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  receiving = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  recvCount = _RAND_44[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLSerdes(
  input          clock,
  input          reset,
  output         auto_in_a_ready,
  input          auto_in_a_valid,
  input  [2:0]   auto_in_a_bits_opcode,
  input  [2:0]   auto_in_a_bits_param,
  input  [2:0]   auto_in_a_bits_size,
  input  [3:0]   auto_in_a_bits_source,
  input  [31:0]  auto_in_a_bits_address,
  input  [31:0]  auto_in_a_bits_mask,
  input  [255:0] auto_in_a_bits_data,
  input          auto_in_b_ready,
  output         auto_in_b_valid,
  output [2:0]   auto_in_b_bits_size,
  output [3:0]   auto_in_b_bits_source,
  output [31:0]  auto_in_b_bits_address,
  output         auto_in_c_ready,
  input          auto_in_c_valid,
  input  [2:0]   auto_in_c_bits_opcode,
  input  [2:0]   auto_in_c_bits_param,
  input  [2:0]   auto_in_c_bits_size,
  input  [3:0]   auto_in_c_bits_source,
  input  [31:0]  auto_in_c_bits_address,
  input  [255:0] auto_in_c_bits_data,
  input          auto_in_d_ready,
  output         auto_in_d_valid,
  output [2:0]   auto_in_d_bits_opcode,
  output [2:0]   auto_in_d_bits_size,
  output [3:0]   auto_in_d_bits_source,
  output [5:0]   auto_in_d_bits_sink,
  output [255:0] auto_in_d_bits_data,
  output         auto_in_e_ready,
  input          auto_in_e_valid,
  input  [5:0]   auto_in_e_bits_sink,
  output         io_ser_0_in_ready,
  input          io_ser_0_in_valid,
  input  [7:0]   io_ser_0_in_bits,
  input          io_ser_0_out_ready,
  output         io_ser_0_out_valid,
  output [7:0]   io_ser_0_out_bits
);
  wire  outArb_clock; // @[Serdes.scala 568:33]
  wire  outArb_reset; // @[Serdes.scala 568:33]
  wire  outArb_io_in_0_ready; // @[Serdes.scala 568:33]
  wire  outArb_io_in_0_valid; // @[Serdes.scala 568:33]
  wire [31:0] outArb_io_in_0_bits_union; // @[Serdes.scala 568:33]
  wire  outArb_io_in_1_ready; // @[Serdes.scala 568:33]
  wire  outArb_io_in_1_valid; // @[Serdes.scala 568:33]
  wire [2:0] outArb_io_in_1_bits_opcode; // @[Serdes.scala 568:33]
  wire [2:0] outArb_io_in_1_bits_param; // @[Serdes.scala 568:33]
  wire [2:0] outArb_io_in_1_bits_size; // @[Serdes.scala 568:33]
  wire [3:0] outArb_io_in_1_bits_source; // @[Serdes.scala 568:33]
  wire [31:0] outArb_io_in_1_bits_address; // @[Serdes.scala 568:33]
  wire [255:0] outArb_io_in_1_bits_data; // @[Serdes.scala 568:33]
  wire  outArb_io_in_2_ready; // @[Serdes.scala 568:33]
  wire  outArb_io_in_2_valid; // @[Serdes.scala 568:33]
  wire [2:0] outArb_io_in_2_bits_opcode; // @[Serdes.scala 568:33]
  wire [2:0] outArb_io_in_2_bits_param; // @[Serdes.scala 568:33]
  wire [2:0] outArb_io_in_2_bits_size; // @[Serdes.scala 568:33]
  wire [3:0] outArb_io_in_2_bits_source; // @[Serdes.scala 568:33]
  wire [31:0] outArb_io_in_2_bits_address; // @[Serdes.scala 568:33]
  wire [255:0] outArb_io_in_2_bits_data; // @[Serdes.scala 568:33]
  wire [31:0] outArb_io_in_2_bits_union; // @[Serdes.scala 568:33]
  wire  outArb_io_out_ready; // @[Serdes.scala 568:33]
  wire  outArb_io_out_valid; // @[Serdes.scala 568:33]
  wire [2:0] outArb_io_out_bits_chanId; // @[Serdes.scala 568:33]
  wire [2:0] outArb_io_out_bits_opcode; // @[Serdes.scala 568:33]
  wire [2:0] outArb_io_out_bits_param; // @[Serdes.scala 568:33]
  wire [2:0] outArb_io_out_bits_size; // @[Serdes.scala 568:33]
  wire [3:0] outArb_io_out_bits_source; // @[Serdes.scala 568:33]
  wire [31:0] outArb_io_out_bits_address; // @[Serdes.scala 568:33]
  wire [255:0] outArb_io_out_bits_data; // @[Serdes.scala 568:33]
  wire [31:0] outArb_io_out_bits_union; // @[Serdes.scala 568:33]
  wire  outArb_io_out_bits_last; // @[Serdes.scala 568:33]
  wire  outSer_clock; // @[Serdes.scala 569:33]
  wire  outSer_reset; // @[Serdes.scala 569:33]
  wire  outSer_io_in_ready; // @[Serdes.scala 569:33]
  wire  outSer_io_in_valid; // @[Serdes.scala 569:33]
  wire [2:0] outSer_io_in_bits_chanId; // @[Serdes.scala 569:33]
  wire [2:0] outSer_io_in_bits_opcode; // @[Serdes.scala 569:33]
  wire [2:0] outSer_io_in_bits_param; // @[Serdes.scala 569:33]
  wire [2:0] outSer_io_in_bits_size; // @[Serdes.scala 569:33]
  wire [3:0] outSer_io_in_bits_source; // @[Serdes.scala 569:33]
  wire [31:0] outSer_io_in_bits_address; // @[Serdes.scala 569:33]
  wire [255:0] outSer_io_in_bits_data; // @[Serdes.scala 569:33]
  wire [31:0] outSer_io_in_bits_union; // @[Serdes.scala 569:33]
  wire  outSer_io_out_ready; // @[Serdes.scala 569:33]
  wire  outSer_io_out_valid; // @[Serdes.scala 569:33]
  wire [7:0] outSer_io_out_bits; // @[Serdes.scala 569:33]
  wire  inDes_clock; // @[Serdes.scala 574:27]
  wire  inDes_reset; // @[Serdes.scala 574:27]
  wire  inDes_io_in_ready; // @[Serdes.scala 574:27]
  wire  inDes_io_in_valid; // @[Serdes.scala 574:27]
  wire [7:0] inDes_io_in_bits; // @[Serdes.scala 574:27]
  wire  inDes_io_out_ready; // @[Serdes.scala 574:27]
  wire  inDes_io_out_valid; // @[Serdes.scala 574:27]
  wire [2:0] inDes_io_out_bits_chanId; // @[Serdes.scala 574:27]
  wire [2:0] inDes_io_out_bits_opcode; // @[Serdes.scala 574:27]
  wire [2:0] inDes_io_out_bits_size; // @[Serdes.scala 574:27]
  wire [3:0] inDes_io_out_bits_source; // @[Serdes.scala 574:27]
  wire [31:0] inDes_io_out_bits_address; // @[Serdes.scala 574:27]
  wire [255:0] inDes_io_out_bits_data; // @[Serdes.scala 574:27]
  wire [31:0] inDes_io_out_bits_union; // @[Serdes.scala 574:27]
  wire [6:0] _outChannels_merged_bits_merged_union_T = {auto_in_e_bits_sink,1'h0}; // @[Cat.scala 33:92]
  wire  _bundleIn_0_b_valid_T = inDes_io_out_bits_chanId == 3'h1; // @[Serdes.scala 235:37]
  wire  _bundleIn_0_d_valid_T = inDes_io_out_bits_chanId == 3'h3; // @[Serdes.scala 237:37]
  wire [31:0] _bundleIn_0_d_bits_d_sink_T = {{1'd0}, inDes_io_out_bits_union[31:1]}; // @[Serdes.scala 486:31]
  HellaPeekingArbiter outArb ( // @[Serdes.scala 568:33]
    .clock(outArb_clock),
    .reset(outArb_reset),
    .io_in_0_ready(outArb_io_in_0_ready),
    .io_in_0_valid(outArb_io_in_0_valid),
    .io_in_0_bits_union(outArb_io_in_0_bits_union),
    .io_in_1_ready(outArb_io_in_1_ready),
    .io_in_1_valid(outArb_io_in_1_valid),
    .io_in_1_bits_opcode(outArb_io_in_1_bits_opcode),
    .io_in_1_bits_param(outArb_io_in_1_bits_param),
    .io_in_1_bits_size(outArb_io_in_1_bits_size),
    .io_in_1_bits_source(outArb_io_in_1_bits_source),
    .io_in_1_bits_address(outArb_io_in_1_bits_address),
    .io_in_1_bits_data(outArb_io_in_1_bits_data),
    .io_in_2_ready(outArb_io_in_2_ready),
    .io_in_2_valid(outArb_io_in_2_valid),
    .io_in_2_bits_opcode(outArb_io_in_2_bits_opcode),
    .io_in_2_bits_param(outArb_io_in_2_bits_param),
    .io_in_2_bits_size(outArb_io_in_2_bits_size),
    .io_in_2_bits_source(outArb_io_in_2_bits_source),
    .io_in_2_bits_address(outArb_io_in_2_bits_address),
    .io_in_2_bits_data(outArb_io_in_2_bits_data),
    .io_in_2_bits_union(outArb_io_in_2_bits_union),
    .io_out_ready(outArb_io_out_ready),
    .io_out_valid(outArb_io_out_valid),
    .io_out_bits_chanId(outArb_io_out_bits_chanId),
    .io_out_bits_opcode(outArb_io_out_bits_opcode),
    .io_out_bits_param(outArb_io_out_bits_param),
    .io_out_bits_size(outArb_io_out_bits_size),
    .io_out_bits_source(outArb_io_out_bits_source),
    .io_out_bits_address(outArb_io_out_bits_address),
    .io_out_bits_data(outArb_io_out_bits_data),
    .io_out_bits_union(outArb_io_out_bits_union),
    .io_out_bits_last(outArb_io_out_bits_last)
  );
  GenericSerializer outSer ( // @[Serdes.scala 569:33]
    .clock(outSer_clock),
    .reset(outSer_reset),
    .io_in_ready(outSer_io_in_ready),
    .io_in_valid(outSer_io_in_valid),
    .io_in_bits_chanId(outSer_io_in_bits_chanId),
    .io_in_bits_opcode(outSer_io_in_bits_opcode),
    .io_in_bits_param(outSer_io_in_bits_param),
    .io_in_bits_size(outSer_io_in_bits_size),
    .io_in_bits_source(outSer_io_in_bits_source),
    .io_in_bits_address(outSer_io_in_bits_address),
    .io_in_bits_data(outSer_io_in_bits_data),
    .io_in_bits_union(outSer_io_in_bits_union),
    .io_out_ready(outSer_io_out_ready),
    .io_out_valid(outSer_io_out_valid),
    .io_out_bits(outSer_io_out_bits)
  );
  GenericDeserializer inDes ( // @[Serdes.scala 574:27]
    .clock(inDes_clock),
    .reset(inDes_reset),
    .io_in_ready(inDes_io_in_ready),
    .io_in_valid(inDes_io_in_valid),
    .io_in_bits(inDes_io_in_bits),
    .io_out_ready(inDes_io_out_ready),
    .io_out_valid(inDes_io_out_valid),
    .io_out_bits_chanId(inDes_io_out_bits_chanId),
    .io_out_bits_opcode(inDes_io_out_bits_opcode),
    .io_out_bits_size(inDes_io_out_bits_size),
    .io_out_bits_source(inDes_io_out_bits_source),
    .io_out_bits_address(inDes_io_out_bits_address),
    .io_out_bits_data(inDes_io_out_bits_data),
    .io_out_bits_union(inDes_io_out_bits_union)
  );
  assign auto_in_a_ready = outArb_io_in_2_ready; // @[Serdes.scala 363:22 570:22]
  assign auto_in_b_valid = inDes_io_out_valid & _bundleIn_0_b_valid_T; // @[Serdes.scala 576:43]
  assign auto_in_b_bits_size = inDes_io_out_bits_size; // @[Serdes.scala 413:17 416:15]
  assign auto_in_b_bits_source = inDes_io_out_bits_source; // @[Serdes.scala 413:17 417:15]
  assign auto_in_b_bits_address = inDes_io_out_bits_address; // @[Serdes.scala 413:17 418:15]
  assign auto_in_c_ready = outArb_io_in_1_ready; // @[Serdes.scala 363:22 570:22]
  assign auto_in_d_valid = inDes_io_out_valid & _bundleIn_0_d_valid_T; // @[Serdes.scala 578:43]
  assign auto_in_d_bits_opcode = inDes_io_out_bits_opcode; // @[Serdes.scala 478:17 479:14]
  assign auto_in_d_bits_size = inDes_io_out_bits_size; // @[Serdes.scala 478:17 481:14]
  assign auto_in_d_bits_source = inDes_io_out_bits_source; // @[Serdes.scala 478:17 482:14]
  assign auto_in_d_bits_sink = _bundleIn_0_d_bits_d_sink_T[5:0]; // @[Serdes.scala 478:17 486:17]
  assign auto_in_d_bits_data = inDes_io_out_bits_data; // @[Serdes.scala 478:17 483:14]
  assign auto_in_e_ready = outArb_io_in_0_ready; // @[Serdes.scala 363:22 570:22]
  assign io_ser_0_in_ready = inDes_io_in_ready; // @[Serdes.scala 575:21]
  assign io_ser_0_out_valid = outSer_io_out_valid; // @[Serdes.scala 572:22]
  assign io_ser_0_out_bits = outSer_io_out_bits; // @[Serdes.scala 572:22]
  assign outArb_clock = clock;
  assign outArb_reset = reset;
  assign outArb_io_in_0_valid = auto_in_e_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign outArb_io_in_0_bits_union = {{25'd0}, _outChannels_merged_bits_merged_union_T}; // @[Serdes.scala 330:22 340:26]
  assign outArb_io_in_1_valid = auto_in_c_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign outArb_io_in_1_bits_opcode = auto_in_c_bits_opcode; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign outArb_io_in_1_bits_param = auto_in_c_bits_param; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign outArb_io_in_1_bits_size = auto_in_c_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign outArb_io_in_1_bits_source = auto_in_c_bits_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign outArb_io_in_1_bits_address = auto_in_c_bits_address; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign outArb_io_in_1_bits_data = auto_in_c_bits_data; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign outArb_io_in_2_valid = auto_in_a_valid; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign outArb_io_in_2_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign outArb_io_in_2_bits_param = auto_in_a_bits_param; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign outArb_io_in_2_bits_size = auto_in_a_bits_size; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign outArb_io_in_2_bits_source = auto_in_a_bits_source; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign outArb_io_in_2_bits_address = auto_in_a_bits_address; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign outArb_io_in_2_bits_data = auto_in_a_bits_data; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign outArb_io_in_2_bits_union = auto_in_a_bits_mask; // @[Nodes.scala 1215:84 LazyModule.scala 366:16]
  assign outArb_io_out_ready = outSer_io_in_ready; // @[Serdes.scala 571:22]
  assign outSer_clock = clock;
  assign outSer_reset = reset;
  assign outSer_io_in_valid = outArb_io_out_valid; // @[Serdes.scala 571:22]
  assign outSer_io_in_bits_chanId = outArb_io_out_bits_chanId; // @[Serdes.scala 571:22]
  assign outSer_io_in_bits_opcode = outArb_io_out_bits_opcode; // @[Serdes.scala 571:22]
  assign outSer_io_in_bits_param = outArb_io_out_bits_param; // @[Serdes.scala 571:22]
  assign outSer_io_in_bits_size = outArb_io_out_bits_size; // @[Serdes.scala 571:22]
  assign outSer_io_in_bits_source = outArb_io_out_bits_source; // @[Serdes.scala 571:22]
  assign outSer_io_in_bits_address = outArb_io_out_bits_address; // @[Serdes.scala 571:22]
  assign outSer_io_in_bits_data = outArb_io_out_bits_data; // @[Serdes.scala 571:22]
  assign outSer_io_in_bits_union = outArb_io_out_bits_union; // @[Serdes.scala 571:22]
  assign outSer_io_out_ready = io_ser_0_out_ready; // @[Serdes.scala 572:22]
  assign inDes_clock = clock;
  assign inDes_reset = reset;
  assign inDes_io_in_valid = io_ser_0_in_valid; // @[Serdes.scala 575:21]
  assign inDes_io_in_bits = io_ser_0_in_bits; // @[Serdes.scala 575:21]
  assign inDes_io_out_ready = 3'h3 == inDes_io_out_bits_chanId ? auto_in_d_ready : 3'h1 == inDes_io_out_bits_chanId &
    auto_in_b_ready; // @[Mux.scala 81:58]
endmodule
module TLTraceBuffer(
  input          clock,
  input          reset,
  output         auto_in_a_ready,
  input          auto_in_a_valid,
  input  [2:0]   auto_in_a_bits_opcode,
  input  [2:0]   auto_in_a_bits_param,
  input  [2:0]   auto_in_a_bits_size,
  input  [3:0]   auto_in_a_bits_source,
  input  [31:0]  auto_in_a_bits_address,
  input  [31:0]  auto_in_a_bits_mask,
  input  [255:0] auto_in_a_bits_data,
  input          auto_in_b_ready,
  output         auto_in_b_valid,
  output [2:0]   auto_in_b_bits_size,
  output [3:0]   auto_in_b_bits_source,
  output [31:0]  auto_in_b_bits_address,
  output         auto_in_c_ready,
  input          auto_in_c_valid,
  input  [2:0]   auto_in_c_bits_opcode,
  input  [2:0]   auto_in_c_bits_param,
  input  [2:0]   auto_in_c_bits_size,
  input  [3:0]   auto_in_c_bits_source,
  input  [31:0]  auto_in_c_bits_address,
  input  [255:0] auto_in_c_bits_data,
  input          auto_in_d_ready,
  output         auto_in_d_valid,
  output [2:0]   auto_in_d_bits_opcode,
  output [2:0]   auto_in_d_bits_size,
  output [3:0]   auto_in_d_bits_source,
  output [5:0]   auto_in_d_bits_sink,
  output [255:0] auto_in_d_bits_data,
  output         auto_in_e_ready,
  input          auto_in_e_valid,
  input  [5:0]   auto_in_e_bits_sink,
  input          auto_out_a_ready,
  output         auto_out_a_valid,
  output [2:0]   auto_out_a_bits_opcode,
  output [2:0]   auto_out_a_bits_param,
  output [2:0]   auto_out_a_bits_size,
  output [3:0]   auto_out_a_bits_source,
  output [31:0]  auto_out_a_bits_address,
  output [31:0]  auto_out_a_bits_mask,
  output [255:0] auto_out_a_bits_data,
  output         auto_out_b_ready,
  input          auto_out_b_valid,
  input  [2:0]   auto_out_b_bits_size,
  input  [3:0]   auto_out_b_bits_source,
  input  [31:0]  auto_out_b_bits_address,
  input          auto_out_c_ready,
  output         auto_out_c_valid,
  output [2:0]   auto_out_c_bits_opcode,
  output [2:0]   auto_out_c_bits_param,
  output [2:0]   auto_out_c_bits_size,
  output [3:0]   auto_out_c_bits_source,
  output [31:0]  auto_out_c_bits_address,
  output [255:0] auto_out_c_bits_data,
  output         auto_out_d_ready,
  input          auto_out_d_valid,
  input  [2:0]   auto_out_d_bits_opcode,
  input  [2:0]   auto_out_d_bits_size,
  input  [3:0]   auto_out_d_bits_source,
  input  [5:0]   auto_out_d_bits_sink,
  input  [255:0] auto_out_d_bits_data,
  input          auto_out_e_ready,
  output         auto_out_e_valid,
  output [5:0]   auto_out_e_bits_sink
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [255:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [255:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [255:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
`endif // RANDOMIZE_REG_INIT
  reg  in_a_scan_valid; // @[Utils.scala 36:20]
  wire  _x1_a_ready_T_1 = auto_out_a_ready & in_a_scan_valid; // @[Decoupled.scala 51:35]
  wire  tl_in_a_ready = ~in_a_scan_valid | _x1_a_ready_T_1; // @[TLTraceBuffer.scala 30:38]
  wire  _in_a_scan_bits_T = tl_in_a_ready & auto_in_a_valid; // @[Decoupled.scala 51:35]
  reg [2:0] in_a_scan_bits_opcode; // @[Reg.scala 35:20]
  reg [2:0] in_a_scan_bits_param; // @[Reg.scala 35:20]
  reg [2:0] in_a_scan_bits_size; // @[Reg.scala 35:20]
  reg [3:0] in_a_scan_bits_source; // @[Reg.scala 35:20]
  reg [31:0] in_a_scan_bits_address; // @[Reg.scala 35:20]
  reg [31:0] in_a_scan_bits_mask; // @[Reg.scala 35:20]
  reg [255:0] in_a_scan_bits_data; // @[Reg.scala 35:20]
  wire  _GEN_8 = _x1_a_ready_T_1 ? 1'h0 : in_a_scan_valid; // @[Utils.scala 38:18 36:20 38:22]
  wire  _GEN_9 = _in_a_scan_bits_T | _GEN_8; // @[Utils.scala 39:{19,23}]
  reg  out_b_scan_valid; // @[Utils.scala 36:20]
  wire  _x1_b_ready_T_1 = auto_in_b_ready & out_b_scan_valid; // @[Decoupled.scala 51:35]
  wire  tl_out_b_ready = ~out_b_scan_valid | _x1_b_ready_T_1; // @[TLTraceBuffer.scala 33:39]
  wire  _out_b_scan_bits_T = tl_out_b_ready & auto_out_b_valid; // @[Decoupled.scala 51:35]
  reg [2:0] out_b_scan_bits_size; // @[Reg.scala 35:20]
  reg [3:0] out_b_scan_bits_source; // @[Reg.scala 35:20]
  reg [31:0] out_b_scan_bits_address; // @[Reg.scala 35:20]
  wire  _GEN_18 = _x1_b_ready_T_1 ? 1'h0 : out_b_scan_valid; // @[Utils.scala 38:18 36:20 38:22]
  wire  _GEN_19 = _out_b_scan_bits_T | _GEN_18; // @[Utils.scala 39:{19,23}]
  reg  in_c_scan_valid; // @[Utils.scala 36:20]
  wire  _x1_c_ready_T_1 = auto_out_c_ready & in_c_scan_valid; // @[Decoupled.scala 51:35]
  wire  tl_in_c_ready = ~in_c_scan_valid | _x1_c_ready_T_1; // @[TLTraceBuffer.scala 36:38]
  wire  _in_c_scan_bits_T = tl_in_c_ready & auto_in_c_valid; // @[Decoupled.scala 51:35]
  reg [2:0] in_c_scan_bits_opcode; // @[Reg.scala 35:20]
  reg [2:0] in_c_scan_bits_param; // @[Reg.scala 35:20]
  reg [2:0] in_c_scan_bits_size; // @[Reg.scala 35:20]
  reg [3:0] in_c_scan_bits_source; // @[Reg.scala 35:20]
  reg [31:0] in_c_scan_bits_address; // @[Reg.scala 35:20]
  reg [255:0] in_c_scan_bits_data; // @[Reg.scala 35:20]
  wire  _GEN_27 = _x1_c_ready_T_1 ? 1'h0 : in_c_scan_valid; // @[Utils.scala 38:18 36:20 38:22]
  wire  _GEN_28 = _in_c_scan_bits_T | _GEN_27; // @[Utils.scala 39:{19,23}]
  reg  out_d_scan_valid; // @[Utils.scala 36:20]
  wire  _x1_d_ready_T_1 = auto_in_d_ready & out_d_scan_valid; // @[Decoupled.scala 51:35]
  wire  tl_out_d_ready = ~out_d_scan_valid | _x1_d_ready_T_1; // @[TLTraceBuffer.scala 39:39]
  wire  _out_d_scan_bits_T = tl_out_d_ready & auto_out_d_valid; // @[Decoupled.scala 51:35]
  reg [2:0] out_d_scan_bits_opcode; // @[Reg.scala 35:20]
  reg [2:0] out_d_scan_bits_size; // @[Reg.scala 35:20]
  reg [3:0] out_d_scan_bits_source; // @[Reg.scala 35:20]
  reg [5:0] out_d_scan_bits_sink; // @[Reg.scala 35:20]
  reg [255:0] out_d_scan_bits_data; // @[Reg.scala 35:20]
  wire  _GEN_37 = _x1_d_ready_T_1 ? 1'h0 : out_d_scan_valid; // @[Utils.scala 38:18 36:20 38:22]
  wire  _GEN_38 = _out_d_scan_bits_T | _GEN_37; // @[Utils.scala 39:{19,23}]
  reg  in_e_scan_valid; // @[Utils.scala 36:20]
  wire  _x1_e_ready_T_1 = auto_out_e_ready & in_e_scan_valid; // @[Decoupled.scala 51:35]
  wire  tl_in_e_ready = ~in_e_scan_valid | _x1_e_ready_T_1; // @[TLTraceBuffer.scala 42:38]
  wire  _in_e_scan_bits_T = tl_in_e_ready & auto_in_e_valid; // @[Decoupled.scala 51:35]
  reg [5:0] in_e_scan_bits_sink; // @[Reg.scala 35:20]
  wire  _GEN_40 = _x1_e_ready_T_1 ? 1'h0 : in_e_scan_valid; // @[Utils.scala 38:18 36:20 38:22]
  wire  _GEN_41 = _in_e_scan_bits_T | _GEN_40; // @[Utils.scala 39:{19,23}]
  assign auto_in_a_ready = ~in_a_scan_valid | _x1_a_ready_T_1; // @[TLTraceBuffer.scala 30:38]
  assign auto_in_b_valid = out_b_scan_valid; // @[Nodes.scala 1215:84 TLTraceBuffer.scala 31:18]
  assign auto_in_b_bits_size = out_b_scan_bits_size; // @[Nodes.scala 1215:84 TLTraceBuffer.scala 32:18]
  assign auto_in_b_bits_source = out_b_scan_bits_source; // @[Nodes.scala 1215:84 TLTraceBuffer.scala 32:18]
  assign auto_in_b_bits_address = out_b_scan_bits_address; // @[Nodes.scala 1215:84 TLTraceBuffer.scala 32:18]
  assign auto_in_c_ready = ~in_c_scan_valid | _x1_c_ready_T_1; // @[TLTraceBuffer.scala 36:38]
  assign auto_in_d_valid = out_d_scan_valid; // @[Nodes.scala 1215:84 TLTraceBuffer.scala 37:18]
  assign auto_in_d_bits_opcode = out_d_scan_bits_opcode; // @[Nodes.scala 1215:84 TLTraceBuffer.scala 38:18]
  assign auto_in_d_bits_size = out_d_scan_bits_size; // @[Nodes.scala 1215:84 TLTraceBuffer.scala 38:18]
  assign auto_in_d_bits_source = out_d_scan_bits_source; // @[Nodes.scala 1215:84 TLTraceBuffer.scala 38:18]
  assign auto_in_d_bits_sink = out_d_scan_bits_sink; // @[Nodes.scala 1215:84 TLTraceBuffer.scala 38:18]
  assign auto_in_d_bits_data = out_d_scan_bits_data; // @[Nodes.scala 1215:84 TLTraceBuffer.scala 38:18]
  assign auto_in_e_ready = ~in_e_scan_valid | _x1_e_ready_T_1; // @[TLTraceBuffer.scala 42:38]
  assign auto_out_a_valid = in_a_scan_valid; // @[Nodes.scala 1212:84 TLTraceBuffer.scala 28:18]
  assign auto_out_a_bits_opcode = in_a_scan_bits_opcode; // @[Nodes.scala 1212:84 TLTraceBuffer.scala 29:18]
  assign auto_out_a_bits_param = in_a_scan_bits_param; // @[Nodes.scala 1212:84 TLTraceBuffer.scala 29:18]
  assign auto_out_a_bits_size = in_a_scan_bits_size; // @[Nodes.scala 1212:84 TLTraceBuffer.scala 29:18]
  assign auto_out_a_bits_source = in_a_scan_bits_source; // @[Nodes.scala 1212:84 TLTraceBuffer.scala 29:18]
  assign auto_out_a_bits_address = in_a_scan_bits_address; // @[Nodes.scala 1212:84 TLTraceBuffer.scala 29:18]
  assign auto_out_a_bits_mask = in_a_scan_bits_mask; // @[Nodes.scala 1212:84 TLTraceBuffer.scala 29:18]
  assign auto_out_a_bits_data = in_a_scan_bits_data; // @[Nodes.scala 1212:84 TLTraceBuffer.scala 29:18]
  assign auto_out_b_ready = ~out_b_scan_valid | _x1_b_ready_T_1; // @[TLTraceBuffer.scala 33:39]
  assign auto_out_c_valid = in_c_scan_valid; // @[Nodes.scala 1212:84 TLTraceBuffer.scala 34:18]
  assign auto_out_c_bits_opcode = in_c_scan_bits_opcode; // @[Nodes.scala 1212:84 TLTraceBuffer.scala 35:18]
  assign auto_out_c_bits_param = in_c_scan_bits_param; // @[Nodes.scala 1212:84 TLTraceBuffer.scala 35:18]
  assign auto_out_c_bits_size = in_c_scan_bits_size; // @[Nodes.scala 1212:84 TLTraceBuffer.scala 35:18]
  assign auto_out_c_bits_source = in_c_scan_bits_source; // @[Nodes.scala 1212:84 TLTraceBuffer.scala 35:18]
  assign auto_out_c_bits_address = in_c_scan_bits_address; // @[Nodes.scala 1212:84 TLTraceBuffer.scala 35:18]
  assign auto_out_c_bits_data = in_c_scan_bits_data; // @[Nodes.scala 1212:84 TLTraceBuffer.scala 35:18]
  assign auto_out_d_ready = ~out_d_scan_valid | _x1_d_ready_T_1; // @[TLTraceBuffer.scala 39:39]
  assign auto_out_e_valid = in_e_scan_valid; // @[Nodes.scala 1212:84 TLTraceBuffer.scala 40:18]
  assign auto_out_e_bits_sink = in_e_scan_bits_sink; // @[Nodes.scala 1212:84 TLTraceBuffer.scala 41:18]
  always @(posedge clock) begin
    if (reset) begin // @[Utils.scala 36:20]
      in_a_scan_valid <= 1'h0; // @[Utils.scala 36:20]
    end else begin
      in_a_scan_valid <= _GEN_9;
    end
    if (reset) begin // @[Reg.scala 35:20]
      in_a_scan_bits_opcode <= 3'h0; // @[Reg.scala 35:20]
    end else if (_in_a_scan_bits_T) begin // @[Reg.scala 36:18]
      in_a_scan_bits_opcode <= auto_in_a_bits_opcode; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      in_a_scan_bits_param <= 3'h0; // @[Reg.scala 35:20]
    end else if (_in_a_scan_bits_T) begin // @[Reg.scala 36:18]
      in_a_scan_bits_param <= auto_in_a_bits_param; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      in_a_scan_bits_size <= 3'h0; // @[Reg.scala 35:20]
    end else if (_in_a_scan_bits_T) begin // @[Reg.scala 36:18]
      in_a_scan_bits_size <= auto_in_a_bits_size; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      in_a_scan_bits_source <= 4'h0; // @[Reg.scala 35:20]
    end else if (_in_a_scan_bits_T) begin // @[Reg.scala 36:18]
      in_a_scan_bits_source <= auto_in_a_bits_source; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      in_a_scan_bits_address <= 32'h0; // @[Reg.scala 35:20]
    end else if (_in_a_scan_bits_T) begin // @[Reg.scala 36:18]
      in_a_scan_bits_address <= auto_in_a_bits_address; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      in_a_scan_bits_mask <= 32'h0; // @[Reg.scala 35:20]
    end else if (_in_a_scan_bits_T) begin // @[Reg.scala 36:18]
      in_a_scan_bits_mask <= auto_in_a_bits_mask; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      in_a_scan_bits_data <= 256'h0; // @[Reg.scala 35:20]
    end else if (_in_a_scan_bits_T) begin // @[Reg.scala 36:18]
      in_a_scan_bits_data <= auto_in_a_bits_data; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Utils.scala 36:20]
      out_b_scan_valid <= 1'h0; // @[Utils.scala 36:20]
    end else begin
      out_b_scan_valid <= _GEN_19;
    end
    if (reset) begin // @[Reg.scala 35:20]
      out_b_scan_bits_size <= 3'h0; // @[Reg.scala 35:20]
    end else if (_out_b_scan_bits_T) begin // @[Reg.scala 36:18]
      out_b_scan_bits_size <= auto_out_b_bits_size; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      out_b_scan_bits_source <= 4'h0; // @[Reg.scala 35:20]
    end else if (_out_b_scan_bits_T) begin // @[Reg.scala 36:18]
      out_b_scan_bits_source <= auto_out_b_bits_source; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      out_b_scan_bits_address <= 32'h0; // @[Reg.scala 35:20]
    end else if (_out_b_scan_bits_T) begin // @[Reg.scala 36:18]
      out_b_scan_bits_address <= auto_out_b_bits_address; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Utils.scala 36:20]
      in_c_scan_valid <= 1'h0; // @[Utils.scala 36:20]
    end else begin
      in_c_scan_valid <= _GEN_28;
    end
    if (reset) begin // @[Reg.scala 35:20]
      in_c_scan_bits_opcode <= 3'h0; // @[Reg.scala 35:20]
    end else if (_in_c_scan_bits_T) begin // @[Reg.scala 36:18]
      in_c_scan_bits_opcode <= auto_in_c_bits_opcode; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      in_c_scan_bits_param <= 3'h0; // @[Reg.scala 35:20]
    end else if (_in_c_scan_bits_T) begin // @[Reg.scala 36:18]
      in_c_scan_bits_param <= auto_in_c_bits_param; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      in_c_scan_bits_size <= 3'h0; // @[Reg.scala 35:20]
    end else if (_in_c_scan_bits_T) begin // @[Reg.scala 36:18]
      in_c_scan_bits_size <= auto_in_c_bits_size; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      in_c_scan_bits_source <= 4'h0; // @[Reg.scala 35:20]
    end else if (_in_c_scan_bits_T) begin // @[Reg.scala 36:18]
      in_c_scan_bits_source <= auto_in_c_bits_source; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      in_c_scan_bits_address <= 32'h0; // @[Reg.scala 35:20]
    end else if (_in_c_scan_bits_T) begin // @[Reg.scala 36:18]
      in_c_scan_bits_address <= auto_in_c_bits_address; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      in_c_scan_bits_data <= 256'h0; // @[Reg.scala 35:20]
    end else if (_in_c_scan_bits_T) begin // @[Reg.scala 36:18]
      in_c_scan_bits_data <= auto_in_c_bits_data; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Utils.scala 36:20]
      out_d_scan_valid <= 1'h0; // @[Utils.scala 36:20]
    end else begin
      out_d_scan_valid <= _GEN_38;
    end
    if (reset) begin // @[Reg.scala 35:20]
      out_d_scan_bits_opcode <= 3'h0; // @[Reg.scala 35:20]
    end else if (_out_d_scan_bits_T) begin // @[Reg.scala 36:18]
      out_d_scan_bits_opcode <= auto_out_d_bits_opcode; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      out_d_scan_bits_size <= 3'h0; // @[Reg.scala 35:20]
    end else if (_out_d_scan_bits_T) begin // @[Reg.scala 36:18]
      out_d_scan_bits_size <= auto_out_d_bits_size; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      out_d_scan_bits_source <= 4'h0; // @[Reg.scala 35:20]
    end else if (_out_d_scan_bits_T) begin // @[Reg.scala 36:18]
      out_d_scan_bits_source <= auto_out_d_bits_source; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      out_d_scan_bits_sink <= 6'h0; // @[Reg.scala 35:20]
    end else if (_out_d_scan_bits_T) begin // @[Reg.scala 36:18]
      out_d_scan_bits_sink <= auto_out_d_bits_sink; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      out_d_scan_bits_data <= 256'h0; // @[Reg.scala 35:20]
    end else if (_out_d_scan_bits_T) begin // @[Reg.scala 36:18]
      out_d_scan_bits_data <= auto_out_d_bits_data; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Utils.scala 36:20]
      in_e_scan_valid <= 1'h0; // @[Utils.scala 36:20]
    end else begin
      in_e_scan_valid <= _GEN_41;
    end
    if (reset) begin // @[Reg.scala 35:20]
      in_e_scan_bits_sink <= 6'h0; // @[Reg.scala 35:20]
    end else if (_in_e_scan_bits_T) begin // @[Reg.scala 36:18]
      in_e_scan_bits_sink <= auto_in_e_bits_sink; // @[Reg.scala 36:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  in_a_scan_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  in_a_scan_bits_opcode = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  in_a_scan_bits_param = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  in_a_scan_bits_size = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  in_a_scan_bits_source = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  in_a_scan_bits_address = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  in_a_scan_bits_mask = _RAND_6[31:0];
  _RAND_7 = {8{`RANDOM}};
  in_a_scan_bits_data = _RAND_7[255:0];
  _RAND_8 = {1{`RANDOM}};
  out_b_scan_valid = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  out_b_scan_bits_size = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  out_b_scan_bits_source = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  out_b_scan_bits_address = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  in_c_scan_valid = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  in_c_scan_bits_opcode = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  in_c_scan_bits_param = _RAND_14[2:0];
  _RAND_15 = {1{`RANDOM}};
  in_c_scan_bits_size = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  in_c_scan_bits_source = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
  in_c_scan_bits_address = _RAND_17[31:0];
  _RAND_18 = {8{`RANDOM}};
  in_c_scan_bits_data = _RAND_18[255:0];
  _RAND_19 = {1{`RANDOM}};
  out_d_scan_valid = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  out_d_scan_bits_opcode = _RAND_20[2:0];
  _RAND_21 = {1{`RANDOM}};
  out_d_scan_bits_size = _RAND_21[2:0];
  _RAND_22 = {1{`RANDOM}};
  out_d_scan_bits_source = _RAND_22[3:0];
  _RAND_23 = {1{`RANDOM}};
  out_d_scan_bits_sink = _RAND_23[5:0];
  _RAND_24 = {8{`RANDOM}};
  out_d_scan_bits_data = _RAND_24[255:0];
  _RAND_25 = {1{`RANDOM}};
  in_e_scan_valid = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  in_e_scan_bits_sink = _RAND_26[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AsyncResetSynchronizerPrimitiveShiftReg_d3_i0(
  input   clock,
  input   reset,
  input   io_d,
  output  io_q
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg  sync_0; // @[SynchronizerReg.scala 51:87]
  reg  sync_1; // @[SynchronizerReg.scala 51:87]
  reg  sync_2; // @[SynchronizerReg.scala 51:87]
  assign io_q = sync_0; // @[SynchronizerReg.scala 59:8]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SynchronizerReg.scala 51:87]
      sync_0 <= 1'h0; // @[SynchronizerReg.scala 51:87]
    end else begin
      sync_0 <= sync_1; // @[SynchronizerReg.scala 57:10]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SynchronizerReg.scala 51:87]
      sync_1 <= 1'h0; // @[SynchronizerReg.scala 51:87]
    end else begin
      sync_1 <= sync_2; // @[SynchronizerReg.scala 57:10]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[SynchronizerReg.scala 54:22]
      sync_2 <= 1'h0;
    end else begin
      sync_2 <= io_d;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sync_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  sync_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  sync_2 = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    sync_0 = 1'h0;
  end
  if (reset) begin
    sync_1 = 1'h0;
  end
  if (reset) begin
    sync_2 = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AsyncResetSynchronizerShiftReg_w4_d3_i0(
  input        clock,
  input        reset,
  input  [3:0] io_d,
  output [3:0] io_q
);
  wire  output_chain_clock; // @[ShiftReg.scala 45:23]
  wire  output_chain_reset; // @[ShiftReg.scala 45:23]
  wire  output_chain_io_d; // @[ShiftReg.scala 45:23]
  wire  output_chain_io_q; // @[ShiftReg.scala 45:23]
  wire  output_chain_1_clock; // @[ShiftReg.scala 45:23]
  wire  output_chain_1_reset; // @[ShiftReg.scala 45:23]
  wire  output_chain_1_io_d; // @[ShiftReg.scala 45:23]
  wire  output_chain_1_io_q; // @[ShiftReg.scala 45:23]
  wire  output_chain_2_clock; // @[ShiftReg.scala 45:23]
  wire  output_chain_2_reset; // @[ShiftReg.scala 45:23]
  wire  output_chain_2_io_d; // @[ShiftReg.scala 45:23]
  wire  output_chain_2_io_q; // @[ShiftReg.scala 45:23]
  wire  output_chain_3_clock; // @[ShiftReg.scala 45:23]
  wire  output_chain_3_reset; // @[ShiftReg.scala 45:23]
  wire  output_chain_3_io_d; // @[ShiftReg.scala 45:23]
  wire  output_chain_3_io_q; // @[ShiftReg.scala 45:23]
  wire  output_1 = output_chain_1_io_q; // @[ShiftReg.scala 48:{24,24}]
  wire  output_0 = output_chain_io_q; // @[ShiftReg.scala 48:{24,24}]
  wire [1:0] io_q_lo = {output_1,output_0}; // @[Cat.scala 33:92]
  wire  output_3 = output_chain_3_io_q; // @[ShiftReg.scala 48:{24,24}]
  wire  output_2 = output_chain_2_io_q; // @[ShiftReg.scala 48:{24,24}]
  wire [1:0] io_q_hi = {output_3,output_2}; // @[Cat.scala 33:92]
  AsyncResetSynchronizerPrimitiveShiftReg_d3_i0 output_chain ( // @[ShiftReg.scala 45:23]
    .clock(output_chain_clock),
    .reset(output_chain_reset),
    .io_d(output_chain_io_d),
    .io_q(output_chain_io_q)
  );
  AsyncResetSynchronizerPrimitiveShiftReg_d3_i0 output_chain_1 ( // @[ShiftReg.scala 45:23]
    .clock(output_chain_1_clock),
    .reset(output_chain_1_reset),
    .io_d(output_chain_1_io_d),
    .io_q(output_chain_1_io_q)
  );
  AsyncResetSynchronizerPrimitiveShiftReg_d3_i0 output_chain_2 ( // @[ShiftReg.scala 45:23]
    .clock(output_chain_2_clock),
    .reset(output_chain_2_reset),
    .io_d(output_chain_2_io_d),
    .io_q(output_chain_2_io_q)
  );
  AsyncResetSynchronizerPrimitiveShiftReg_d3_i0 output_chain_3 ( // @[ShiftReg.scala 45:23]
    .clock(output_chain_3_clock),
    .reset(output_chain_3_reset),
    .io_d(output_chain_3_io_d),
    .io_q(output_chain_3_io_q)
  );
  assign io_q = {io_q_hi,io_q_lo}; // @[Cat.scala 33:92]
  assign output_chain_clock = clock;
  assign output_chain_reset = reset; // @[SynchronizerReg.scala 86:21]
  assign output_chain_io_d = io_d[0]; // @[SynchronizerReg.scala 87:41]
  assign output_chain_1_clock = clock;
  assign output_chain_1_reset = reset; // @[SynchronizerReg.scala 86:21]
  assign output_chain_1_io_d = io_d[1]; // @[SynchronizerReg.scala 87:41]
  assign output_chain_2_clock = clock;
  assign output_chain_2_reset = reset; // @[SynchronizerReg.scala 86:21]
  assign output_chain_2_io_d = io_d[2]; // @[SynchronizerReg.scala 87:41]
  assign output_chain_3_clock = clock;
  assign output_chain_3_reset = reset; // @[SynchronizerReg.scala 86:21]
  assign output_chain_3_io_d = io_d[3]; // @[SynchronizerReg.scala 87:41]
endmodule
module AsyncResetSynchronizerShiftReg_w1_d3_i0(
  input   clock,
  input   reset,
  input   io_d,
  output  io_q
);
  wire  output_chain_clock; // @[ShiftReg.scala 45:23]
  wire  output_chain_reset; // @[ShiftReg.scala 45:23]
  wire  output_chain_io_d; // @[ShiftReg.scala 45:23]
  wire  output_chain_io_q; // @[ShiftReg.scala 45:23]
  AsyncResetSynchronizerPrimitiveShiftReg_d3_i0 output_chain ( // @[ShiftReg.scala 45:23]
    .clock(output_chain_clock),
    .reset(output_chain_reset),
    .io_d(output_chain_io_d),
    .io_q(output_chain_io_q)
  );
  assign io_q = output_chain_io_q; // @[ShiftReg.scala 48:{24,24}]
  assign output_chain_clock = clock;
  assign output_chain_reset = reset; // @[SynchronizerReg.scala 86:21]
  assign output_chain_io_d = io_d; // @[SynchronizerReg.scala 87:41]
endmodule
module AsyncValidSync(
  input   io_in,
  output  io_out,
  input   clock,
  input   reset
);
  wire  io_out_source_valid_0_clock; // @[ShiftReg.scala 45:23]
  wire  io_out_source_valid_0_reset; // @[ShiftReg.scala 45:23]
  wire  io_out_source_valid_0_io_d; // @[ShiftReg.scala 45:23]
  wire  io_out_source_valid_0_io_q; // @[ShiftReg.scala 45:23]
  AsyncResetSynchronizerShiftReg_w1_d3_i0 io_out_source_valid_0 ( // @[ShiftReg.scala 45:23]
    .clock(io_out_source_valid_0_clock),
    .reset(io_out_source_valid_0_reset),
    .io_d(io_out_source_valid_0_io_d),
    .io_q(io_out_source_valid_0_io_q)
  );
  assign io_out = io_out_source_valid_0_io_q; // @[ShiftReg.scala 48:{24,24}]
  assign io_out_source_valid_0_clock = clock;
  assign io_out_source_valid_0_reset = reset;
  assign io_out_source_valid_0_io_d = io_in; // @[ShiftReg.scala 47:16]
endmodule
module AsyncQueueSource(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [7:0] io_enq_bits,
  output [7:0] io_async_mem_0,
  output [7:0] io_async_mem_1,
  output [7:0] io_async_mem_2,
  output [7:0] io_async_mem_3,
  output [7:0] io_async_mem_4,
  output [7:0] io_async_mem_5,
  output [7:0] io_async_mem_6,
  output [7:0] io_async_mem_7,
  input  [3:0] io_async_ridx,
  output [3:0] io_async_widx,
  input        io_async_safe_ridx_valid,
  output       io_async_safe_widx_valid,
  output       io_async_safe_source_reset_n,
  input        io_async_safe_sink_reset_n
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire  ridx_ridx_gray_clock; // @[ShiftReg.scala 45:23]
  wire  ridx_ridx_gray_reset; // @[ShiftReg.scala 45:23]
  wire [3:0] ridx_ridx_gray_io_d; // @[ShiftReg.scala 45:23]
  wire [3:0] ridx_ridx_gray_io_q; // @[ShiftReg.scala 45:23]
  wire  source_valid_0_io_in; // @[AsyncQueue.scala 100:32]
  wire  source_valid_0_io_out; // @[AsyncQueue.scala 100:32]
  wire  source_valid_0_clock; // @[AsyncQueue.scala 100:32]
  wire  source_valid_0_reset; // @[AsyncQueue.scala 100:32]
  wire  source_valid_1_io_in; // @[AsyncQueue.scala 101:32]
  wire  source_valid_1_io_out; // @[AsyncQueue.scala 101:32]
  wire  source_valid_1_clock; // @[AsyncQueue.scala 101:32]
  wire  source_valid_1_reset; // @[AsyncQueue.scala 101:32]
  wire  sink_extend_io_in; // @[AsyncQueue.scala 103:30]
  wire  sink_extend_io_out; // @[AsyncQueue.scala 103:30]
  wire  sink_extend_clock; // @[AsyncQueue.scala 103:30]
  wire  sink_extend_reset; // @[AsyncQueue.scala 103:30]
  wire  sink_valid_io_in; // @[AsyncQueue.scala 104:30]
  wire  sink_valid_io_out; // @[AsyncQueue.scala 104:30]
  wire  sink_valid_clock; // @[AsyncQueue.scala 104:30]
  wire  sink_valid_reset; // @[AsyncQueue.scala 104:30]
  reg [7:0] mem_0; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_1; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_2; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_3; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_4; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_5; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_6; // @[AsyncQueue.scala 80:16]
  reg [7:0] mem_7; // @[AsyncQueue.scala 80:16]
  wire  _widx_T_1 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 51:35]
  wire  sink_ready = sink_valid_io_out; // @[AsyncQueue.scala 120:16 79:28]
  wire  _widx_T_2 = ~sink_ready; // @[AsyncQueue.scala 81:79]
  reg [3:0] widx_widx_bin; // @[AsyncQueue.scala 52:25]
  wire [3:0] _GEN_16 = {{3'd0}, _widx_T_1}; // @[AsyncQueue.scala 53:43]
  wire [3:0] _widx_incremented_T_1 = widx_widx_bin + _GEN_16; // @[AsyncQueue.scala 53:43]
  wire [3:0] widx_incremented = _widx_T_2 ? 4'h0 : _widx_incremented_T_1; // @[AsyncQueue.scala 53:23]
  wire [3:0] _GEN_17 = {{1'd0}, widx_incremented[3:1]}; // @[AsyncQueue.scala 54:17]
  wire [3:0] widx = widx_incremented ^ _GEN_17; // @[AsyncQueue.scala 54:17]
  wire [3:0] ridx = ridx_ridx_gray_io_q; // @[ShiftReg.scala 48:{24,24}]
  wire [3:0] _ready_T = ridx ^ 4'hc; // @[AsyncQueue.scala 83:44]
  wire [2:0] _index_T_2 = {io_async_widx[3], 2'h0}; // @[AsyncQueue.scala 85:93]
  wire [2:0] index = io_async_widx[2:0] ^ _index_T_2; // @[AsyncQueue.scala 85:64]
  reg  ready_reg; // @[AsyncQueue.scala 88:56]
  reg [3:0] widx_gray; // @[AsyncQueue.scala 91:55]
  AsyncResetSynchronizerShiftReg_w4_d3_i0 ridx_ridx_gray ( // @[ShiftReg.scala 45:23]
    .clock(ridx_ridx_gray_clock),
    .reset(ridx_ridx_gray_reset),
    .io_d(ridx_ridx_gray_io_d),
    .io_q(ridx_ridx_gray_io_q)
  );
  AsyncValidSync source_valid_0 ( // @[AsyncQueue.scala 100:32]
    .io_in(source_valid_0_io_in),
    .io_out(source_valid_0_io_out),
    .clock(source_valid_0_clock),
    .reset(source_valid_0_reset)
  );
  AsyncValidSync source_valid_1 ( // @[AsyncQueue.scala 101:32]
    .io_in(source_valid_1_io_in),
    .io_out(source_valid_1_io_out),
    .clock(source_valid_1_clock),
    .reset(source_valid_1_reset)
  );
  AsyncValidSync sink_extend ( // @[AsyncQueue.scala 103:30]
    .io_in(sink_extend_io_in),
    .io_out(sink_extend_io_out),
    .clock(sink_extend_clock),
    .reset(sink_extend_reset)
  );
  AsyncValidSync sink_valid ( // @[AsyncQueue.scala 104:30]
    .io_in(sink_valid_io_in),
    .io_out(sink_valid_io_out),
    .clock(sink_valid_clock),
    .reset(sink_valid_reset)
  );
  assign io_enq_ready = ready_reg & sink_ready; // @[AsyncQueue.scala 89:29]
  assign io_async_mem_0 = mem_0; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_1 = mem_1; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_2 = mem_2; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_3 = mem_3; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_4 = mem_4; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_5 = mem_5; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_6 = mem_6; // @[AsyncQueue.scala 96:31]
  assign io_async_mem_7 = mem_7; // @[AsyncQueue.scala 96:31]
  assign io_async_widx = widx_gray; // @[AsyncQueue.scala 92:17]
  assign io_async_safe_widx_valid = source_valid_1_io_out; // @[AsyncQueue.scala 117:20]
  assign io_async_safe_source_reset_n = ~reset; // @[AsyncQueue.scala 121:27]
  assign ridx_ridx_gray_clock = clock;
  assign ridx_ridx_gray_reset = reset;
  assign ridx_ridx_gray_io_d = io_async_ridx; // @[ShiftReg.scala 47:16]
  assign source_valid_0_io_in = 1'h1; // @[AsyncQueue.scala 115:26]
  assign source_valid_0_clock = clock; // @[AsyncQueue.scala 110:26]
  assign source_valid_0_reset = reset | ~io_async_safe_sink_reset_n; // @[AsyncQueue.scala 105:65]
  assign source_valid_1_io_in = source_valid_0_io_out; // @[AsyncQueue.scala 116:26]
  assign source_valid_1_clock = clock; // @[AsyncQueue.scala 111:26]
  assign source_valid_1_reset = reset | ~io_async_safe_sink_reset_n; // @[AsyncQueue.scala 106:65]
  assign sink_extend_io_in = io_async_safe_ridx_valid; // @[AsyncQueue.scala 118:23]
  assign sink_extend_clock = clock; // @[AsyncQueue.scala 112:26]
  assign sink_extend_reset = reset | ~io_async_safe_sink_reset_n; // @[AsyncQueue.scala 107:65]
  assign sink_valid_io_in = sink_extend_io_out; // @[AsyncQueue.scala 119:22]
  assign sink_valid_clock = clock; // @[AsyncQueue.scala 113:26]
  assign sink_valid_reset = reset; // @[AsyncQueue.scala 108:35]
  always @(posedge clock) begin
    if (_widx_T_1) begin // @[AsyncQueue.scala 86:24]
      if (3'h0 == index) begin // @[AsyncQueue.scala 86:37]
        mem_0 <= io_enq_bits; // @[AsyncQueue.scala 86:37]
      end
    end
    if (_widx_T_1) begin // @[AsyncQueue.scala 86:24]
      if (3'h1 == index) begin // @[AsyncQueue.scala 86:37]
        mem_1 <= io_enq_bits; // @[AsyncQueue.scala 86:37]
      end
    end
    if (_widx_T_1) begin // @[AsyncQueue.scala 86:24]
      if (3'h2 == index) begin // @[AsyncQueue.scala 86:37]
        mem_2 <= io_enq_bits; // @[AsyncQueue.scala 86:37]
      end
    end
    if (_widx_T_1) begin // @[AsyncQueue.scala 86:24]
      if (3'h3 == index) begin // @[AsyncQueue.scala 86:37]
        mem_3 <= io_enq_bits; // @[AsyncQueue.scala 86:37]
      end
    end
    if (_widx_T_1) begin // @[AsyncQueue.scala 86:24]
      if (3'h4 == index) begin // @[AsyncQueue.scala 86:37]
        mem_4 <= io_enq_bits; // @[AsyncQueue.scala 86:37]
      end
    end
    if (_widx_T_1) begin // @[AsyncQueue.scala 86:24]
      if (3'h5 == index) begin // @[AsyncQueue.scala 86:37]
        mem_5 <= io_enq_bits; // @[AsyncQueue.scala 86:37]
      end
    end
    if (_widx_T_1) begin // @[AsyncQueue.scala 86:24]
      if (3'h6 == index) begin // @[AsyncQueue.scala 86:37]
        mem_6 <= io_enq_bits; // @[AsyncQueue.scala 86:37]
      end
    end
    if (_widx_T_1) begin // @[AsyncQueue.scala 86:24]
      if (3'h7 == index) begin // @[AsyncQueue.scala 86:37]
        mem_7 <= io_enq_bits; // @[AsyncQueue.scala 86:37]
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsyncQueue.scala 53:23]
      widx_widx_bin <= 4'h0;
    end else if (_widx_T_2) begin
      widx_widx_bin <= 4'h0;
    end else begin
      widx_widx_bin <= _widx_incremented_T_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsyncQueue.scala 83:26]
      ready_reg <= 1'h0;
    end else begin
      ready_reg <= sink_ready & widx != _ready_T;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsyncQueue.scala 54:17]
      widx_gray <= 4'h0;
    end else begin
      widx_gray <= widx_incremented ^ _GEN_17;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mem_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  mem_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  mem_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  mem_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  mem_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  mem_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  mem_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  mem_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  widx_widx_bin = _RAND_8[3:0];
  _RAND_9 = {1{`RANDOM}};
  ready_reg = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  widx_gray = _RAND_10[3:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    widx_widx_bin = 4'h0;
  end
  if (reset) begin
    ready_reg = 1'h0;
  end
  if (reset) begin
    widx_gray = 4'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ClockCrossingReg_w8(
  input        clock,
  input  [7:0] io_d,
  output [7:0] io_q,
  input        io_en
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] cdc_reg; // @[Reg.scala 19:16]
  assign io_q = cdc_reg; // @[SynchronizerReg.scala 202:8]
  always @(posedge clock) begin
    if (io_en) begin // @[Reg.scala 20:18]
      cdc_reg <= io_d; // @[Reg.scala 20:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cdc_reg = _RAND_0[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AsyncQueueSink(
  input        clock,
  input        reset,
  input        io_deq_ready,
  output       io_deq_valid,
  output [7:0] io_deq_bits,
  input  [7:0] io_async_mem_0,
  input  [7:0] io_async_mem_1,
  input  [7:0] io_async_mem_2,
  input  [7:0] io_async_mem_3,
  input  [7:0] io_async_mem_4,
  input  [7:0] io_async_mem_5,
  input  [7:0] io_async_mem_6,
  input  [7:0] io_async_mem_7,
  output [3:0] io_async_ridx,
  input  [3:0] io_async_widx,
  output       io_async_safe_ridx_valid,
  input        io_async_safe_widx_valid,
  input        io_async_safe_source_reset_n,
  output       io_async_safe_sink_reset_n
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  widx_widx_gray_clock; // @[ShiftReg.scala 45:23]
  wire  widx_widx_gray_reset; // @[ShiftReg.scala 45:23]
  wire [3:0] widx_widx_gray_io_d; // @[ShiftReg.scala 45:23]
  wire [3:0] widx_widx_gray_io_q; // @[ShiftReg.scala 45:23]
  wire  io_deq_bits_deq_bits_reg_clock; // @[SynchronizerReg.scala 207:25]
  wire [7:0] io_deq_bits_deq_bits_reg_io_d; // @[SynchronizerReg.scala 207:25]
  wire [7:0] io_deq_bits_deq_bits_reg_io_q; // @[SynchronizerReg.scala 207:25]
  wire  io_deq_bits_deq_bits_reg_io_en; // @[SynchronizerReg.scala 207:25]
  wire  sink_valid_0_io_in; // @[AsyncQueue.scala 168:33]
  wire  sink_valid_0_io_out; // @[AsyncQueue.scala 168:33]
  wire  sink_valid_0_clock; // @[AsyncQueue.scala 168:33]
  wire  sink_valid_0_reset; // @[AsyncQueue.scala 168:33]
  wire  sink_valid_1_io_in; // @[AsyncQueue.scala 169:33]
  wire  sink_valid_1_io_out; // @[AsyncQueue.scala 169:33]
  wire  sink_valid_1_clock; // @[AsyncQueue.scala 169:33]
  wire  sink_valid_1_reset; // @[AsyncQueue.scala 169:33]
  wire  source_extend_io_in; // @[AsyncQueue.scala 171:31]
  wire  source_extend_io_out; // @[AsyncQueue.scala 171:31]
  wire  source_extend_clock; // @[AsyncQueue.scala 171:31]
  wire  source_extend_reset; // @[AsyncQueue.scala 171:31]
  wire  source_valid_io_in; // @[AsyncQueue.scala 172:31]
  wire  source_valid_io_out; // @[AsyncQueue.scala 172:31]
  wire  source_valid_clock; // @[AsyncQueue.scala 172:31]
  wire  source_valid_reset; // @[AsyncQueue.scala 172:31]
  wire  _ridx_T_1 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 51:35]
  wire  source_ready = source_valid_io_out; // @[AsyncQueue.scala 143:30 188:18]
  wire  _ridx_T_2 = ~source_ready; // @[AsyncQueue.scala 144:79]
  reg [3:0] ridx_ridx_bin; // @[AsyncQueue.scala 52:25]
  wire [3:0] _GEN_8 = {{3'd0}, _ridx_T_1}; // @[AsyncQueue.scala 53:43]
  wire [3:0] _ridx_incremented_T_1 = ridx_ridx_bin + _GEN_8; // @[AsyncQueue.scala 53:43]
  wire [3:0] ridx_incremented = _ridx_T_2 ? 4'h0 : _ridx_incremented_T_1; // @[AsyncQueue.scala 53:23]
  wire [3:0] _GEN_9 = {{1'd0}, ridx_incremented[3:1]}; // @[AsyncQueue.scala 54:17]
  wire [3:0] ridx = ridx_incremented ^ _GEN_9; // @[AsyncQueue.scala 54:17]
  wire [3:0] widx = widx_widx_gray_io_q; // @[ShiftReg.scala 48:{24,24}]
  wire [2:0] _index_T_2 = {ridx[3], 2'h0}; // @[AsyncQueue.scala 152:75]
  wire [2:0] index = ridx[2:0] ^ _index_T_2; // @[AsyncQueue.scala 152:55]
  wire [7:0] _GEN_1 = 3'h1 == index ? io_async_mem_1 : io_async_mem_0; // @[SynchronizerReg.scala 209:{18,18}]
  wire [7:0] _GEN_2 = 3'h2 == index ? io_async_mem_2 : _GEN_1; // @[SynchronizerReg.scala 209:{18,18}]
  wire [7:0] _GEN_3 = 3'h3 == index ? io_async_mem_3 : _GEN_2; // @[SynchronizerReg.scala 209:{18,18}]
  wire [7:0] _GEN_4 = 3'h4 == index ? io_async_mem_4 : _GEN_3; // @[SynchronizerReg.scala 209:{18,18}]
  wire [7:0] _GEN_5 = 3'h5 == index ? io_async_mem_5 : _GEN_4; // @[SynchronizerReg.scala 209:{18,18}]
  wire [7:0] _GEN_6 = 3'h6 == index ? io_async_mem_6 : _GEN_5; // @[SynchronizerReg.scala 209:{18,18}]
  reg  valid_reg; // @[AsyncQueue.scala 161:56]
  reg [3:0] ridx_gray; // @[AsyncQueue.scala 164:55]
  AsyncResetSynchronizerShiftReg_w4_d3_i0 widx_widx_gray ( // @[ShiftReg.scala 45:23]
    .clock(widx_widx_gray_clock),
    .reset(widx_widx_gray_reset),
    .io_d(widx_widx_gray_io_d),
    .io_q(widx_widx_gray_io_q)
  );
  ClockCrossingReg_w8 io_deq_bits_deq_bits_reg ( // @[SynchronizerReg.scala 207:25]
    .clock(io_deq_bits_deq_bits_reg_clock),
    .io_d(io_deq_bits_deq_bits_reg_io_d),
    .io_q(io_deq_bits_deq_bits_reg_io_q),
    .io_en(io_deq_bits_deq_bits_reg_io_en)
  );
  AsyncValidSync sink_valid_0 ( // @[AsyncQueue.scala 168:33]
    .io_in(sink_valid_0_io_in),
    .io_out(sink_valid_0_io_out),
    .clock(sink_valid_0_clock),
    .reset(sink_valid_0_reset)
  );
  AsyncValidSync sink_valid_1 ( // @[AsyncQueue.scala 169:33]
    .io_in(sink_valid_1_io_in),
    .io_out(sink_valid_1_io_out),
    .clock(sink_valid_1_clock),
    .reset(sink_valid_1_reset)
  );
  AsyncValidSync source_extend ( // @[AsyncQueue.scala 171:31]
    .io_in(source_extend_io_in),
    .io_out(source_extend_io_out),
    .clock(source_extend_clock),
    .reset(source_extend_reset)
  );
  AsyncValidSync source_valid ( // @[AsyncQueue.scala 172:31]
    .io_in(source_valid_io_in),
    .io_out(source_valid_io_out),
    .clock(source_valid_clock),
    .reset(source_valid_reset)
  );
  assign io_deq_valid = valid_reg & source_ready; // @[AsyncQueue.scala 162:29]
  assign io_deq_bits = io_deq_bits_deq_bits_reg_io_q; // @[SynchronizerReg.scala 211:{26,26}]
  assign io_async_ridx = ridx_gray; // @[AsyncQueue.scala 165:17]
  assign io_async_safe_ridx_valid = sink_valid_1_io_out; // @[AsyncQueue.scala 185:20]
  assign io_async_safe_sink_reset_n = ~reset; // @[AsyncQueue.scala 189:25]
  assign widx_widx_gray_clock = clock;
  assign widx_widx_gray_reset = reset;
  assign widx_widx_gray_io_d = io_async_widx; // @[ShiftReg.scala 47:16]
  assign io_deq_bits_deq_bits_reg_clock = clock;
  assign io_deq_bits_deq_bits_reg_io_d = 3'h7 == index ? io_async_mem_7 : _GEN_6; // @[SynchronizerReg.scala 209:{18,18}]
  assign io_deq_bits_deq_bits_reg_io_en = source_ready & ridx != widx; // @[AsyncQueue.scala 146:28]
  assign sink_valid_0_io_in = 1'h1; // @[AsyncQueue.scala 183:24]
  assign sink_valid_0_clock = clock; // @[AsyncQueue.scala 178:25]
  assign sink_valid_0_reset = reset | ~io_async_safe_source_reset_n; // @[AsyncQueue.scala 173:66]
  assign sink_valid_1_io_in = sink_valid_0_io_out; // @[AsyncQueue.scala 184:24]
  assign sink_valid_1_clock = clock; // @[AsyncQueue.scala 179:25]
  assign sink_valid_1_reset = reset | ~io_async_safe_source_reset_n; // @[AsyncQueue.scala 174:66]
  assign source_extend_io_in = io_async_safe_widx_valid; // @[AsyncQueue.scala 186:25]
  assign source_extend_clock = clock; // @[AsyncQueue.scala 180:25]
  assign source_extend_reset = reset | ~io_async_safe_source_reset_n; // @[AsyncQueue.scala 175:66]
  assign source_valid_io_in = source_extend_io_out; // @[AsyncQueue.scala 187:24]
  assign source_valid_clock = clock; // @[AsyncQueue.scala 181:25]
  assign source_valid_reset = reset; // @[AsyncQueue.scala 176:34]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsyncQueue.scala 53:23]
      ridx_ridx_bin <= 4'h0;
    end else if (_ridx_T_2) begin
      ridx_ridx_bin <= 4'h0;
    end else begin
      ridx_ridx_bin <= _ridx_incremented_T_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsyncQueue.scala 146:28]
      valid_reg <= 1'h0;
    end else begin
      valid_reg <= source_ready & ridx != widx;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsyncQueue.scala 54:17]
      ridx_gray <= 4'h0;
    end else begin
      ridx_gray <= ridx_incremented ^ _GEN_9;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ridx_ridx_bin = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  valid_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  ridx_gray = _RAND_2[3:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    ridx_ridx_bin = 4'h0;
  end
  if (reset) begin
    valid_reg = 1'h0;
  end
  if (reset) begin
    ridx_gray = 4'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AsyncQueue(
  input        io_enq_clock,
  input        io_enq_reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [7:0] io_enq_bits,
  input        io_deq_clock,
  input        io_deq_reset,
  input        io_deq_ready,
  output       io_deq_valid,
  output [7:0] io_deq_bits
);
  wire  source_clock; // @[AsyncQueue.scala 224:22]
  wire  source_reset; // @[AsyncQueue.scala 224:22]
  wire  source_io_enq_ready; // @[AsyncQueue.scala 224:22]
  wire  source_io_enq_valid; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_enq_bits; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_0; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_1; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_2; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_3; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_4; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_5; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_6; // @[AsyncQueue.scala 224:22]
  wire [7:0] source_io_async_mem_7; // @[AsyncQueue.scala 224:22]
  wire [3:0] source_io_async_ridx; // @[AsyncQueue.scala 224:22]
  wire [3:0] source_io_async_widx; // @[AsyncQueue.scala 224:22]
  wire  source_io_async_safe_ridx_valid; // @[AsyncQueue.scala 224:22]
  wire  source_io_async_safe_widx_valid; // @[AsyncQueue.scala 224:22]
  wire  source_io_async_safe_source_reset_n; // @[AsyncQueue.scala 224:22]
  wire  source_io_async_safe_sink_reset_n; // @[AsyncQueue.scala 224:22]
  wire  sink_clock; // @[AsyncQueue.scala 225:22]
  wire  sink_reset; // @[AsyncQueue.scala 225:22]
  wire  sink_io_deq_ready; // @[AsyncQueue.scala 225:22]
  wire  sink_io_deq_valid; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_deq_bits; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_0; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_1; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_2; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_3; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_4; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_5; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_6; // @[AsyncQueue.scala 225:22]
  wire [7:0] sink_io_async_mem_7; // @[AsyncQueue.scala 225:22]
  wire [3:0] sink_io_async_ridx; // @[AsyncQueue.scala 225:22]
  wire [3:0] sink_io_async_widx; // @[AsyncQueue.scala 225:22]
  wire  sink_io_async_safe_ridx_valid; // @[AsyncQueue.scala 225:22]
  wire  sink_io_async_safe_widx_valid; // @[AsyncQueue.scala 225:22]
  wire  sink_io_async_safe_source_reset_n; // @[AsyncQueue.scala 225:22]
  wire  sink_io_async_safe_sink_reset_n; // @[AsyncQueue.scala 225:22]
  AsyncQueueSource source ( // @[AsyncQueue.scala 224:22]
    .clock(source_clock),
    .reset(source_reset),
    .io_enq_ready(source_io_enq_ready),
    .io_enq_valid(source_io_enq_valid),
    .io_enq_bits(source_io_enq_bits),
    .io_async_mem_0(source_io_async_mem_0),
    .io_async_mem_1(source_io_async_mem_1),
    .io_async_mem_2(source_io_async_mem_2),
    .io_async_mem_3(source_io_async_mem_3),
    .io_async_mem_4(source_io_async_mem_4),
    .io_async_mem_5(source_io_async_mem_5),
    .io_async_mem_6(source_io_async_mem_6),
    .io_async_mem_7(source_io_async_mem_7),
    .io_async_ridx(source_io_async_ridx),
    .io_async_widx(source_io_async_widx),
    .io_async_safe_ridx_valid(source_io_async_safe_ridx_valid),
    .io_async_safe_widx_valid(source_io_async_safe_widx_valid),
    .io_async_safe_source_reset_n(source_io_async_safe_source_reset_n),
    .io_async_safe_sink_reset_n(source_io_async_safe_sink_reset_n)
  );
  AsyncQueueSink sink ( // @[AsyncQueue.scala 225:22]
    .clock(sink_clock),
    .reset(sink_reset),
    .io_deq_ready(sink_io_deq_ready),
    .io_deq_valid(sink_io_deq_valid),
    .io_deq_bits(sink_io_deq_bits),
    .io_async_mem_0(sink_io_async_mem_0),
    .io_async_mem_1(sink_io_async_mem_1),
    .io_async_mem_2(sink_io_async_mem_2),
    .io_async_mem_3(sink_io_async_mem_3),
    .io_async_mem_4(sink_io_async_mem_4),
    .io_async_mem_5(sink_io_async_mem_5),
    .io_async_mem_6(sink_io_async_mem_6),
    .io_async_mem_7(sink_io_async_mem_7),
    .io_async_ridx(sink_io_async_ridx),
    .io_async_widx(sink_io_async_widx),
    .io_async_safe_ridx_valid(sink_io_async_safe_ridx_valid),
    .io_async_safe_widx_valid(sink_io_async_safe_widx_valid),
    .io_async_safe_source_reset_n(sink_io_async_safe_source_reset_n),
    .io_async_safe_sink_reset_n(sink_io_async_safe_sink_reset_n)
  );
  assign io_enq_ready = source_io_enq_ready; // @[AsyncQueue.scala 232:17]
  assign io_deq_valid = sink_io_deq_valid; // @[AsyncQueue.scala 233:10]
  assign io_deq_bits = sink_io_deq_bits; // @[AsyncQueue.scala 233:10]
  assign source_clock = io_enq_clock; // @[AsyncQueue.scala 227:16]
  assign source_reset = io_enq_reset; // @[AsyncQueue.scala 228:16]
  assign source_io_enq_valid = io_enq_valid; // @[AsyncQueue.scala 232:17]
  assign source_io_enq_bits = io_enq_bits; // @[AsyncQueue.scala 232:17]
  assign source_io_async_ridx = sink_io_async_ridx; // @[AsyncQueue.scala 234:17]
  assign source_io_async_safe_ridx_valid = sink_io_async_safe_ridx_valid; // @[AsyncQueue.scala 234:17]
  assign source_io_async_safe_sink_reset_n = sink_io_async_safe_sink_reset_n; // @[AsyncQueue.scala 234:17]
  assign sink_clock = io_deq_clock; // @[AsyncQueue.scala 229:14]
  assign sink_reset = io_deq_reset; // @[AsyncQueue.scala 230:14]
  assign sink_io_deq_ready = io_deq_ready; // @[AsyncQueue.scala 233:10]
  assign sink_io_async_mem_0 = source_io_async_mem_0; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_1 = source_io_async_mem_1; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_2 = source_io_async_mem_2; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_3 = source_io_async_mem_3; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_4 = source_io_async_mem_4; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_5 = source_io_async_mem_5; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_6 = source_io_async_mem_6; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_mem_7 = source_io_async_mem_7; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_widx = source_io_async_widx; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_safe_widx_valid = source_io_async_safe_widx_valid; // @[AsyncQueue.scala 234:17]
  assign sink_io_async_safe_source_reset_n = source_io_async_safe_source_reset_n; // @[AsyncQueue.scala 234:17]
endmodule
module SoC(
  input        clock,
  input        reset,
  output       io_in_ready,
  input        io_in_valid,
  input  [7:0] io_in_bits,
  input        io_out_ready,
  output       io_out_valid,
  output [7:0] io_out_bits,
  input        io_io_clock,
  input        io_io_reset,
  input        io_intr_mtip,
  input        io_intr_msip,
  input        io_intr_meip,
  input        io_intr_seip
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  wire  soc_imp_clock; // @[SoC.scala 81:27]
  wire  soc_imp_reset; // @[SoC.scala 81:27]
  wire  soc_imp_auto_out_a_ready; // @[SoC.scala 81:27]
  wire  soc_imp_auto_out_a_valid; // @[SoC.scala 81:27]
  wire [2:0] soc_imp_auto_out_a_bits_opcode; // @[SoC.scala 81:27]
  wire [2:0] soc_imp_auto_out_a_bits_param; // @[SoC.scala 81:27]
  wire [2:0] soc_imp_auto_out_a_bits_size; // @[SoC.scala 81:27]
  wire [3:0] soc_imp_auto_out_a_bits_source; // @[SoC.scala 81:27]
  wire [31:0] soc_imp_auto_out_a_bits_address; // @[SoC.scala 81:27]
  wire [31:0] soc_imp_auto_out_a_bits_mask; // @[SoC.scala 81:27]
  wire [255:0] soc_imp_auto_out_a_bits_data; // @[SoC.scala 81:27]
  wire  soc_imp_auto_out_b_ready; // @[SoC.scala 81:27]
  wire  soc_imp_auto_out_b_valid; // @[SoC.scala 81:27]
  wire [2:0] soc_imp_auto_out_b_bits_size; // @[SoC.scala 81:27]
  wire [3:0] soc_imp_auto_out_b_bits_source; // @[SoC.scala 81:27]
  wire [31:0] soc_imp_auto_out_b_bits_address; // @[SoC.scala 81:27]
  wire  soc_imp_auto_out_c_ready; // @[SoC.scala 81:27]
  wire  soc_imp_auto_out_c_valid; // @[SoC.scala 81:27]
  wire [2:0] soc_imp_auto_out_c_bits_opcode; // @[SoC.scala 81:27]
  wire [2:0] soc_imp_auto_out_c_bits_param; // @[SoC.scala 81:27]
  wire [2:0] soc_imp_auto_out_c_bits_size; // @[SoC.scala 81:27]
  wire [3:0] soc_imp_auto_out_c_bits_source; // @[SoC.scala 81:27]
  wire [31:0] soc_imp_auto_out_c_bits_address; // @[SoC.scala 81:27]
  wire [255:0] soc_imp_auto_out_c_bits_data; // @[SoC.scala 81:27]
  wire  soc_imp_auto_out_d_ready; // @[SoC.scala 81:27]
  wire  soc_imp_auto_out_d_valid; // @[SoC.scala 81:27]
  wire [2:0] soc_imp_auto_out_d_bits_opcode; // @[SoC.scala 81:27]
  wire [2:0] soc_imp_auto_out_d_bits_size; // @[SoC.scala 81:27]
  wire [3:0] soc_imp_auto_out_d_bits_source; // @[SoC.scala 81:27]
  wire [5:0] soc_imp_auto_out_d_bits_sink; // @[SoC.scala 81:27]
  wire [255:0] soc_imp_auto_out_d_bits_data; // @[SoC.scala 81:27]
  wire  soc_imp_auto_out_e_ready; // @[SoC.scala 81:27]
  wire  soc_imp_auto_out_e_valid; // @[SoC.scala 81:27]
  wire [5:0] soc_imp_auto_out_e_bits_sink; // @[SoC.scala 81:27]
  wire  soc_imp_io_intr_mtip; // @[SoC.scala 81:27]
  wire  soc_imp_io_intr_msip; // @[SoC.scala 81:27]
  wire  soc_imp_io_intr_meip; // @[SoC.scala 81:27]
  wire  soc_imp_io_intr_seip; // @[SoC.scala 81:27]
  wire  serdes_clock; // @[SoC.scala 87:26]
  wire  serdes_reset; // @[SoC.scala 87:26]
  wire  serdes_auto_in_a_ready; // @[SoC.scala 87:26]
  wire  serdes_auto_in_a_valid; // @[SoC.scala 87:26]
  wire [2:0] serdes_auto_in_a_bits_opcode; // @[SoC.scala 87:26]
  wire [2:0] serdes_auto_in_a_bits_param; // @[SoC.scala 87:26]
  wire [2:0] serdes_auto_in_a_bits_size; // @[SoC.scala 87:26]
  wire [3:0] serdes_auto_in_a_bits_source; // @[SoC.scala 87:26]
  wire [31:0] serdes_auto_in_a_bits_address; // @[SoC.scala 87:26]
  wire [31:0] serdes_auto_in_a_bits_mask; // @[SoC.scala 87:26]
  wire [255:0] serdes_auto_in_a_bits_data; // @[SoC.scala 87:26]
  wire  serdes_auto_in_b_ready; // @[SoC.scala 87:26]
  wire  serdes_auto_in_b_valid; // @[SoC.scala 87:26]
  wire [2:0] serdes_auto_in_b_bits_size; // @[SoC.scala 87:26]
  wire [3:0] serdes_auto_in_b_bits_source; // @[SoC.scala 87:26]
  wire [31:0] serdes_auto_in_b_bits_address; // @[SoC.scala 87:26]
  wire  serdes_auto_in_c_ready; // @[SoC.scala 87:26]
  wire  serdes_auto_in_c_valid; // @[SoC.scala 87:26]
  wire [2:0] serdes_auto_in_c_bits_opcode; // @[SoC.scala 87:26]
  wire [2:0] serdes_auto_in_c_bits_param; // @[SoC.scala 87:26]
  wire [2:0] serdes_auto_in_c_bits_size; // @[SoC.scala 87:26]
  wire [3:0] serdes_auto_in_c_bits_source; // @[SoC.scala 87:26]
  wire [31:0] serdes_auto_in_c_bits_address; // @[SoC.scala 87:26]
  wire [255:0] serdes_auto_in_c_bits_data; // @[SoC.scala 87:26]
  wire  serdes_auto_in_d_ready; // @[SoC.scala 87:26]
  wire  serdes_auto_in_d_valid; // @[SoC.scala 87:26]
  wire [2:0] serdes_auto_in_d_bits_opcode; // @[SoC.scala 87:26]
  wire [2:0] serdes_auto_in_d_bits_size; // @[SoC.scala 87:26]
  wire [3:0] serdes_auto_in_d_bits_source; // @[SoC.scala 87:26]
  wire [5:0] serdes_auto_in_d_bits_sink; // @[SoC.scala 87:26]
  wire [255:0] serdes_auto_in_d_bits_data; // @[SoC.scala 87:26]
  wire  serdes_auto_in_e_ready; // @[SoC.scala 87:26]
  wire  serdes_auto_in_e_valid; // @[SoC.scala 87:26]
  wire [5:0] serdes_auto_in_e_bits_sink; // @[SoC.scala 87:26]
  wire  serdes_io_ser_0_in_ready; // @[SoC.scala 87:26]
  wire  serdes_io_ser_0_in_valid; // @[SoC.scala 87:26]
  wire [7:0] serdes_io_ser_0_in_bits; // @[SoC.scala 87:26]
  wire  serdes_io_ser_0_out_ready; // @[SoC.scala 87:26]
  wire  serdes_io_ser_0_out_valid; // @[SoC.scala 87:26]
  wire [7:0] serdes_io_ser_0_out_bits; // @[SoC.scala 87:26]
  wire  trace_buffer_clock; // @[TLTraceBuffer.scala 47:34]
  wire  trace_buffer_reset; // @[TLTraceBuffer.scala 47:34]
  wire  trace_buffer_auto_in_a_ready; // @[TLTraceBuffer.scala 47:34]
  wire  trace_buffer_auto_in_a_valid; // @[TLTraceBuffer.scala 47:34]
  wire [2:0] trace_buffer_auto_in_a_bits_opcode; // @[TLTraceBuffer.scala 47:34]
  wire [2:0] trace_buffer_auto_in_a_bits_param; // @[TLTraceBuffer.scala 47:34]
  wire [2:0] trace_buffer_auto_in_a_bits_size; // @[TLTraceBuffer.scala 47:34]
  wire [3:0] trace_buffer_auto_in_a_bits_source; // @[TLTraceBuffer.scala 47:34]
  wire [31:0] trace_buffer_auto_in_a_bits_address; // @[TLTraceBuffer.scala 47:34]
  wire [31:0] trace_buffer_auto_in_a_bits_mask; // @[TLTraceBuffer.scala 47:34]
  wire [255:0] trace_buffer_auto_in_a_bits_data; // @[TLTraceBuffer.scala 47:34]
  wire  trace_buffer_auto_in_b_ready; // @[TLTraceBuffer.scala 47:34]
  wire  trace_buffer_auto_in_b_valid; // @[TLTraceBuffer.scala 47:34]
  wire [2:0] trace_buffer_auto_in_b_bits_size; // @[TLTraceBuffer.scala 47:34]
  wire [3:0] trace_buffer_auto_in_b_bits_source; // @[TLTraceBuffer.scala 47:34]
  wire [31:0] trace_buffer_auto_in_b_bits_address; // @[TLTraceBuffer.scala 47:34]
  wire  trace_buffer_auto_in_c_ready; // @[TLTraceBuffer.scala 47:34]
  wire  trace_buffer_auto_in_c_valid; // @[TLTraceBuffer.scala 47:34]
  wire [2:0] trace_buffer_auto_in_c_bits_opcode; // @[TLTraceBuffer.scala 47:34]
  wire [2:0] trace_buffer_auto_in_c_bits_param; // @[TLTraceBuffer.scala 47:34]
  wire [2:0] trace_buffer_auto_in_c_bits_size; // @[TLTraceBuffer.scala 47:34]
  wire [3:0] trace_buffer_auto_in_c_bits_source; // @[TLTraceBuffer.scala 47:34]
  wire [31:0] trace_buffer_auto_in_c_bits_address; // @[TLTraceBuffer.scala 47:34]
  wire [255:0] trace_buffer_auto_in_c_bits_data; // @[TLTraceBuffer.scala 47:34]
  wire  trace_buffer_auto_in_d_ready; // @[TLTraceBuffer.scala 47:34]
  wire  trace_buffer_auto_in_d_valid; // @[TLTraceBuffer.scala 47:34]
  wire [2:0] trace_buffer_auto_in_d_bits_opcode; // @[TLTraceBuffer.scala 47:34]
  wire [2:0] trace_buffer_auto_in_d_bits_size; // @[TLTraceBuffer.scala 47:34]
  wire [3:0] trace_buffer_auto_in_d_bits_source; // @[TLTraceBuffer.scala 47:34]
  wire [5:0] trace_buffer_auto_in_d_bits_sink; // @[TLTraceBuffer.scala 47:34]
  wire [255:0] trace_buffer_auto_in_d_bits_data; // @[TLTraceBuffer.scala 47:34]
  wire  trace_buffer_auto_in_e_ready; // @[TLTraceBuffer.scala 47:34]
  wire  trace_buffer_auto_in_e_valid; // @[TLTraceBuffer.scala 47:34]
  wire [5:0] trace_buffer_auto_in_e_bits_sink; // @[TLTraceBuffer.scala 47:34]
  wire  trace_buffer_auto_out_a_ready; // @[TLTraceBuffer.scala 47:34]
  wire  trace_buffer_auto_out_a_valid; // @[TLTraceBuffer.scala 47:34]
  wire [2:0] trace_buffer_auto_out_a_bits_opcode; // @[TLTraceBuffer.scala 47:34]
  wire [2:0] trace_buffer_auto_out_a_bits_param; // @[TLTraceBuffer.scala 47:34]
  wire [2:0] trace_buffer_auto_out_a_bits_size; // @[TLTraceBuffer.scala 47:34]
  wire [3:0] trace_buffer_auto_out_a_bits_source; // @[TLTraceBuffer.scala 47:34]
  wire [31:0] trace_buffer_auto_out_a_bits_address; // @[TLTraceBuffer.scala 47:34]
  wire [31:0] trace_buffer_auto_out_a_bits_mask; // @[TLTraceBuffer.scala 47:34]
  wire [255:0] trace_buffer_auto_out_a_bits_data; // @[TLTraceBuffer.scala 47:34]
  wire  trace_buffer_auto_out_b_ready; // @[TLTraceBuffer.scala 47:34]
  wire  trace_buffer_auto_out_b_valid; // @[TLTraceBuffer.scala 47:34]
  wire [2:0] trace_buffer_auto_out_b_bits_size; // @[TLTraceBuffer.scala 47:34]
  wire [3:0] trace_buffer_auto_out_b_bits_source; // @[TLTraceBuffer.scala 47:34]
  wire [31:0] trace_buffer_auto_out_b_bits_address; // @[TLTraceBuffer.scala 47:34]
  wire  trace_buffer_auto_out_c_ready; // @[TLTraceBuffer.scala 47:34]
  wire  trace_buffer_auto_out_c_valid; // @[TLTraceBuffer.scala 47:34]
  wire [2:0] trace_buffer_auto_out_c_bits_opcode; // @[TLTraceBuffer.scala 47:34]
  wire [2:0] trace_buffer_auto_out_c_bits_param; // @[TLTraceBuffer.scala 47:34]
  wire [2:0] trace_buffer_auto_out_c_bits_size; // @[TLTraceBuffer.scala 47:34]
  wire [3:0] trace_buffer_auto_out_c_bits_source; // @[TLTraceBuffer.scala 47:34]
  wire [31:0] trace_buffer_auto_out_c_bits_address; // @[TLTraceBuffer.scala 47:34]
  wire [255:0] trace_buffer_auto_out_c_bits_data; // @[TLTraceBuffer.scala 47:34]
  wire  trace_buffer_auto_out_d_ready; // @[TLTraceBuffer.scala 47:34]
  wire  trace_buffer_auto_out_d_valid; // @[TLTraceBuffer.scala 47:34]
  wire [2:0] trace_buffer_auto_out_d_bits_opcode; // @[TLTraceBuffer.scala 47:34]
  wire [2:0] trace_buffer_auto_out_d_bits_size; // @[TLTraceBuffer.scala 47:34]
  wire [3:0] trace_buffer_auto_out_d_bits_source; // @[TLTraceBuffer.scala 47:34]
  wire [5:0] trace_buffer_auto_out_d_bits_sink; // @[TLTraceBuffer.scala 47:34]
  wire [255:0] trace_buffer_auto_out_d_bits_data; // @[TLTraceBuffer.scala 47:34]
  wire  trace_buffer_auto_out_e_ready; // @[TLTraceBuffer.scala 47:34]
  wire  trace_buffer_auto_out_e_valid; // @[TLTraceBuffer.scala 47:34]
  wire [5:0] trace_buffer_auto_out_e_bits_sink; // @[TLTraceBuffer.scala 47:34]
  wire  in_fifo_io_enq_clock; // @[SoC.scala 111:26]
  wire  in_fifo_io_enq_reset; // @[SoC.scala 111:26]
  wire  in_fifo_io_enq_ready; // @[SoC.scala 111:26]
  wire  in_fifo_io_enq_valid; // @[SoC.scala 111:26]
  wire [7:0] in_fifo_io_enq_bits; // @[SoC.scala 111:26]
  wire  in_fifo_io_deq_clock; // @[SoC.scala 111:26]
  wire  in_fifo_io_deq_reset; // @[SoC.scala 111:26]
  wire  in_fifo_io_deq_ready; // @[SoC.scala 111:26]
  wire  in_fifo_io_deq_valid; // @[SoC.scala 111:26]
  wire [7:0] in_fifo_io_deq_bits; // @[SoC.scala 111:26]
  wire  out_fifo_io_enq_clock; // @[SoC.scala 112:26]
  wire  out_fifo_io_enq_reset; // @[SoC.scala 112:26]
  wire  out_fifo_io_enq_ready; // @[SoC.scala 112:26]
  wire  out_fifo_io_enq_valid; // @[SoC.scala 112:26]
  wire [7:0] out_fifo_io_enq_bits; // @[SoC.scala 112:26]
  wire  out_fifo_io_deq_clock; // @[SoC.scala 112:26]
  wire  out_fifo_io_deq_reset; // @[SoC.scala 112:26]
  wire  out_fifo_io_deq_ready; // @[SoC.scala 112:26]
  wire  out_fifo_io_deq_valid; // @[SoC.scala 112:26]
  wire [7:0] out_fifo_io_deq_bits; // @[SoC.scala 112:26]
  reg  sync_dff_0_mtip; // @[SoC.scala 127:27]
  reg  sync_dff_0_msip; // @[SoC.scala 127:27]
  reg  sync_dff_0_meip; // @[SoC.scala 127:27]
  reg  sync_dff_0_seip; // @[SoC.scala 127:27]
  reg  sync_dff_1_mtip; // @[SoC.scala 127:27]
  reg  sync_dff_1_msip; // @[SoC.scala 127:27]
  reg  sync_dff_1_meip; // @[SoC.scala 127:27]
  reg  sync_dff_1_seip; // @[SoC.scala 127:27]
  reg  sync_dff_2_mtip; // @[SoC.scala 127:27]
  reg  sync_dff_2_msip; // @[SoC.scala 127:27]
  reg  sync_dff_2_meip; // @[SoC.scala 127:27]
  reg  sync_dff_2_seip; // @[SoC.scala 127:27]
  SoCImp soc_imp ( // @[SoC.scala 81:27]
    .clock(soc_imp_clock),
    .reset(soc_imp_reset),
    .auto_out_a_ready(soc_imp_auto_out_a_ready),
    .auto_out_a_valid(soc_imp_auto_out_a_valid),
    .auto_out_a_bits_opcode(soc_imp_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(soc_imp_auto_out_a_bits_param),
    .auto_out_a_bits_size(soc_imp_auto_out_a_bits_size),
    .auto_out_a_bits_source(soc_imp_auto_out_a_bits_source),
    .auto_out_a_bits_address(soc_imp_auto_out_a_bits_address),
    .auto_out_a_bits_mask(soc_imp_auto_out_a_bits_mask),
    .auto_out_a_bits_data(soc_imp_auto_out_a_bits_data),
    .auto_out_b_ready(soc_imp_auto_out_b_ready),
    .auto_out_b_valid(soc_imp_auto_out_b_valid),
    .auto_out_b_bits_size(soc_imp_auto_out_b_bits_size),
    .auto_out_b_bits_source(soc_imp_auto_out_b_bits_source),
    .auto_out_b_bits_address(soc_imp_auto_out_b_bits_address),
    .auto_out_c_ready(soc_imp_auto_out_c_ready),
    .auto_out_c_valid(soc_imp_auto_out_c_valid),
    .auto_out_c_bits_opcode(soc_imp_auto_out_c_bits_opcode),
    .auto_out_c_bits_param(soc_imp_auto_out_c_bits_param),
    .auto_out_c_bits_size(soc_imp_auto_out_c_bits_size),
    .auto_out_c_bits_source(soc_imp_auto_out_c_bits_source),
    .auto_out_c_bits_address(soc_imp_auto_out_c_bits_address),
    .auto_out_c_bits_data(soc_imp_auto_out_c_bits_data),
    .auto_out_d_ready(soc_imp_auto_out_d_ready),
    .auto_out_d_valid(soc_imp_auto_out_d_valid),
    .auto_out_d_bits_opcode(soc_imp_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(soc_imp_auto_out_d_bits_size),
    .auto_out_d_bits_source(soc_imp_auto_out_d_bits_source),
    .auto_out_d_bits_sink(soc_imp_auto_out_d_bits_sink),
    .auto_out_d_bits_data(soc_imp_auto_out_d_bits_data),
    .auto_out_e_ready(soc_imp_auto_out_e_ready),
    .auto_out_e_valid(soc_imp_auto_out_e_valid),
    .auto_out_e_bits_sink(soc_imp_auto_out_e_bits_sink),
    .io_intr_mtip(soc_imp_io_intr_mtip),
    .io_intr_msip(soc_imp_io_intr_msip),
    .io_intr_meip(soc_imp_io_intr_meip),
    .io_intr_seip(soc_imp_io_intr_seip)
  );
  TLSerdes serdes ( // @[SoC.scala 87:26]
    .clock(serdes_clock),
    .reset(serdes_reset),
    .auto_in_a_ready(serdes_auto_in_a_ready),
    .auto_in_a_valid(serdes_auto_in_a_valid),
    .auto_in_a_bits_opcode(serdes_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(serdes_auto_in_a_bits_param),
    .auto_in_a_bits_size(serdes_auto_in_a_bits_size),
    .auto_in_a_bits_source(serdes_auto_in_a_bits_source),
    .auto_in_a_bits_address(serdes_auto_in_a_bits_address),
    .auto_in_a_bits_mask(serdes_auto_in_a_bits_mask),
    .auto_in_a_bits_data(serdes_auto_in_a_bits_data),
    .auto_in_b_ready(serdes_auto_in_b_ready),
    .auto_in_b_valid(serdes_auto_in_b_valid),
    .auto_in_b_bits_size(serdes_auto_in_b_bits_size),
    .auto_in_b_bits_source(serdes_auto_in_b_bits_source),
    .auto_in_b_bits_address(serdes_auto_in_b_bits_address),
    .auto_in_c_ready(serdes_auto_in_c_ready),
    .auto_in_c_valid(serdes_auto_in_c_valid),
    .auto_in_c_bits_opcode(serdes_auto_in_c_bits_opcode),
    .auto_in_c_bits_param(serdes_auto_in_c_bits_param),
    .auto_in_c_bits_size(serdes_auto_in_c_bits_size),
    .auto_in_c_bits_source(serdes_auto_in_c_bits_source),
    .auto_in_c_bits_address(serdes_auto_in_c_bits_address),
    .auto_in_c_bits_data(serdes_auto_in_c_bits_data),
    .auto_in_d_ready(serdes_auto_in_d_ready),
    .auto_in_d_valid(serdes_auto_in_d_valid),
    .auto_in_d_bits_opcode(serdes_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(serdes_auto_in_d_bits_size),
    .auto_in_d_bits_source(serdes_auto_in_d_bits_source),
    .auto_in_d_bits_sink(serdes_auto_in_d_bits_sink),
    .auto_in_d_bits_data(serdes_auto_in_d_bits_data),
    .auto_in_e_ready(serdes_auto_in_e_ready),
    .auto_in_e_valid(serdes_auto_in_e_valid),
    .auto_in_e_bits_sink(serdes_auto_in_e_bits_sink),
    .io_ser_0_in_ready(serdes_io_ser_0_in_ready),
    .io_ser_0_in_valid(serdes_io_ser_0_in_valid),
    .io_ser_0_in_bits(serdes_io_ser_0_in_bits),
    .io_ser_0_out_ready(serdes_io_ser_0_out_ready),
    .io_ser_0_out_valid(serdes_io_ser_0_out_valid),
    .io_ser_0_out_bits(serdes_io_ser_0_out_bits)
  );
  TLTraceBuffer trace_buffer ( // @[TLTraceBuffer.scala 47:34]
    .clock(trace_buffer_clock),
    .reset(trace_buffer_reset),
    .auto_in_a_ready(trace_buffer_auto_in_a_ready),
    .auto_in_a_valid(trace_buffer_auto_in_a_valid),
    .auto_in_a_bits_opcode(trace_buffer_auto_in_a_bits_opcode),
    .auto_in_a_bits_param(trace_buffer_auto_in_a_bits_param),
    .auto_in_a_bits_size(trace_buffer_auto_in_a_bits_size),
    .auto_in_a_bits_source(trace_buffer_auto_in_a_bits_source),
    .auto_in_a_bits_address(trace_buffer_auto_in_a_bits_address),
    .auto_in_a_bits_mask(trace_buffer_auto_in_a_bits_mask),
    .auto_in_a_bits_data(trace_buffer_auto_in_a_bits_data),
    .auto_in_b_ready(trace_buffer_auto_in_b_ready),
    .auto_in_b_valid(trace_buffer_auto_in_b_valid),
    .auto_in_b_bits_size(trace_buffer_auto_in_b_bits_size),
    .auto_in_b_bits_source(trace_buffer_auto_in_b_bits_source),
    .auto_in_b_bits_address(trace_buffer_auto_in_b_bits_address),
    .auto_in_c_ready(trace_buffer_auto_in_c_ready),
    .auto_in_c_valid(trace_buffer_auto_in_c_valid),
    .auto_in_c_bits_opcode(trace_buffer_auto_in_c_bits_opcode),
    .auto_in_c_bits_param(trace_buffer_auto_in_c_bits_param),
    .auto_in_c_bits_size(trace_buffer_auto_in_c_bits_size),
    .auto_in_c_bits_source(trace_buffer_auto_in_c_bits_source),
    .auto_in_c_bits_address(trace_buffer_auto_in_c_bits_address),
    .auto_in_c_bits_data(trace_buffer_auto_in_c_bits_data),
    .auto_in_d_ready(trace_buffer_auto_in_d_ready),
    .auto_in_d_valid(trace_buffer_auto_in_d_valid),
    .auto_in_d_bits_opcode(trace_buffer_auto_in_d_bits_opcode),
    .auto_in_d_bits_size(trace_buffer_auto_in_d_bits_size),
    .auto_in_d_bits_source(trace_buffer_auto_in_d_bits_source),
    .auto_in_d_bits_sink(trace_buffer_auto_in_d_bits_sink),
    .auto_in_d_bits_data(trace_buffer_auto_in_d_bits_data),
    .auto_in_e_ready(trace_buffer_auto_in_e_ready),
    .auto_in_e_valid(trace_buffer_auto_in_e_valid),
    .auto_in_e_bits_sink(trace_buffer_auto_in_e_bits_sink),
    .auto_out_a_ready(trace_buffer_auto_out_a_ready),
    .auto_out_a_valid(trace_buffer_auto_out_a_valid),
    .auto_out_a_bits_opcode(trace_buffer_auto_out_a_bits_opcode),
    .auto_out_a_bits_param(trace_buffer_auto_out_a_bits_param),
    .auto_out_a_bits_size(trace_buffer_auto_out_a_bits_size),
    .auto_out_a_bits_source(trace_buffer_auto_out_a_bits_source),
    .auto_out_a_bits_address(trace_buffer_auto_out_a_bits_address),
    .auto_out_a_bits_mask(trace_buffer_auto_out_a_bits_mask),
    .auto_out_a_bits_data(trace_buffer_auto_out_a_bits_data),
    .auto_out_b_ready(trace_buffer_auto_out_b_ready),
    .auto_out_b_valid(trace_buffer_auto_out_b_valid),
    .auto_out_b_bits_size(trace_buffer_auto_out_b_bits_size),
    .auto_out_b_bits_source(trace_buffer_auto_out_b_bits_source),
    .auto_out_b_bits_address(trace_buffer_auto_out_b_bits_address),
    .auto_out_c_ready(trace_buffer_auto_out_c_ready),
    .auto_out_c_valid(trace_buffer_auto_out_c_valid),
    .auto_out_c_bits_opcode(trace_buffer_auto_out_c_bits_opcode),
    .auto_out_c_bits_param(trace_buffer_auto_out_c_bits_param),
    .auto_out_c_bits_size(trace_buffer_auto_out_c_bits_size),
    .auto_out_c_bits_source(trace_buffer_auto_out_c_bits_source),
    .auto_out_c_bits_address(trace_buffer_auto_out_c_bits_address),
    .auto_out_c_bits_data(trace_buffer_auto_out_c_bits_data),
    .auto_out_d_ready(trace_buffer_auto_out_d_ready),
    .auto_out_d_valid(trace_buffer_auto_out_d_valid),
    .auto_out_d_bits_opcode(trace_buffer_auto_out_d_bits_opcode),
    .auto_out_d_bits_size(trace_buffer_auto_out_d_bits_size),
    .auto_out_d_bits_source(trace_buffer_auto_out_d_bits_source),
    .auto_out_d_bits_sink(trace_buffer_auto_out_d_bits_sink),
    .auto_out_d_bits_data(trace_buffer_auto_out_d_bits_data),
    .auto_out_e_ready(trace_buffer_auto_out_e_ready),
    .auto_out_e_valid(trace_buffer_auto_out_e_valid),
    .auto_out_e_bits_sink(trace_buffer_auto_out_e_bits_sink)
  );
  AsyncQueue in_fifo ( // @[SoC.scala 111:26]
    .io_enq_clock(in_fifo_io_enq_clock),
    .io_enq_reset(in_fifo_io_enq_reset),
    .io_enq_ready(in_fifo_io_enq_ready),
    .io_enq_valid(in_fifo_io_enq_valid),
    .io_enq_bits(in_fifo_io_enq_bits),
    .io_deq_clock(in_fifo_io_deq_clock),
    .io_deq_reset(in_fifo_io_deq_reset),
    .io_deq_ready(in_fifo_io_deq_ready),
    .io_deq_valid(in_fifo_io_deq_valid),
    .io_deq_bits(in_fifo_io_deq_bits)
  );
  AsyncQueue out_fifo ( // @[SoC.scala 112:26]
    .io_enq_clock(out_fifo_io_enq_clock),
    .io_enq_reset(out_fifo_io_enq_reset),
    .io_enq_ready(out_fifo_io_enq_ready),
    .io_enq_valid(out_fifo_io_enq_valid),
    .io_enq_bits(out_fifo_io_enq_bits),
    .io_deq_clock(out_fifo_io_deq_clock),
    .io_deq_reset(out_fifo_io_deq_reset),
    .io_deq_ready(out_fifo_io_deq_ready),
    .io_deq_valid(out_fifo_io_deq_valid),
    .io_deq_bits(out_fifo_io_deq_bits)
  );
  assign io_in_ready = in_fifo_io_enq_ready; // @[SoC.scala 113:27]
  assign io_out_valid = out_fifo_io_deq_valid; // @[SoC.scala 122:27]
  assign io_out_bits = out_fifo_io_deq_bits; // @[SoC.scala 122:27]
  assign soc_imp_clock = clock;
  assign soc_imp_reset = reset;
  assign soc_imp_auto_out_a_ready = trace_buffer_auto_in_a_ready; // @[LazyModule.scala 355:16]
  assign soc_imp_auto_out_b_valid = trace_buffer_auto_in_b_valid; // @[LazyModule.scala 355:16]
  assign soc_imp_auto_out_b_bits_size = trace_buffer_auto_in_b_bits_size; // @[LazyModule.scala 355:16]
  assign soc_imp_auto_out_b_bits_source = trace_buffer_auto_in_b_bits_source; // @[LazyModule.scala 355:16]
  assign soc_imp_auto_out_b_bits_address = trace_buffer_auto_in_b_bits_address; // @[LazyModule.scala 355:16]
  assign soc_imp_auto_out_c_ready = trace_buffer_auto_in_c_ready; // @[LazyModule.scala 355:16]
  assign soc_imp_auto_out_d_valid = trace_buffer_auto_in_d_valid; // @[LazyModule.scala 355:16]
  assign soc_imp_auto_out_d_bits_opcode = trace_buffer_auto_in_d_bits_opcode; // @[LazyModule.scala 355:16]
  assign soc_imp_auto_out_d_bits_size = trace_buffer_auto_in_d_bits_size; // @[LazyModule.scala 355:16]
  assign soc_imp_auto_out_d_bits_source = trace_buffer_auto_in_d_bits_source; // @[LazyModule.scala 355:16]
  assign soc_imp_auto_out_d_bits_sink = trace_buffer_auto_in_d_bits_sink; // @[LazyModule.scala 355:16]
  assign soc_imp_auto_out_d_bits_data = trace_buffer_auto_in_d_bits_data; // @[LazyModule.scala 355:16]
  assign soc_imp_auto_out_e_ready = trace_buffer_auto_in_e_ready; // @[LazyModule.scala 355:16]
  assign soc_imp_io_intr_mtip = sync_dff_2_mtip; // @[SoC.scala 131:28]
  assign soc_imp_io_intr_msip = sync_dff_2_msip; // @[SoC.scala 131:28]
  assign soc_imp_io_intr_meip = sync_dff_2_meip; // @[SoC.scala 131:28]
  assign soc_imp_io_intr_seip = sync_dff_2_seip; // @[SoC.scala 131:28]
  assign serdes_clock = clock;
  assign serdes_reset = reset;
  assign serdes_auto_in_a_valid = trace_buffer_auto_out_a_valid; // @[LazyModule.scala 353:16]
  assign serdes_auto_in_a_bits_opcode = trace_buffer_auto_out_a_bits_opcode; // @[LazyModule.scala 353:16]
  assign serdes_auto_in_a_bits_param = trace_buffer_auto_out_a_bits_param; // @[LazyModule.scala 353:16]
  assign serdes_auto_in_a_bits_size = trace_buffer_auto_out_a_bits_size; // @[LazyModule.scala 353:16]
  assign serdes_auto_in_a_bits_source = trace_buffer_auto_out_a_bits_source; // @[LazyModule.scala 353:16]
  assign serdes_auto_in_a_bits_address = trace_buffer_auto_out_a_bits_address; // @[LazyModule.scala 353:16]
  assign serdes_auto_in_a_bits_mask = trace_buffer_auto_out_a_bits_mask; // @[LazyModule.scala 353:16]
  assign serdes_auto_in_a_bits_data = trace_buffer_auto_out_a_bits_data; // @[LazyModule.scala 353:16]
  assign serdes_auto_in_b_ready = trace_buffer_auto_out_b_ready; // @[LazyModule.scala 353:16]
  assign serdes_auto_in_c_valid = trace_buffer_auto_out_c_valid; // @[LazyModule.scala 353:16]
  assign serdes_auto_in_c_bits_opcode = trace_buffer_auto_out_c_bits_opcode; // @[LazyModule.scala 353:16]
  assign serdes_auto_in_c_bits_param = trace_buffer_auto_out_c_bits_param; // @[LazyModule.scala 353:16]
  assign serdes_auto_in_c_bits_size = trace_buffer_auto_out_c_bits_size; // @[LazyModule.scala 353:16]
  assign serdes_auto_in_c_bits_source = trace_buffer_auto_out_c_bits_source; // @[LazyModule.scala 353:16]
  assign serdes_auto_in_c_bits_address = trace_buffer_auto_out_c_bits_address; // @[LazyModule.scala 353:16]
  assign serdes_auto_in_c_bits_data = trace_buffer_auto_out_c_bits_data; // @[LazyModule.scala 353:16]
  assign serdes_auto_in_d_ready = trace_buffer_auto_out_d_ready; // @[LazyModule.scala 353:16]
  assign serdes_auto_in_e_valid = trace_buffer_auto_out_e_valid; // @[LazyModule.scala 353:16]
  assign serdes_auto_in_e_bits_sink = trace_buffer_auto_out_e_bits_sink; // @[LazyModule.scala 353:16]
  assign serdes_io_ser_0_in_valid = in_fifo_io_deq_valid; // @[SoC.scala 116:27]
  assign serdes_io_ser_0_in_bits = in_fifo_io_deq_bits; // @[SoC.scala 116:27]
  assign serdes_io_ser_0_out_ready = out_fifo_io_enq_ready; // @[SoC.scala 119:27]
  assign trace_buffer_clock = clock;
  assign trace_buffer_reset = reset;
  assign trace_buffer_auto_in_a_valid = soc_imp_auto_out_a_valid; // @[LazyModule.scala 355:16]
  assign trace_buffer_auto_in_a_bits_opcode = soc_imp_auto_out_a_bits_opcode; // @[LazyModule.scala 355:16]
  assign trace_buffer_auto_in_a_bits_param = soc_imp_auto_out_a_bits_param; // @[LazyModule.scala 355:16]
  assign trace_buffer_auto_in_a_bits_size = soc_imp_auto_out_a_bits_size; // @[LazyModule.scala 355:16]
  assign trace_buffer_auto_in_a_bits_source = soc_imp_auto_out_a_bits_source; // @[LazyModule.scala 355:16]
  assign trace_buffer_auto_in_a_bits_address = soc_imp_auto_out_a_bits_address; // @[LazyModule.scala 355:16]
  assign trace_buffer_auto_in_a_bits_mask = soc_imp_auto_out_a_bits_mask; // @[LazyModule.scala 355:16]
  assign trace_buffer_auto_in_a_bits_data = soc_imp_auto_out_a_bits_data; // @[LazyModule.scala 355:16]
  assign trace_buffer_auto_in_b_ready = soc_imp_auto_out_b_ready; // @[LazyModule.scala 355:16]
  assign trace_buffer_auto_in_c_valid = soc_imp_auto_out_c_valid; // @[LazyModule.scala 355:16]
  assign trace_buffer_auto_in_c_bits_opcode = soc_imp_auto_out_c_bits_opcode; // @[LazyModule.scala 355:16]
  assign trace_buffer_auto_in_c_bits_param = soc_imp_auto_out_c_bits_param; // @[LazyModule.scala 355:16]
  assign trace_buffer_auto_in_c_bits_size = soc_imp_auto_out_c_bits_size; // @[LazyModule.scala 355:16]
  assign trace_buffer_auto_in_c_bits_source = soc_imp_auto_out_c_bits_source; // @[LazyModule.scala 355:16]
  assign trace_buffer_auto_in_c_bits_address = soc_imp_auto_out_c_bits_address; // @[LazyModule.scala 355:16]
  assign trace_buffer_auto_in_c_bits_data = soc_imp_auto_out_c_bits_data; // @[LazyModule.scala 355:16]
  assign trace_buffer_auto_in_d_ready = soc_imp_auto_out_d_ready; // @[LazyModule.scala 355:16]
  assign trace_buffer_auto_in_e_valid = soc_imp_auto_out_e_valid; // @[LazyModule.scala 355:16]
  assign trace_buffer_auto_in_e_bits_sink = soc_imp_auto_out_e_bits_sink; // @[LazyModule.scala 355:16]
  assign trace_buffer_auto_out_a_ready = serdes_auto_in_a_ready; // @[LazyModule.scala 353:16]
  assign trace_buffer_auto_out_b_valid = serdes_auto_in_b_valid; // @[LazyModule.scala 353:16]
  assign trace_buffer_auto_out_b_bits_size = serdes_auto_in_b_bits_size; // @[LazyModule.scala 353:16]
  assign trace_buffer_auto_out_b_bits_source = serdes_auto_in_b_bits_source; // @[LazyModule.scala 353:16]
  assign trace_buffer_auto_out_b_bits_address = serdes_auto_in_b_bits_address; // @[LazyModule.scala 353:16]
  assign trace_buffer_auto_out_c_ready = serdes_auto_in_c_ready; // @[LazyModule.scala 353:16]
  assign trace_buffer_auto_out_d_valid = serdes_auto_in_d_valid; // @[LazyModule.scala 353:16]
  assign trace_buffer_auto_out_d_bits_opcode = serdes_auto_in_d_bits_opcode; // @[LazyModule.scala 353:16]
  assign trace_buffer_auto_out_d_bits_size = serdes_auto_in_d_bits_size; // @[LazyModule.scala 353:16]
  assign trace_buffer_auto_out_d_bits_source = serdes_auto_in_d_bits_source; // @[LazyModule.scala 353:16]
  assign trace_buffer_auto_out_d_bits_sink = serdes_auto_in_d_bits_sink; // @[LazyModule.scala 353:16]
  assign trace_buffer_auto_out_d_bits_data = serdes_auto_in_d_bits_data; // @[LazyModule.scala 353:16]
  assign trace_buffer_auto_out_e_ready = serdes_auto_in_e_ready; // @[LazyModule.scala 353:16]
  assign in_fifo_io_enq_clock = io_io_clock; // @[SoC.scala 114:27]
  assign in_fifo_io_enq_reset = io_io_reset; // @[SoC.scala 115:27]
  assign in_fifo_io_enq_valid = io_in_valid; // @[SoC.scala 113:27]
  assign in_fifo_io_enq_bits = io_in_bits; // @[SoC.scala 113:27]
  assign in_fifo_io_deq_clock = clock; // @[SoC.scala 117:27]
  assign in_fifo_io_deq_reset = reset; // @[SoC.scala 118:27]
  assign in_fifo_io_deq_ready = serdes_io_ser_0_in_ready; // @[SoC.scala 116:27]
  assign out_fifo_io_enq_clock = clock; // @[SoC.scala 120:27]
  assign out_fifo_io_enq_reset = reset; // @[SoC.scala 121:27]
  assign out_fifo_io_enq_valid = serdes_io_ser_0_out_valid; // @[SoC.scala 119:27]
  assign out_fifo_io_enq_bits = serdes_io_ser_0_out_bits; // @[SoC.scala 119:27]
  assign out_fifo_io_deq_clock = io_io_clock; // @[SoC.scala 123:27]
  assign out_fifo_io_deq_reset = io_io_reset; // @[SoC.scala 124:27]
  assign out_fifo_io_deq_ready = io_out_ready; // @[SoC.scala 122:27]
  always @(posedge clock) begin
    if (reset) begin // @[SoC.scala 127:27]
      sync_dff_0_mtip <= 1'h0; // @[SoC.scala 127:27]
    end else begin
      sync_dff_0_mtip <= io_intr_mtip; // @[SoC.scala 128:28]
    end
    if (reset) begin // @[SoC.scala 127:27]
      sync_dff_0_msip <= 1'h0; // @[SoC.scala 127:27]
    end else begin
      sync_dff_0_msip <= io_intr_msip; // @[SoC.scala 128:28]
    end
    if (reset) begin // @[SoC.scala 127:27]
      sync_dff_0_meip <= 1'h0; // @[SoC.scala 127:27]
    end else begin
      sync_dff_0_meip <= io_intr_meip; // @[SoC.scala 128:28]
    end
    if (reset) begin // @[SoC.scala 127:27]
      sync_dff_0_seip <= 1'h0; // @[SoC.scala 127:27]
    end else begin
      sync_dff_0_seip <= io_intr_seip; // @[SoC.scala 128:28]
    end
    if (reset) begin // @[SoC.scala 127:27]
      sync_dff_1_mtip <= 1'h0; // @[SoC.scala 127:27]
    end else begin
      sync_dff_1_mtip <= sync_dff_0_mtip; // @[SoC.scala 129:28]
    end
    if (reset) begin // @[SoC.scala 127:27]
      sync_dff_1_msip <= 1'h0; // @[SoC.scala 127:27]
    end else begin
      sync_dff_1_msip <= sync_dff_0_msip; // @[SoC.scala 129:28]
    end
    if (reset) begin // @[SoC.scala 127:27]
      sync_dff_1_meip <= 1'h0; // @[SoC.scala 127:27]
    end else begin
      sync_dff_1_meip <= sync_dff_0_meip; // @[SoC.scala 129:28]
    end
    if (reset) begin // @[SoC.scala 127:27]
      sync_dff_1_seip <= 1'h0; // @[SoC.scala 127:27]
    end else begin
      sync_dff_1_seip <= sync_dff_0_seip; // @[SoC.scala 129:28]
    end
    if (reset) begin // @[SoC.scala 127:27]
      sync_dff_2_mtip <= 1'h0; // @[SoC.scala 127:27]
    end else begin
      sync_dff_2_mtip <= sync_dff_1_mtip; // @[SoC.scala 130:28]
    end
    if (reset) begin // @[SoC.scala 127:27]
      sync_dff_2_msip <= 1'h0; // @[SoC.scala 127:27]
    end else begin
      sync_dff_2_msip <= sync_dff_1_msip; // @[SoC.scala 130:28]
    end
    if (reset) begin // @[SoC.scala 127:27]
      sync_dff_2_meip <= 1'h0; // @[SoC.scala 127:27]
    end else begin
      sync_dff_2_meip <= sync_dff_1_meip; // @[SoC.scala 130:28]
    end
    if (reset) begin // @[SoC.scala 127:27]
      sync_dff_2_seip <= 1'h0; // @[SoC.scala 127:27]
    end else begin
      sync_dff_2_seip <= sync_dff_1_seip; // @[SoC.scala 130:28]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sync_dff_0_mtip = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  sync_dff_0_msip = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  sync_dff_0_meip = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  sync_dff_0_seip = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  sync_dff_1_mtip = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  sync_dff_1_msip = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  sync_dff_1_meip = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  sync_dff_1_seip = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  sync_dff_2_mtip = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  sync_dff_2_msip = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  sync_dff_2_meip = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  sync_dff_2_seip = _RAND_11[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
